

    module v$ROM1_3190(q, a, clk);
    output reg [15:0] q;
    input clk;
    input [9:0] a;
    reg [15:0] rom [1023:0];
    always @(posedge clk) q <= rom[a];
    integer i;
    initial
    begin
        for (i=0; i < 1024; i=i+1)
        begin
            rom[i] = 0;
        end
    
        
    end
    endmodule
     

    module v$ROM1_7586(q, a, clk);
    output reg [15:0] q;
    input clk;
    input [9:0] a;
    reg [15:0] rom [1023:0];
    always @(posedge clk) q <= rom[a];
    integer i;
    initial
    begin
        for (i=0; i < 1024; i=i+1)
        begin
            rom[i] = 0;
        end
    
        
    end
    endmodule
     

    module v$RAM1_13483(q, a, d, we, clk);
    output reg [15:0] q;
    input [15:0] d;
    input [11:0] a;
    input we, clk;
    reg [15:0] ram [4095:0];
     always @(posedge clk) begin
         if (we)
             ram[a] <= d;
         q <= ram[a];
     end

    integer i;
    initial
    begin
        for (i=0; i < 4096; i=i+1)
        begin
            ram[i] = 0;
        end

        ram[0] = 4080;
ram[1] = 4059;
ram[2] = 16201;
ram[3] = 43691;
ram[4] = 15914;
ram[5] = 0;
ram[6] = 0;
ram[7] = 34953;
ram[8] = 15368;
ram[9] = 0;
ram[10] = 0;
ram[11] = 5120;
ram[12] = 14672;
ram[13] = 0;
ram[14] = 0;
ram[15] = 0;
ram[18] = 15944;
ram[19] = 12629;
ram[20] = 0;
ram[21] = 8260;
ram[22] = 0;
ram[23] = 5120;
ram[4080] = 14920;
ram[4081] = 12629;
ram[4082] = 0;
ram[4083] = 8260;
ram[4084] = 0;
ram[4085] = 0;
    end
    endmodule

    

    module v$AROM1_16768(q, a);
    output[43:0] q;
    input [5:0] a;
    reg [43:0] rom [63:0];

    assign q = rom[a];
    integer i;
    initial
    begin
        for (i=0; i < 64; i=i+1)
        begin
            rom[i] = 0;
        end
    
        rom[0] = 1030792151295;
rom[1] = 64424509695;
rom[2] = 1095216660735;
rom[3] = 4026532095;
rom[4] = 1034818683135;
rom[5] = 68451041535;
rom[6] = 1099243192575;
rom[7] = 251658495;
rom[8] = 1031043809535;
rom[9] = 64676167935;
rom[10] = 0;
    end
    endmodule
     

    module v$AROM1_16769(q, a);
    output[43:0] q;
    input [5:0] a;
    reg [43:0] rom [63:0];

    assign q = rom[a];
    integer i;
    initial
    begin
        for (i=0; i < 64; i=i+1)
        begin
            rom[i] = 0;
        end
    
        rom[0] = 1030792151295;
rom[1] = 64424509695;
rom[2] = 1095216660735;
rom[3] = 4026532095;
rom[4] = 1034818683135;
rom[5] = 68451041535;
rom[6] = 1099243192575;
rom[7] = 251658495;
rom[8] = 1031043809535;
rom[9] = 64676167935;
rom[10] = 0;
    end
    endmodule
     
module main (
	clk,
	v$PC0_8220_out0,
	v$PC1_12778_out0);
input clk;
output  [11:0] v$PC0_8220_out0;
output  [11:0] v$PC1_12778_out0;
reg  [11:0] v$INT0_16488_out0 = 12'h0;
reg  [11:0] v$INT0_16489_out0 = 12'h0;
reg  [11:0] v$INT1_19145_out0 = 12'h0;
reg  [11:0] v$INT1_19146_out0 = 12'h0;
reg  [11:0] v$INT2_265_out0 = 12'h0;
reg  [11:0] v$INT2_266_out0 = 12'h0;
reg  [11:0] v$INT3_281_out0 = 12'h0;
reg  [11:0] v$INT3_282_out0 = 12'h0;
reg  [11:0] v$PCINTERRUPT_18413_out0 = 12'h0;
reg  [11:0] v$PCINTERRUPT_18414_out0 = 12'h0;
reg  [11:0] v$PCNORMAL_13337_out0 = 12'h0;
reg  [11:0] v$PCNORMAL_13338_out0 = 12'h0;
reg  [11:0] v$REG12_3553_out0 = 12'h0;
reg  [11:0] v$REG9_16701_out0 = 12'h0;
reg  [15:0] v$REG0_16864_out0 = 16'h0;
reg  [15:0] v$REG0_16865_out0 = 16'h0;
reg  [15:0] v$REG10_17089_out0 = 16'h0;
reg  [15:0] v$REG11_10004_out0 = 16'h0;
reg  [15:0] v$REG1_1309_out0 = 16'h0;
reg  [15:0] v$REG1_1310_out0 = 16'h0;
reg  [15:0] v$REG1_14166_out0 = 16'h0;
reg  [15:0] v$REG1_14167_out0 = 16'h0;
reg  [15:0] v$REG1_14711_out0 = 16'h0;
reg  [15:0] v$REG1_14712_out0 = 16'h0;
reg  [15:0] v$REG1_5110_out0 = 16'h0;
reg  [15:0] v$REG1_5111_out0 = 16'h0;
reg  [15:0] v$REG2_15622_out0 = 16'h0;
reg  [15:0] v$REG2_15623_out0 = 16'h0;
reg  [15:0] v$REG2_16210_out0 = 16'h0;
reg  [15:0] v$REG2_16211_out0 = 16'h0;
reg  [15:0] v$REG2_16962_out0 = 16'h0;
reg  [15:0] v$REG2_16963_out0 = 16'h0;
reg  [15:0] v$REG2_18120_out0 = 16'h0;
reg  [15:0] v$REG2_18121_out0 = 16'h0;
reg  [15:0] v$REG3_11509_out0 = 16'h0;
reg  [15:0] v$REG3_11510_out0 = 16'h0;
reg  [15:0] v$REG3_12336_out0 = 16'h0;
reg  [15:0] v$REG3_12337_out0 = 16'h0;
reg  [15:0] v$REG3_3046_out0 = 16'h0;
reg  [15:0] v$REG3_3047_out0 = 16'h0;
reg  [15:0] v$REG4_6885_out0 = 16'h0;
reg  [15:0] v$REG4_6886_out0 = 16'h0;
reg  [1:0] v$REG1_11407_out0 = 2'h0;
reg  [1:0] v$REG1_11408_out0 = 2'h0;
reg  [1:0] v$REG4_11270_out0 = 2'h0;
reg  [1:0] v$REG4_11271_out0 = 2'h0;
reg  [23:0] v$REG1_12653_out0 = 24'h0;
reg  [23:0] v$REG1_12654_out0 = 24'h0;
reg  [23:0] v$REG2_17420_out0 = 24'h0;
reg  [23:0] v$REG2_17421_out0 = 24'h0;
reg  [31:0] v$REG1_8170_out0 = 32'h0;
reg  [31:0] v$REG1_8171_out0 = 32'h0;
reg  [31:0] v$REG2_4204_out0 = 32'h0;
reg  [31:0] v$REG2_4205_out0 = 32'h0;
reg  [3:0] v$REG1_19272_out0 = 4'h0;
reg  [3:0] v$REG1_19273_out0 = 4'h0;
reg  [3:0] v$REG1_9225_out0 = 4'h0;
reg  [3:0] v$REG1_9226_out0 = 4'h0;
reg  [4:0] v$REG1_14701_out0 = 5'h0;
reg  [4:0] v$REG1_14702_out0 = 5'h0;
reg  [5:0] v$REG1_15444_out0 = 6'h0;
reg  [5:0] v$REG1_15445_out0 = 6'h0;
reg  [5:0] v$REG2_718_out0 = 6'h0;
reg  [5:0] v$REG2_719_out0 = 6'h0;
reg  [7:0] v$REG1_10757_out0 = 8'h0;
reg  [7:0] v$REG1_10758_out0 = 8'h0;
reg  [7:0] v$REG1_4200_out0 = 8'h0;
reg  [7:0] v$REG1_4201_out0 = 8'h0;
reg v$FF0_4488_out0 = 1'b0;
reg v$FF0_4489_out0 = 1'b0;
reg v$FF0_5223_out0 = 1'b0;
reg v$FF0_5224_out0 = 1'b0;
reg v$FF0_716_out0 = 1'b0;
reg v$FF0_717_out0 = 1'b0;
reg v$FF0_9775_out0 = 1'b0;
reg v$FF0_9776_out0 = 1'b0;
reg v$FF10_14804_out0 = 1'b0;
reg v$FF10_14805_out0 = 1'b0;
reg v$FF10_8216_out0 = 1'b0;
reg v$FF10_8217_out0 = 1'b0;
reg v$FF11_2642_out0 = 1'b0;
reg v$FF11_2643_out0 = 1'b0;
reg v$FF12_17048_out0 = 1'b0;
reg v$FF12_17049_out0 = 1'b0;
reg v$FF13_19153_out0 = 1'b0;
reg v$FF13_19154_out0 = 1'b0;
reg v$FF14_11409_out0 = 1'b0;
reg v$FF14_11410_out0 = 1'b0;
reg v$FF15_13286_out0 = 1'b0;
reg v$FF15_13287_out0 = 1'b0;
reg v$FF1_10012_out0 = 1'b0;
reg v$FF1_10013_out0 = 1'b0;
reg v$FF1_10761_out0 = 1'b0;
reg v$FF1_10762_out0 = 1'b0;
reg v$FF1_11566_out0 = 1'b0;
reg v$FF1_11567_out0 = 1'b0;
reg v$FF1_1325_out0 = 1'b0;
reg v$FF1_1326_out0 = 1'b0;
reg v$FF1_13671_out0 = 1'b0;
reg v$FF1_13672_out0 = 1'b0;
reg v$FF1_14261_out0 = 1'b0;
reg v$FF1_14262_out0 = 1'b0;
reg v$FF1_1539_out0 = 1'b0;
reg v$FF1_1540_out0 = 1'b0;
reg v$FF1_16687_out0 = 1'b0;
reg v$FF1_16688_out0 = 1'b0;
reg v$FF1_16689_out0 = 1'b0;
reg v$FF1_16690_out0 = 1'b0;
reg v$FF1_16691_out0 = 1'b0;
reg v$FF1_16692_out0 = 1'b0;
reg v$FF1_16693_out0 = 1'b0;
reg v$FF1_16694_out0 = 1'b0;
reg v$FF1_16695_out0 = 1'b0;
reg v$FF1_16696_out0 = 1'b0;
reg v$FF1_16697_out0 = 1'b0;
reg v$FF1_16698_out0 = 1'b0;
reg v$FF1_16797_out0 = 1'b0;
reg v$FF1_16798_out0 = 1'b0;
reg v$FF1_16930_out0 = 1'b0;
reg v$FF1_16931_out0 = 1'b0;
reg v$FF1_194_out0 = 1'b0;
reg v$FF1_195_out0 = 1'b0;
reg v$FF1_2722_out0 = 1'b0;
reg v$FF1_2723_out0 = 1'b0;
reg v$FF1_2_out0 = 1'b0;
reg v$FF1_3_out0 = 1'b0;
reg v$FF1_4502_out0 = 1'b0;
reg v$FF1_4503_out0 = 1'b0;
reg v$FF1_5439_out0 = 1'b0;
reg v$FF1_5440_out0 = 1'b0;
reg v$FF1_5441_out0 = 1'b0;
reg v$FF1_5442_out0 = 1'b0;
reg v$FF1_5443_out0 = 1'b0;
reg v$FF1_5444_out0 = 1'b0;
reg v$FF1_5688_out0 = 1'b0;
reg v$FF1_6306_out0 = 1'b0;
reg v$FF1_6307_out0 = 1'b0;
reg v$FF1_6414_out0 = 1'b0;
reg v$FF1_6415_out0 = 1'b0;
reg v$FF1_8531_out0 = 1'b0;
reg v$FF1_8532_out0 = 1'b0;
reg v$FF1_9797_out0 = 1'b0;
reg v$FF1_9798_out0 = 1'b0;
reg v$FF1_9988_out0 = 1'b0;
reg v$FF1_9989_out0 = 1'b0;
reg v$FF2_1327_out0 = 1'b0;
reg v$FF2_1328_out0 = 1'b0;
reg v$FF2_13615_out0 = 1'b0;
reg v$FF2_13616_out0 = 1'b0;
reg v$FF2_13617_out0 = 1'b0;
reg v$FF2_13618_out0 = 1'b0;
reg v$FF2_13619_out0 = 1'b0;
reg v$FF2_13620_out0 = 1'b0;
reg v$FF2_13621_out0 = 1'b0;
reg v$FF2_13622_out0 = 1'b0;
reg v$FF2_13623_out0 = 1'b0;
reg v$FF2_13624_out0 = 1'b0;
reg v$FF2_13625_out0 = 1'b0;
reg v$FF2_13626_out0 = 1'b0;
reg v$FF2_13627_out0 = 1'b0;
reg v$FF2_13628_out0 = 1'b0;
reg v$FF2_13629_out0 = 1'b0;
reg v$FF2_13630_out0 = 1'b0;
reg v$FF2_13631_out0 = 1'b0;
reg v$FF2_13632_out0 = 1'b0;
reg v$FF2_13633_out0 = 1'b0;
reg v$FF2_13634_out0 = 1'b0;
reg v$FF2_13635_out0 = 1'b0;
reg v$FF2_13636_out0 = 1'b0;
reg v$FF2_14043_out0 = 1'b0;
reg v$FF2_15233_out0 = 1'b0;
reg v$FF2_15234_out0 = 1'b0;
reg v$FF2_15390_out0 = 1'b0;
reg v$FF2_15391_out0 = 1'b0;
reg v$FF2_15392_out0 = 1'b0;
reg v$FF2_15393_out0 = 1'b0;
reg v$FF2_15394_out0 = 1'b0;
reg v$FF2_15395_out0 = 1'b0;
reg v$FF2_15396_out0 = 1'b0;
reg v$FF2_15397_out0 = 1'b0;
reg v$FF2_15398_out0 = 1'b0;
reg v$FF2_15399_out0 = 1'b0;
reg v$FF2_15400_out0 = 1'b0;
reg v$FF2_15401_out0 = 1'b0;
reg v$FF2_16070_out0 = 1'b0;
reg v$FF2_16071_out0 = 1'b0;
reg v$FF2_16954_out0 = 1'b0;
reg v$FF2_16955_out0 = 1'b0;
reg v$FF2_17272_out0 = 1'b0;
reg v$FF2_17273_out0 = 1'b0;
reg v$FF2_1729_out0 = 1'b0;
reg v$FF2_1730_out0 = 1'b0;
reg v$FF2_3160_out0 = 1'b0;
reg v$FF2_3161_out0 = 1'b0;
reg v$FF2_4510_out0 = 1'b0;
reg v$FF2_4511_out0 = 1'b0;
reg v$FF2_9793_out0 = 1'b0;
reg v$FF2_9794_out0 = 1'b0;
reg v$FF3_10396_out0 = 1'b0;
reg v$FF3_10397_out0 = 1'b0;
reg v$FF3_10398_out0 = 1'b0;
reg v$FF3_10399_out0 = 1'b0;
reg v$FF3_10400_out0 = 1'b0;
reg v$FF3_10401_out0 = 1'b0;
reg v$FF3_10402_out0 = 1'b0;
reg v$FF3_10403_out0 = 1'b0;
reg v$FF3_10404_out0 = 1'b0;
reg v$FF3_10405_out0 = 1'b0;
reg v$FF3_10406_out0 = 1'b0;
reg v$FF3_10407_out0 = 1'b0;
reg v$FF3_11419_out0 = 1'b0;
reg v$FF3_11420_out0 = 1'b0;
reg v$FF3_1456_out0 = 1'b0;
reg v$FF3_1457_out0 = 1'b0;
reg v$FF3_15648_out0 = 1'b0;
reg v$FF3_15649_out0 = 1'b0;
reg v$FF3_16564_out0 = 1'b0;
reg v$FF3_16565_out0 = 1'b0;
reg v$FF3_18727_out0 = 1'b0;
reg v$FF3_18728_out0 = 1'b0;
reg v$FF3_271_out0 = 1'b0;
reg v$FF3_272_out0 = 1'b0;
reg v$FF3_3598_out0 = 1'b0;
reg v$FF3_7649_out0 = 1'b0;
reg v$FF3_7650_out0 = 1'b0;
reg v$FF3_7887_out0 = 1'b0;
reg v$FF3_7888_out0 = 1'b0;
reg v$FF4_14125_out0 = 1'b0;
reg v$FF4_16584_out0 = 1'b0;
reg v$FF4_16585_out0 = 1'b0;
reg v$FF4_16586_out0 = 1'b0;
reg v$FF4_16587_out0 = 1'b0;
reg v$FF4_16588_out0 = 1'b0;
reg v$FF4_16589_out0 = 1'b0;
reg v$FF4_16590_out0 = 1'b0;
reg v$FF4_16591_out0 = 1'b0;
reg v$FF4_16592_out0 = 1'b0;
reg v$FF4_16593_out0 = 1'b0;
reg v$FF4_16594_out0 = 1'b0;
reg v$FF4_16595_out0 = 1'b0;
reg v$FF4_18456_out0 = 1'b0;
reg v$FF4_18457_out0 = 1'b0;
reg v$FF4_19047_out0 = 1'b0;
reg v$FF4_19048_out0 = 1'b0;
reg v$FF4_2541_out0 = 1'b0;
reg v$FF4_2542_out0 = 1'b0;
reg v$FF4_3963_out0 = 1'b0;
reg v$FF4_3964_out0 = 1'b0;
reg v$FF4_7301_out0 = 1'b0;
reg v$FF4_7302_out0 = 1'b0;
reg v$FF4_8369_out0 = 1'b0;
reg v$FF4_8370_out0 = 1'b0;
reg v$FF4_8562_out0 = 1'b0;
reg v$FF4_8563_out0 = 1'b0;
reg v$FF5_16956_out0 = 1'b0;
reg v$FF5_16957_out0 = 1'b0;
reg v$FF5_17047_out0 = 1'b0;
reg v$FF5_19083_out0 = 1'b0;
reg v$FF5_19084_out0 = 1'b0;
reg v$FF5_1915_out0 = 1'b0;
reg v$FF5_1916_out0 = 1'b0;
reg v$FF5_1917_out0 = 1'b0;
reg v$FF5_1918_out0 = 1'b0;
reg v$FF5_1919_out0 = 1'b0;
reg v$FF5_1920_out0 = 1'b0;
reg v$FF5_1921_out0 = 1'b0;
reg v$FF5_1922_out0 = 1'b0;
reg v$FF5_1923_out0 = 1'b0;
reg v$FF5_1924_out0 = 1'b0;
reg v$FF5_1925_out0 = 1'b0;
reg v$FF5_1926_out0 = 1'b0;
reg v$FF5_4957_out0 = 1'b0;
reg v$FF5_4958_out0 = 1'b0;
reg v$FF6_15909_out0 = 1'b0;
reg v$FF6_15910_out0 = 1'b0;
reg v$FF6_16780_out0 = 1'b0;
reg v$FF6_2817_out0 = 1'b0;
reg v$FF6_2818_out0 = 1'b0;
reg v$FF6_2819_out0 = 1'b0;
reg v$FF6_2820_out0 = 1'b0;
reg v$FF6_2821_out0 = 1'b0;
reg v$FF6_2822_out0 = 1'b0;
reg v$FF6_2823_out0 = 1'b0;
reg v$FF6_2824_out0 = 1'b0;
reg v$FF6_2825_out0 = 1'b0;
reg v$FF6_2826_out0 = 1'b0;
reg v$FF6_2827_out0 = 1'b0;
reg v$FF6_2828_out0 = 1'b0;
reg v$FF6_9289_out0 = 1'b0;
reg v$FF6_9290_out0 = 1'b0;
reg v$FF7_13325_out0 = 1'b0;
reg v$FF7_13326_out0 = 1'b0;
reg v$FF7_15152_out0 = 1'b0;
reg v$FF7_15153_out0 = 1'b0;
reg v$FF7_18731_out0 = 1'b0;
reg v$FF7_18732_out0 = 1'b0;
reg v$FF7_8401_out0 = 1'b0;
reg v$FF7_8402_out0 = 1'b0;
reg v$FF7_8609_out0 = 1'b0;
reg v$FF7_8610_out0 = 1'b0;
reg v$FF7_8611_out0 = 1'b0;
reg v$FF7_8612_out0 = 1'b0;
reg v$FF7_8613_out0 = 1'b0;
reg v$FF7_8614_out0 = 1'b0;
reg v$FF7_8615_out0 = 1'b0;
reg v$FF7_8616_out0 = 1'b0;
reg v$FF7_8617_out0 = 1'b0;
reg v$FF7_8618_out0 = 1'b0;
reg v$FF7_8619_out0 = 1'b0;
reg v$FF7_8620_out0 = 1'b0;
reg v$FF8_10797_out0 = 1'b0;
reg v$FF8_10798_out0 = 1'b0;
reg v$FF8_15064_out0 = 1'b0;
reg v$FF8_15065_out0 = 1'b0;
reg v$FF8_15066_out0 = 1'b0;
reg v$FF8_15067_out0 = 1'b0;
reg v$FF8_15068_out0 = 1'b0;
reg v$FF8_15069_out0 = 1'b0;
reg v$FF8_15070_out0 = 1'b0;
reg v$FF8_15071_out0 = 1'b0;
reg v$FF8_15072_out0 = 1'b0;
reg v$FF8_15073_out0 = 1'b0;
reg v$FF8_15074_out0 = 1'b0;
reg v$FF8_15075_out0 = 1'b0;
reg v$FF8_17348_out0 = 1'b0;
reg v$FF8_17349_out0 = 1'b0;
reg v$FF8_8346_out0 = 1'b0;
reg v$FF8_8347_out0 = 1'b0;
reg v$FF9_11158_out0 = 1'b0;
reg v$FF9_11159_out0 = 1'b0;
reg v$FF9_16635_out0 = 1'b0;
reg v$FF9_16636_out0 = 1'b0;
reg v$LSB$FF_19125_out0 = 1'b0;
reg v$LSB$FF_19126_out0 = 1'b0;
reg v$REG13_308_out0 = 1'b0;
reg v$REG14_5698_out0 = 1'b0;
reg v$REG1_7363_out0 = 1'b0;
reg v$REG1_9169_out0 = 1'b0;
reg v$REG2_12370_out0 = 1'b0;
reg v$REG2_12371_out0 = 1'b0;
reg v$REG2_5345_out0 = 1'b0;
reg v$REG3_18364_out0 = 1'b0;
reg v$REG3_18365_out0 = 1'b0;
reg v$REG4_11502_out0 = 1'b0;
reg v$REG7_6442_out0 = 1'b0;
reg v$REG8_4264_out0 = 1'b0;
reg v$S$FF_11312_out0 = 1'b0;
reg v$S$FF_11313_out0 = 1'b0;
wire  [10:0] v$C1_16407_out0;
wire  [10:0] v$C1_16408_out0;
wire  [10:0] v$SEL5_16783_out0;
wire  [10:0] v$SEL5_16784_out0;
wire  [11:0] v$A1_15427_out0;
wire  [11:0] v$A1_15428_out0;
wire  [11:0] v$ADDRESS_15794_out0;
wire  [11:0] v$ADDRESS_16504_out0;
wire  [11:0] v$ADDRESS_16505_out0;
wire  [11:0] v$ADDRESS_2829_out0;
wire  [11:0] v$ADDRESS_6098_out0;
wire  [11:0] v$ADDRESS_6099_out0;
wire  [11:0] v$ADD_3164_out0;
wire  [11:0] v$ADD_3165_out0;
wire  [11:0] v$A_2739_out0;
wire  [11:0] v$A_2740_out0;
wire  [11:0] v$A_2741_out0;
wire  [11:0] v$A_2742_out0;
wire  [11:0] v$B_12696_out0;
wire  [11:0] v$B_12697_out0;
wire  [11:0] v$B_12698_out0;
wire  [11:0] v$B_12699_out0;
wire  [11:0] v$C1_16546_out0;
wire  [11:0] v$C1_16547_out0;
wire  [11:0] v$C4_16509_out0;
wire  [11:0] v$C4_16510_out0;
wire  [11:0] v$END_17218_out0;
wire  [11:0] v$END_17219_out0;
wire  [11:0] v$MUX1_2011_out0;
wire  [11:0] v$MUX2_3903_out0;
wire  [11:0] v$MUX2_3904_out0;
wire  [11:0] v$MUX3_9451_out0;
wire  [11:0] v$MUX4_1731_out0;
wire  [11:0] v$MUX4_1732_out0;
wire  [11:0] v$MUX5_17586_out0;
wire  [11:0] v$MUX5_17587_out0;
wire  [11:0] v$MUX6_15024_out0;
wire  [11:0] v$MUX6_15025_out0;
wire  [11:0] v$MUX6_7182_out0;
wire  [11:0] v$MUX7_1279_out0;
wire  [11:0] v$MUX7_1280_out0;
wire  [11:0] v$MUX8_12853_out0;
wire  [11:0] v$MUX8_12854_out0;
wire  [11:0] v$N$VIEWER_1771_out0;
wire  [11:0] v$N$VIEWER_1772_out0;
wire  [11:0] v$NEXTINSTRUCTIONADDRESS_19015_out0;
wire  [11:0] v$NEXTINSTRUCTIONADDRESS_19016_out0;
wire  [11:0] v$N_12322_out0;
wire  [11:0] v$N_12323_out0;
wire  [11:0] v$N_12539_out0;
wire  [11:0] v$N_12540_out0;
wire  [11:0] v$N_15106_out0;
wire  [11:0] v$N_15107_out0;
wire  [11:0] v$N_15454_out0;
wire  [11:0] v$N_15455_out0;
wire  [11:0] v$N_1777_out0;
wire  [11:0] v$N_1778_out0;
wire  [11:0] v$N_18551_out0;
wire  [11:0] v$N_18552_out0;
wire  [11:0] v$N_18899_out0;
wire  [11:0] v$N_18900_out0;
wire  [11:0] v$N_8578_out0;
wire  [11:0] v$N_8579_out0;
wire  [11:0] v$PC$NEXT0_2098_out0;
wire  [11:0] v$PC$NEXT1_3697_out0;
wire  [11:0] v$PCNEXT$VIEWER_16373_out0;
wire  [11:0] v$PCNEXT$VIEWER_16374_out0;
wire  [11:0] v$PCNEXT_6889_out0;
wire  [11:0] v$PCNEXT_6890_out0;
wire  [11:0] v$PC_3365_out0;
wire  [11:0] v$PC_3366_out0;
wire  [11:0] v$RAM$ADDR$VIEWER_16540_out0;
wire  [11:0] v$RAM$ADDR$VIEWER_16541_out0;
wire  [11:0] v$RAM$ADDR0_13120_out0;
wire  [11:0] v$RAM$ADDR1_6700_out0;
wire  [11:0] v$RAM$ADDR_15811_out0;
wire  [11:0] v$RAM$ADDR_15812_out0;
wire  [11:0] v$RAM$ADDR_6656_out0;
wire  [11:0] v$RAM$ADDR_6657_out0;
wire  [11:0] v$RAMADDR0_17579_out0;
wire  [11:0] v$RAMADDR1_13239_out0;
wire  [11:0] v$RAMADDRESS_13291_out0;
wire  [11:0] v$RAMADDRESS_13292_out0;
wire  [11:0] v$RAMADDRESS_7270_out0;
wire  [11:0] v$RAMADDRESS_7271_out0;
wire  [11:0] v$RAMADDRMUX_14981_out0;
wire  [11:0] v$RAMADDRMUX_14982_out0;
wire  [11:0] v$RAMADDRMUX_437_out0;
wire  [11:0] v$RAMADDRMUX_438_out0;
wire  [11:0] v$RAMADDRMUX_4959_out0;
wire  [11:0] v$RAMADDRMUX_4960_out0;
wire  [11:0] v$RAMADDRMUX_5029_out0;
wire  [11:0] v$RAMADDRMUX_5030_out0;
wire  [11:0] v$RAMADDR_14184_out0;
wire  [11:0] v$RAMADDR_19265_out0;
wire  [11:0] v$RAMADDR_9116_out0;
wire  [11:0] v$RAMAddress_2469_out0;
wire  [11:0] v$RAMAddress_2470_out0;
wire  [11:0] v$SEL1_12547_out0;
wire  [11:0] v$SEL1_12548_out0;
wire  [11:0] v$SEL1_3473_out0;
wire  [11:0] v$SEL1_3474_out0;
wire  [11:0] v$SEL2_14330_out0;
wire  [11:0] v$SEL2_14331_out0;
wire  [11:0] v$SEL3_1405_out0;
wire  [11:0] v$SEL3_1406_out0;
wire  [11:0] v$SEL4_1527_out0;
wire  [11:0] v$SEL4_1528_out0;
wire  [11:0] v$SUM_14246_out0;
wire  [11:0] v$SUM_14247_out0;
wire  [11:0] v$_14634_out0;
wire  [11:0] v$_14635_out0;
wire  [11:0] v$_15203_out0;
wire  [11:0] v$_15207_out0;
wire  [11:0] v$_15239_out0;
wire  [11:0] v$_15243_out0;
wire  [11:0] v$_16985_out0;
wire  [11:0] v$_16986_out0;
wire  [11:0] v$_17370_out0;
wire  [11:0] v$_17374_out0;
wire  [11:0] v$_4140_out0;
wire  [11:0] v$_4140_out1;
wire  [11:0] v$_4141_out0;
wire  [11:0] v$_4141_out1;
wire  [11:0] v$_4142_out0;
wire  [11:0] v$_4142_out1;
wire  [11:0] v$_4143_out0;
wire  [11:0] v$_4143_out1;
wire  [11:0] v$_4144_out0;
wire  [11:0] v$_4144_out1;
wire  [11:0] v$_4145_out0;
wire  [11:0] v$_4145_out1;
wire  [11:0] v$_5015_out0;
wire  [11:0] v$_5019_out0;
wire  [11:0] v$_7860_out0;
wire  [11:0] v$_7860_out1;
wire  [11:0] v$_7861_out0;
wire  [11:0] v$_7861_out1;
wire  [11:0] v$_7862_out0;
wire  [11:0] v$_7862_out1;
wire  [11:0] v$_7863_out0;
wire  [11:0] v$_7863_out1;
wire  [11:0] v$_7864_out0;
wire  [11:0] v$_7864_out1;
wire  [11:0] v$_7865_out0;
wire  [11:0] v$_7865_out1;
wire  [11:0] v$_8037_out0;
wire  [11:0] v$_8038_out0;
wire  [12:0] v$C10_9279_out0;
wire  [12:0] v$C10_9280_out0;
wire  [12:0] v$C4_2644_out0;
wire  [12:0] v$C4_2645_out0;
wire  [12:0] v$C6_1689_out0;
wire  [12:0] v$C6_1690_out0;
wire  [12:0] v$C7_6318_out0;
wire  [12:0] v$C7_6319_out0;
wire  [12:0] v$C8_8515_out0;
wire  [12:0] v$C8_8516_out0;
wire  [13:0] v$_15202_out0;
wire  [13:0] v$_15206_out0;
wire  [13:0] v$_15238_out0;
wire  [13:0] v$_15242_out0;
wire  [13:0] v$_17369_out0;
wire  [13:0] v$_17373_out0;
wire  [13:0] v$_5014_out0;
wire  [13:0] v$_5018_out0;
wire  [14:0] v$C2_18617_out0;
wire  [14:0] v$C2_18618_out0;
wire  [14:0] v$C4_8566_out0;
wire  [14:0] v$C4_8568_out0;
wire  [14:0] v$MUX2_14208_out0;
wire  [14:0] v$MUX2_14210_out0;
wire  [14:0] v$SEL2_6430_out0;
wire  [14:0] v$SEL2_6431_out0;
wire  [14:0] v$_11912_out0;
wire  [14:0] v$_11913_out0;
wire  [14:0] v$_15201_out0;
wire  [14:0] v$_15205_out0;
wire  [14:0] v$_15237_out0;
wire  [14:0] v$_15241_out0;
wire  [14:0] v$_15764_out0;
wire  [14:0] v$_15765_out0;
wire  [14:0] v$_16450_out0;
wire  [14:0] v$_16452_out0;
wire  [14:0] v$_17368_out0;
wire  [14:0] v$_17372_out0;
wire  [14:0] v$_5013_out0;
wire  [14:0] v$_5017_out0;
wire  [15:0] v$A$COMPARATOR$IN_1619_out0;
wire  [15:0] v$A$COMPARATOR$IN_1620_out0;
wire  [15:0] v$A$IN$MULTIPLIER_4232_out0;
wire  [15:0] v$A$IN$MULTIPLIER_4233_out0;
wire  [15:0] v$A$SAVED$PIPELINED_17144_out0;
wire  [15:0] v$A$SAVED$PIPELINED_17145_out0;
wire  [15:0] v$A$SAVED_10392_out0;
wire  [15:0] v$A$SAVED_10393_out0;
wire  [15:0] v$A$SAVED_15235_out0;
wire  [15:0] v$A$SAVED_15236_out0;
wire  [15:0] v$A$SAVED_3877_out0;
wire  [15:0] v$A$SAVED_3878_out0;
wire  [15:0] v$A$VIEW_16922_out0;
wire  [15:0] v$A$VIEW_16923_out0;
wire  [15:0] v$A1_14282_out0;
wire  [15:0] v$A1_14283_out0;
wire  [15:0] v$A1_6652_out0;
wire  [15:0] v$A1_6653_out0;
wire  [15:0] v$A1_9805_out0;
wire  [15:0] v$A1_9806_out0;
wire  [15:0] v$ADDEROUT_3704_out0;
wire  [15:0] v$ADDEROUT_3705_out0;
wire  [15:0] v$ALUOUT$LOADSTORE_19243_out0;
wire  [15:0] v$ALUOUT$LOADSTORE_19244_out0;
wire  [15:0] v$ALUOUT_10671_out0;
wire  [15:0] v$ALUOUT_10672_out0;
wire  [15:0] v$ALUOUT_17162_out0;
wire  [15:0] v$ALUOUT_17163_out0;
wire  [15:0] v$ALUOUT_18679_out0;
wire  [15:0] v$ALUOUT_18680_out0;
wire  [15:0] v$ALUOUT_6045_out0;
wire  [15:0] v$ALUOUT_6046_out0;
wire  [15:0] v$ALUOUT_7203_out0;
wire  [15:0] v$ALUOUT_7204_out0;
wire  [15:0] v$ANDOUT_7689_out0;
wire  [15:0] v$ANDOUT_7690_out0;
wire  [15:0] v$A_11554_out0;
wire  [15:0] v$A_11555_out0;
wire  [15:0] v$A_14399_out0;
wire  [15:0] v$A_14401_out0;
wire  [15:0] v$A_14403_out0;
wire  [15:0] v$A_14405_out0;
wire  [15:0] v$A_17040_out0;
wire  [15:0] v$A_17041_out0;
wire  [15:0] v$A_17640_out0;
wire  [15:0] v$A_17641_out0;
wire  [15:0] v$A_18897_out0;
wire  [15:0] v$A_18898_out0;
wire  [15:0] v$A_2497_out0;
wire  [15:0] v$A_2498_out0;
wire  [15:0] v$A_2743_out0;
wire  [15:0] v$A_2744_out0;
wire  [15:0] v$A_3465_out0;
wire  [15:0] v$A_3466_out0;
wire  [15:0] v$A_4354_out0;
wire  [15:0] v$A_4355_out0;
wire  [15:0] v$A_9044_out0;
wire  [15:0] v$A_9045_out0;
wire  [15:0] v$A_9779_out0;
wire  [15:0] v$A_9780_out0;
wire  [15:0] v$B$COMPARATOR$IN_18577_out0;
wire  [15:0] v$B$COMPARATOR$IN_18578_out0;
wire  [15:0] v$B$IN$MULTIPLIER_16058_out0;
wire  [15:0] v$B$IN$MULTIPLIER_16059_out0;
wire  [15:0] v$B$IN_12212_out0;
wire  [15:0] v$B$IN_12213_out0;
wire  [15:0] v$B$MERGE_17206_out0;
wire  [15:0] v$B$MERGE_17207_out0;
wire  [15:0] v$B$SAVED$PIPELINED_18338_out0;
wire  [15:0] v$B$SAVED$PIPELINED_18339_out0;
wire  [15:0] v$B$SAVED_4066_out0;
wire  [15:0] v$B$SAVED_4067_out0;
wire  [15:0] v$B$SAVED_4522_out0;
wire  [15:0] v$B$SAVED_4523_out0;
wire  [15:0] v$B$SAVED_4961_out0;
wire  [15:0] v$B$SAVED_4962_out0;
wire  [15:0] v$B_10432_out0;
wire  [15:0] v$B_10433_out0;
wire  [15:0] v$B_12288_out0;
wire  [15:0] v$B_12289_out0;
wire  [15:0] v$B_14677_out0;
wire  [15:0] v$B_14678_out0;
wire  [15:0] v$B_17646_out0;
wire  [15:0] v$B_17647_out0;
wire  [15:0] v$B_18356_out0;
wire  [15:0] v$B_18357_out0;
wire  [15:0] v$B_18591_out0;
wire  [15:0] v$B_18592_out0;
wire  [15:0] v$B_18707_out0;
wire  [15:0] v$B_18708_out0;
wire  [15:0] v$B_3590_out0;
wire  [15:0] v$B_3591_out0;
wire  [15:0] v$B_5038_out0;
wire  [15:0] v$B_5040_out0;
wire  [15:0] v$B_5042_out0;
wire  [15:0] v$B_5044_out0;
wire  [15:0] v$B_6781_out0;
wire  [15:0] v$B_6782_out0;
wire  [15:0] v$C10_6624_out0;
wire  [15:0] v$C10_6625_out0;
wire  [15:0] v$C1_16938_out0;
wire  [15:0] v$C1_16939_out0;
wire  [15:0] v$C1_18809_out0;
wire  [15:0] v$C1_18810_out0;
wire  [15:0] v$C1_6242_out0;
wire  [15:0] v$C1_6247_out0;
wire  [15:0] v$C1_6252_out0;
wire  [15:0] v$C1_6260_out0;
wire  [15:0] v$C1_6262_out0;
wire  [15:0] v$C1_6270_out0;
wire  [15:0] v$C1_6273_out0;
wire  [15:0] v$C1_6278_out0;
wire  [15:0] v$C1_6283_out0;
wire  [15:0] v$C1_6291_out0;
wire  [15:0] v$C1_6293_out0;
wire  [15:0] v$C1_6301_out0;
wire  [15:0] v$C2_10434_out0;
wire  [15:0] v$C2_10435_out0;
wire  [15:0] v$C2_104_out0;
wire  [15:0] v$C2_109_out0;
wire  [15:0] v$C2_114_out0;
wire  [15:0] v$C2_122_out0;
wire  [15:0] v$C2_124_out0;
wire  [15:0] v$C2_12772_out0;
wire  [15:0] v$C2_12773_out0;
wire  [15:0] v$C2_132_out0;
wire  [15:0] v$C2_135_out0;
wire  [15:0] v$C2_140_out0;
wire  [15:0] v$C2_145_out0;
wire  [15:0] v$C2_153_out0;
wire  [15:0] v$C2_155_out0;
wire  [15:0] v$C2_163_out0;
wire  [15:0] v$C3_12770_out0;
wire  [15:0] v$C3_12771_out0;
wire  [15:0] v$C7_1867_out0;
wire  [15:0] v$C7_1868_out0;
wire  [15:0] v$C9_19371_out0;
wire  [15:0] v$C9_19372_out0;
wire  [15:0] v$C9_3525_out0;
wire  [15:0] v$C9_3526_out0;
wire  [15:0] v$COUNTERTHRESHOLD_18563_out0;
wire  [15:0] v$COUNTERTHRESHOLD_18564_out0;
wire  [15:0] v$COUNTERVALUE_3197_out0;
wire  [15:0] v$COUNTERVALUE_3198_out0;
wire  [15:0] v$C_18715_out0;
wire  [15:0] v$C_18716_out0;
wire  [15:0] v$DATA$IN0_10855_out0;
wire  [15:0] v$DATA$IN1_15866_out0;
wire  [15:0] v$DATA$IN_1763_out0;
wire  [15:0] v$DATA$IN_1764_out0;
wire  [15:0] v$DATA$IN_7364_out0;
wire  [15:0] v$DATA$IN_7365_out0;
wire  [15:0] v$DATA$OUT0_12867_out0;
wire  [15:0] v$DATA$OUT1_16195_out0;
wire  [15:0] v$DATA$OUT_1468_out0;
wire  [15:0] v$DATA$OUT_1469_out0;
wire  [15:0] v$DATA$OUT_7936_out0;
wire  [15:0] v$DATA$OUT_7937_out0;
wire  [15:0] v$DATAIN0_11570_out0;
wire  [15:0] v$DATAIN1_10016_out0;
wire  [15:0] v$DATAINCP_11498_out0;
wire  [15:0] v$DATAINCP_11499_out0;
wire  [15:0] v$DATA_14697_out0;
wire  [15:0] v$DATA_14698_out0;
wire  [15:0] v$DATA_4518_out0;
wire  [15:0] v$DATA_4519_out0;
wire  [15:0] v$DIN$FIRST$MUX_7812_out0;
wire  [15:0] v$DIN$FIRST$MUX_7813_out0;
wire  [15:0] v$DIN3$VIEWER_2412_out0;
wire  [15:0] v$DIN3$VIEWER_2413_out0;
wire  [15:0] v$DIN3_15022_out0;
wire  [15:0] v$DIN3_15023_out0;
wire  [15:0] v$DIN_1883_out0;
wire  [15:0] v$DIN_1884_out0;
wire  [15:0] v$DIN_1965_out0;
wire  [15:0] v$DIN_1966_out0;
wire  [15:0] v$DM1_8182_out0;
wire  [15:0] v$DM1_8182_out1;
wire  [15:0] v$DOUT1_3375_out0;
wire  [15:0] v$DOUT1_3376_out0;
wire  [15:0] v$DOUT2_3714_out0;
wire  [15:0] v$DOUT2_3715_out0;
wire  [15:0] v$FPU$A_16484_out0;
wire  [15:0] v$FPU$A_16485_out0;
wire  [15:0] v$FPU$B$EN_7295_out0;
wire  [15:0] v$FPU$B$EN_7296_out0;
wire  [15:0] v$FPU$OUT_17605_out0;
wire  [15:0] v$FPU$OUT_17606_out0;
wire  [15:0] v$FPU$OUT_8053_out0;
wire  [15:0] v$FPU$OUT_8054_out0;
wire  [15:0] v$HAZ$DECTECTOR$A_18565_out0;
wire  [15:0] v$HAZ$DECTECTOR$A_18566_out0;
wire  [15:0] v$HAZ$DETECTOR$B_5289_out0;
wire  [15:0] v$HAZ$DETECTOR$B_5290_out0;
wire  [15:0] v$INSTR$READ0_14785_out0;
wire  [15:0] v$INSTR$READ1_12546_out0;
wire  [15:0] v$INSTR$READ_15505_out0;
wire  [15:0] v$INSTR$READ_15506_out0;
wire  [15:0] v$INSTR$READ_7535_out0;
wire  [15:0] v$INSTR$READ_7536_out0;
wire  [15:0] v$IN_14141_out0;
wire  [15:0] v$IN_14143_out0;
wire  [15:0] v$IN_14145_out0;
wire  [15:0] v$IN_14147_out0;
wire  [15:0] v$IN_196_out0;
wire  [15:0] v$IN_197_out0;
wire  [15:0] v$IN_4524_out0;
wire  [15:0] v$IN_4525_out0;
wire  [15:0] v$IN_4526_out0;
wire  [15:0] v$IN_4527_out0;
wire  [15:0] v$IN_4528_out0;
wire  [15:0] v$IN_4529_out0;
wire  [15:0] v$IN_4530_out0;
wire  [15:0] v$IN_4531_out0;
wire  [15:0] v$IN_9946_out0;
wire  [15:0] v$IN_9947_out0;
wire  [15:0] v$IN_9948_out0;
wire  [15:0] v$IN_9949_out0;
wire  [15:0] v$IN_9950_out0;
wire  [15:0] v$IN_9951_out0;
wire  [15:0] v$IN_9952_out0;
wire  [15:0] v$IN_9953_out0;
wire  [15:0] v$IR$READ$IN$PREV$CYCLE_6449_out0;
wire  [15:0] v$IR$READ$IN$PREV$CYCLE_6450_out0;
wire  [15:0] v$IR1$VIEWER_7746_out0;
wire  [15:0] v$IR1$VIEWER_7747_out0;
wire  [15:0] v$IR1_13974_out0;
wire  [15:0] v$IR1_13975_out0;
wire  [15:0] v$IR1_16608_out0;
wire  [15:0] v$IR1_16609_out0;
wire  [15:0] v$IR1_17302_out0;
wire  [15:0] v$IR1_17303_out0;
wire  [15:0] v$IR1_18639_out0;
wire  [15:0] v$IR1_18640_out0;
wire  [15:0] v$IR1_22_out0;
wire  [15:0] v$IR1_23_out0;
wire  [15:0] v$IR1_4315_out0;
wire  [15:0] v$IR1_4316_out0;
wire  [15:0] v$IR1_706_out0;
wire  [15:0] v$IR1_707_out0;
wire  [15:0] v$IR1_7941_out0;
wire  [15:0] v$IR1_7942_out0;
wire  [15:0] v$IR2$VIEWER_16914_out0;
wire  [15:0] v$IR2$VIEWER_16915_out0;
wire  [15:0] v$IR2_17178_out0;
wire  [15:0] v$IR2_17179_out0;
wire  [15:0] v$IR2_18567_out0;
wire  [15:0] v$IR2_18568_out0;
wire  [15:0] v$IR2_1911_out0;
wire  [15:0] v$IR2_1912_out0;
wire  [15:0] v$IR2_2422_out0;
wire  [15:0] v$IR2_2423_out0;
wire  [15:0] v$IR2_3141_out0;
wire  [15:0] v$IR2_3142_out0;
wire  [15:0] v$IR2_3511_out0;
wire  [15:0] v$IR2_3512_out0;
wire  [15:0] v$IR2_4118_out0;
wire  [15:0] v$IR2_4119_out0;
wire  [15:0] v$IR2_8094_out0;
wire  [15:0] v$IR2_8095_out0;
wire  [15:0] v$LDST$RAMDOUT_1305_out0;
wire  [15:0] v$LDST$RAMDOUT_1306_out0;
wire  [15:0] v$LDST$RMN_8045_out0;
wire  [15:0] v$LDST$RMN_8046_out0;
wire  [15:0] v$LDSTN_3253_out0;
wire  [15:0] v$LDSTN_3254_out0;
wire  [15:0] v$LDSTRM_7973_out0;
wire  [15:0] v$LDSTRM_7974_out0;
wire  [15:0] v$LOAD$STORE$OUT_18198_out0;
wire  [15:0] v$LOAD$STORE$OUT_18199_out0;
wire  [15:0] v$LOWER$PART_7796_out0;
wire  [15:0] v$LOWER$PART_7797_out0;
wire  [15:0] v$MULTIPLY$DENORMALIZATION$16$BIT_12284_out0;
wire  [15:0] v$MULTIPLY$DENORMALIZATION$16$BIT_12285_out0;
wire  [15:0] v$MUX10_17440_out0;
wire  [15:0] v$MUX10_17441_out0;
wire  [15:0] v$MUX11_9016_out0;
wire  [15:0] v$MUX11_9017_out0;
wire  [15:0] v$MUX13_2745_out0;
wire  [15:0] v$MUX13_2746_out0;
wire  [15:0] v$MUX14_19331_out0;
wire  [15:0] v$MUX14_19332_out0;
wire  [15:0] v$MUX15_7291_out0;
wire  [15:0] v$MUX15_7292_out0;
wire  [15:0] v$MUX16_19139_out0;
wire  [15:0] v$MUX16_19140_out0;
wire  [15:0] v$MUX1_12320_out0;
wire  [15:0] v$MUX1_12321_out0;
wire  [15:0] v$MUX1_15845_out0;
wire  [15:0] v$MUX1_15846_out0;
wire  [15:0] v$MUX1_18336_out0;
wire  [15:0] v$MUX1_18337_out0;
wire  [15:0] v$MUX1_18934_out0;
wire  [15:0] v$MUX1_18935_out0;
wire  [15:0] v$MUX1_1973_out0;
wire  [15:0] v$MUX1_1974_out0;
wire  [15:0] v$MUX1_2159_out0;
wire  [15:0] v$MUX1_2160_out0;
wire  [15:0] v$MUX1_2798_out0;
wire  [15:0] v$MUX1_2799_out0;
wire  [15:0] v$MUX1_4198_out0;
wire  [15:0] v$MUX1_4199_out0;
wire  [15:0] v$MUX1_6106_out0;
wire  [15:0] v$MUX1_6107_out0;
wire  [15:0] v$MUX1_6914_out0;
wire  [15:0] v$MUX1_6915_out0;
wire  [15:0] v$MUX1_6916_out0;
wire  [15:0] v$MUX1_6917_out0;
wire  [15:0] v$MUX1_6918_out0;
wire  [15:0] v$MUX1_6919_out0;
wire  [15:0] v$MUX1_6920_out0;
wire  [15:0] v$MUX1_6921_out0;
wire  [15:0] v$MUX2_11162_out0;
wire  [15:0] v$MUX2_11163_out0;
wire  [15:0] v$MUX2_12557_out0;
wire  [15:0] v$MUX2_12558_out0;
wire  [15:0] v$MUX2_12603_out0;
wire  [15:0] v$MUX2_12604_out0;
wire  [15:0] v$MUX2_12605_out0;
wire  [15:0] v$MUX2_12606_out0;
wire  [15:0] v$MUX2_12607_out0;
wire  [15:0] v$MUX2_12608_out0;
wire  [15:0] v$MUX2_12609_out0;
wire  [15:0] v$MUX2_12610_out0;
wire  [15:0] v$MUX2_15790_out0;
wire  [15:0] v$MUX2_15791_out0;
wire  [15:0] v$MUX2_16447_out0;
wire  [15:0] v$MUX3_1741_out0;
wire  [15:0] v$MUX3_1742_out0;
wire  [15:0] v$MUX3_18992_out0;
wire  [15:0] v$MUX3_18993_out0;
wire  [15:0] v$MUX3_2122_out0;
wire  [15:0] v$MUX3_2123_out0;
wire  [15:0] v$MUX3_2124_out0;
wire  [15:0] v$MUX3_2125_out0;
wire  [15:0] v$MUX3_2126_out0;
wire  [15:0] v$MUX3_2127_out0;
wire  [15:0] v$MUX3_2128_out0;
wire  [15:0] v$MUX3_2129_out0;
wire  [15:0] v$MUX3_4062_out0;
wire  [15:0] v$MUX3_4063_out0;
wire  [15:0] v$MUX4_16600_out0;
wire  [15:0] v$MUX4_16601_out0;
wire  [15:0] v$MUX4_16602_out0;
wire  [15:0] v$MUX4_16603_out0;
wire  [15:0] v$MUX4_16604_out0;
wire  [15:0] v$MUX4_16605_out0;
wire  [15:0] v$MUX4_16606_out0;
wire  [15:0] v$MUX4_16607_out0;
wire  [15:0] v$MUX4_1809_out0;
wire  [15:0] v$MUX4_1810_out0;
wire  [15:0] v$MUX4_18328_out0;
wire  [15:0] v$MUX4_18329_out0;
wire  [15:0] v$MUX4_4023_out0;
wire  [15:0] v$MUX4_46_out0;
wire  [15:0] v$MUX4_47_out0;
wire  [15:0] v$MUX4_6214_out0;
wire  [15:0] v$MUX4_6215_out0;
wire  [15:0] v$MUX5_11398_out0;
wire  [15:0] v$MUX5_12517_out0;
wire  [15:0] v$MUX5_12518_out0;
wire  [15:0] v$MUX5_14693_out0;
wire  [15:0] v$MUX5_14694_out0;
wire  [15:0] v$MUX6_5267_out0;
wire  [15:0] v$MUX6_5268_out0;
wire  [15:0] v$MUX6_7758_out0;
wire  [15:0] v$MUX6_7759_out0;
wire  [15:0] v$MUX9_18555_out0;
wire  [15:0] v$MUX9_18556_out0;
wire  [15:0] v$NEXTENDED_14977_out0;
wire  [15:0] v$NEXTENDED_14978_out0;
wire  [15:0] v$NEXTENDED_2072_out0;
wire  [15:0] v$NEXTENDED_2073_out0;
wire  [15:0] v$OP1_15807_out0;
wire  [15:0] v$OP1_15808_out0;
wire  [15:0] v$OP1_5658_out0;
wire  [15:0] v$OP1_5659_out0;
wire  [15:0] v$OP2_10643_out0;
wire  [15:0] v$OP2_10644_out0;
wire  [15:0] v$OP2_14603_out0;
wire  [15:0] v$OP2_14604_out0;
wire  [15:0] v$OP2_15675_out0;
wire  [15:0] v$OP2_15676_out0;
wire  [15:0] v$OP2_7906_out0;
wire  [15:0] v$OP2_7907_out0;
wire  [15:0] v$OUT_13072_out0;
wire  [15:0] v$OUT_13074_out0;
wire  [15:0] v$OUT_1483_out0;
wire  [15:0] v$OUT_1484_out0;
wire  [15:0] v$OUT_15104_out0;
wire  [15:0] v$OUT_15105_out0;
wire  [15:0] v$OUT_3397_out0;
wire  [15:0] v$OUT_3398_out0;
wire  [15:0] v$OUT_3399_out0;
wire  [15:0] v$OUT_3400_out0;
wire  [15:0] v$OUT_3401_out0;
wire  [15:0] v$OUT_3402_out0;
wire  [15:0] v$OUT_3403_out0;
wire  [15:0] v$OUT_3404_out0;
wire  [15:0] v$OUT_5477_out0;
wire  [15:0] v$OUT_8651_out0;
wire  [15:0] v$PIN_3143_out0;
wire  [15:0] v$PIN_3144_out0;
wire  [15:0] v$R0TEST_14651_out0;
wire  [15:0] v$R0TEST_14652_out0;
wire  [15:0] v$R0TEST_8545_out0;
wire  [15:0] v$R0TEST_8546_out0;
wire  [15:0] v$R0_3503_out0;
wire  [15:0] v$R0_3504_out0;
wire  [15:0] v$R1TEST_15756_out0;
wire  [15:0] v$R1TEST_15757_out0;
wire  [15:0] v$R1TEST_8559_out0;
wire  [15:0] v$R1TEST_8560_out0;
wire  [15:0] v$R1_14351_out0;
wire  [15:0] v$R1_14352_out0;
wire  [15:0] v$R2TEST_16315_out0;
wire  [15:0] v$R2TEST_16316_out0;
wire  [15:0] v$R2TEST_16409_out0;
wire  [15:0] v$R2TEST_16410_out0;
wire  [15:0] v$R2_8285_out0;
wire  [15:0] v$R2_8286_out0;
wire  [15:0] v$R3TEST_12376_out0;
wire  [15:0] v$R3TEST_12377_out0;
wire  [15:0] v$R3TEST_7858_out0;
wire  [15:0] v$R3TEST_7859_out0;
wire  [15:0] v$R3_11234_out0;
wire  [15:0] v$R3_11235_out0;
wire  [15:0] v$RAM1_13483_out0;
wire  [15:0] v$RAMDIN_7323_out0;
wire  [15:0] v$RAMDIN_7324_out0;
wire  [15:0] v$RAMDOUT$DATAPATH_702_out0;
wire  [15:0] v$RAMDOUT$DATAPATH_703_out0;
wire  [15:0] v$RAMDOUT0_9426_out0;
wire  [15:0] v$RAMDOUT1_8627_out0;
wire  [15:0] v$RAMDOUT_17399_out0;
wire  [15:0] v$RAMDOUT_17400_out0;
wire  [15:0] v$RAMDOUT_5664_out0;
wire  [15:0] v$RAMDOUT_5665_out0;
wire  [15:0] v$RAMDOUT_68_out0;
wire  [15:0] v$RAMDOUT_69_out0;
wire  [15:0] v$RAMDOUT_8245_out0;
wire  [15:0] v$RAMDOUT_8246_out0;
wire  [15:0] v$RAMDOutOut_3407_out0;
wire  [15:0] v$RAMDOutOut_3408_out0;
wire  [15:0] v$RDOUT_10807_out0;
wire  [15:0] v$RDOUT_10808_out0;
wire  [15:0] v$RD_2432_out0;
wire  [15:0] v$RD_2433_out0;
wire  [15:0] v$REGDIN_17124_out0;
wire  [15:0] v$REGDIN_17125_out0;
wire  [15:0] v$REGDIN_18984_out0;
wire  [15:0] v$REGDIN_18985_out0;
wire  [15:0] v$RMN_6420_out0;
wire  [15:0] v$RMN_6421_out0;
wire  [15:0] v$RMORIGINAL_13550_out0;
wire  [15:0] v$RMORIGINAL_13551_out0;
wire  [15:0] v$RM_10695_out0;
wire  [15:0] v$RM_10696_out0;
wire  [15:0] v$RM_16803_out0;
wire  [15:0] v$RM_16804_out0;
wire  [15:0] v$RM_18797_out0;
wire  [15:0] v$RM_18798_out0;
wire  [15:0] v$RM_19205_out0;
wire  [15:0] v$RM_19206_out0;
wire  [15:0] v$RM_9801_out0;
wire  [15:0] v$RM_9802_out0;
wire  [15:0] v$ROM1_3190_out0;
wire  [15:0] v$ROM1_7586_out0;
wire  [15:0] v$R_18958_out0;
wire  [15:0] v$R_18959_out0;
wire  [15:0] v$R_60_out0;
wire  [15:0] v$R_61_out0;
wire  [15:0] v$SEL11_3883_out0;
wire  [15:0] v$SEL11_3884_out0;
wire  [15:0] v$SEL12_1339_out0;
wire  [15:0] v$SEL12_1340_out0;
wire  [15:0] v$SEL1_15975_out0;
wire  [15:0] v$SEL1_15980_out0;
wire  [15:0] v$SEL1_15985_out0;
wire  [15:0] v$SEL1_15990_out0;
wire  [15:0] v$SEL1_15995_out0;
wire  [15:0] v$SEL1_16000_out0;
wire  [15:0] v$SEL1_16006_out0;
wire  [15:0] v$SEL1_16011_out0;
wire  [15:0] v$SEL1_16016_out0;
wire  [15:0] v$SEL1_16021_out0;
wire  [15:0] v$SEL1_16026_out0;
wire  [15:0] v$SEL1_16031_out0;
wire  [15:0] v$SEL1_9047_out0;
wire  [15:0] v$SEL1_9052_out0;
wire  [15:0] v$SEL1_9057_out0;
wire  [15:0] v$SEL1_9062_out0;
wire  [15:0] v$SEL1_9067_out0;
wire  [15:0] v$SEL1_9072_out0;
wire  [15:0] v$SEL1_9078_out0;
wire  [15:0] v$SEL1_9083_out0;
wire  [15:0] v$SEL1_9088_out0;
wire  [15:0] v$SEL1_9093_out0;
wire  [15:0] v$SEL1_9098_out0;
wire  [15:0] v$SEL1_9103_out0;
wire  [15:0] v$SEL2_6634_out0;
wire  [15:0] v$SEL2_6635_out0;
wire  [15:0] v$SEL2_6636_out0;
wire  [15:0] v$SEL2_6637_out0;
wire  [15:0] v$SEL4_9936_out0;
wire  [15:0] v$SEL4_9937_out0;
wire  [15:0] v$SEL5_14164_out0;
wire  [15:0] v$SEL5_14165_out0;
wire  [15:0] v$SHIFT1OUT_7908_out0;
wire  [15:0] v$SHIFT1OUT_7909_out0;
wire  [15:0] v$SHIFT2OUT_16274_out0;
wire  [15:0] v$SHIFT2OUT_16275_out0;
wire  [15:0] v$SHIFT4OUT_6222_out0;
wire  [15:0] v$SHIFT4OUT_6223_out0;
wire  [15:0] v$SHIFT8OUT_8329_out0;
wire  [15:0] v$SHIFT8OUT_8330_out0;
wire  [15:0] v$SUM_10759_out0;
wire  [15:0] v$SUM_10760_out0;
wire  [15:0] v$THRESHOLD_16123_out0;
wire  [15:0] v$THRESHOLD_16124_out0;
wire  [15:0] v$UART$DOUT_18104_out0;
wire  [15:0] v$UART$DOUT_18105_out0;
wire  [15:0] v$XOR1_5297_out0;
wire  [15:0] v$XOR1_5298_out0;
wire  [15:0] v$XOR1_9920_out0;
wire  [15:0] v$XOR1_9921_out0;
wire  [15:0] v$_10354_out1;
wire  [15:0] v$_10355_out1;
wire  [15:0] v$_12208_out0;
wire  [15:0] v$_12209_out0;
wire  [15:0] v$_12326_out0;
wire  [15:0] v$_12327_out0;
wire  [15:0] v$_12380_out0;
wire  [15:0] v$_12381_out0;
wire  [15:0] v$_12382_out0;
wire  [15:0] v$_12383_out0;
wire  [15:0] v$_12384_out0;
wire  [15:0] v$_12385_out0;
wire  [15:0] v$_12386_out0;
wire  [15:0] v$_12387_out0;
wire  [15:0] v$_12795_out0;
wire  [15:0] v$_12796_out0;
wire  [15:0] v$_13890_out0;
wire  [15:0] v$_13891_out0;
wire  [15:0] v$_13892_out0;
wire  [15:0] v$_13893_out0;
wire  [15:0] v$_13894_out0;
wire  [15:0] v$_13895_out0;
wire  [15:0] v$_13896_out0;
wire  [15:0] v$_13897_out0;
wire  [15:0] v$_1629_out0;
wire  [15:0] v$_1630_out0;
wire  [15:0] v$_1631_out0;
wire  [15:0] v$_1632_out0;
wire  [15:0] v$_1633_out0;
wire  [15:0] v$_1634_out0;
wire  [15:0] v$_1635_out0;
wire  [15:0] v$_1636_out0;
wire  [15:0] v$_1649_out0;
wire  [15:0] v$_1650_out0;
wire  [15:0] v$_16985_out1;
wire  [15:0] v$_16986_out1;
wire  [15:0] v$_16987_out0;
wire  [15:0] v$_16988_out0;
wire  [15:0] v$_18118_out0;
wire  [15:0] v$_18119_out0;
wire  [15:0] v$_18834_out0;
wire  [15:0] v$_18835_out0;
wire  [15:0] v$_18836_out0;
wire  [15:0] v$_18837_out0;
wire  [15:0] v$_18838_out0;
wire  [15:0] v$_18839_out0;
wire  [15:0] v$_19023_out0;
wire  [15:0] v$_19025_out0;
wire  [15:0] v$_5082_out0;
wire  [15:0] v$_5083_out0;
wire  [15:0] v$_5084_out0;
wire  [15:0] v$_5085_out0;
wire  [15:0] v$_5086_out0;
wire  [15:0] v$_5087_out0;
wire  [15:0] v$_7193_out0;
wire  [15:0] v$_7194_out0;
wire  [15:0] v$_9819_out0;
wire  [15:0] v$_9820_out0;
wire  [15:0] v$_9821_out0;
wire  [15:0] v$_9822_out0;
wire  [15:0] v$_9823_out0;
wire  [15:0] v$_9824_out0;
wire  [15:0] v$_9825_out0;
wire  [15:0] v$_9826_out0;
wire  [19:0] v$SEL1_15977_out0;
wire  [19:0] v$SEL1_15982_out0;
wire  [19:0] v$SEL1_15987_out0;
wire  [19:0] v$SEL1_15991_out0;
wire  [19:0] v$SEL1_15997_out0;
wire  [19:0] v$SEL1_16001_out0;
wire  [19:0] v$SEL1_16008_out0;
wire  [19:0] v$SEL1_16013_out0;
wire  [19:0] v$SEL1_16018_out0;
wire  [19:0] v$SEL1_16022_out0;
wire  [19:0] v$SEL1_16028_out0;
wire  [19:0] v$SEL1_16032_out0;
wire  [19:0] v$SEL1_9049_out0;
wire  [19:0] v$SEL1_9054_out0;
wire  [19:0] v$SEL1_9059_out0;
wire  [19:0] v$SEL1_9063_out0;
wire  [19:0] v$SEL1_9069_out0;
wire  [19:0] v$SEL1_9073_out0;
wire  [19:0] v$SEL1_9080_out0;
wire  [19:0] v$SEL1_9085_out0;
wire  [19:0] v$SEL1_9090_out0;
wire  [19:0] v$SEL1_9094_out0;
wire  [19:0] v$SEL1_9100_out0;
wire  [19:0] v$SEL1_9104_out0;
wire  [1:0] v$2_13308_out0;
wire  [1:0] v$2_13309_out0;
wire  [1:0] v$5_7828_out0;
wire  [1:0] v$5_7829_out0;
wire  [1:0] v$7_14618_out0;
wire  [1:0] v$7_14619_out0;
wire  [1:0] v$8_1341_out0;
wire  [1:0] v$8_1342_out0;
wire  [1:0] v$AD1VIEWER_7293_out0;
wire  [1:0] v$AD1VIEWER_7294_out0;
wire  [1:0] v$AD1_19284_out0;
wire  [1:0] v$AD1_19285_out0;
wire  [1:0] v$AD1_2001_out0;
wire  [1:0] v$AD1_2002_out0;
wire  [1:0] v$AD1_6891_out0;
wire  [1:0] v$AD1_6892_out0;
wire  [1:0] v$AD1_7932_out0;
wire  [1:0] v$AD1_7933_out0;
wire  [1:0] v$AD2$viewer_16349_out0;
wire  [1:0] v$AD2$viewer_16350_out0;
wire  [1:0] v$AD2_16254_out0;
wire  [1:0] v$AD2_16255_out0;
wire  [1:0] v$AD2_4108_out0;
wire  [1:0] v$AD2_4109_out0;
wire  [1:0] v$AD2_6644_out0;
wire  [1:0] v$AD2_6645_out0;
wire  [1:0] v$AD2_9422_out0;
wire  [1:0] v$AD2_9423_out0;
wire  [1:0] v$AD3$VIEWER_8630_out0;
wire  [1:0] v$AD3$VIEWER_8631_out0;
wire  [1:0] v$AD3_13721_out0;
wire  [1:0] v$AD3_13722_out0;
wire  [1:0] v$AD3_15754_out0;
wire  [1:0] v$AD3_15755_out0;
wire  [1:0] v$C1_14855_out0;
wire  [1:0] v$C1_14856_out0;
wire  [1:0] v$C1_3229_out0;
wire  [1:0] v$C1_3230_out0;
wire  [1:0] v$C1_6246_out0;
wire  [1:0] v$C1_6251_out0;
wire  [1:0] v$C1_6256_out0;
wire  [1:0] v$C1_6261_out0;
wire  [1:0] v$C1_6266_out0;
wire  [1:0] v$C1_6271_out0;
wire  [1:0] v$C1_6277_out0;
wire  [1:0] v$C1_6282_out0;
wire  [1:0] v$C1_6287_out0;
wire  [1:0] v$C1_6292_out0;
wire  [1:0] v$C1_6297_out0;
wire  [1:0] v$C1_6302_out0;
wire  [1:0] v$C1_8041_out0;
wire  [1:0] v$C1_8042_out0;
wire  [1:0] v$C1_8288_out0;
wire  [1:0] v$C1_8292_out0;
wire  [1:0] v$C2_108_out0;
wire  [1:0] v$C2_113_out0;
wire  [1:0] v$C2_118_out0;
wire  [1:0] v$C2_123_out0;
wire  [1:0] v$C2_128_out0;
wire  [1:0] v$C2_133_out0;
wire  [1:0] v$C2_13971_out0;
wire  [1:0] v$C2_13972_out0;
wire  [1:0] v$C2_139_out0;
wire  [1:0] v$C2_144_out0;
wire  [1:0] v$C2_149_out0;
wire  [1:0] v$C2_154_out0;
wire  [1:0] v$C2_159_out0;
wire  [1:0] v$C2_164_out0;
wire  [1:0] v$C3_3527_out0;
wire  [1:0] v$C3_3528_out0;
wire  [1:0] v$C3_3529_out0;
wire  [1:0] v$C3_3530_out0;
wire  [1:0] v$C4_16916_out0;
wire  [1:0] v$C4_16917_out0;
wire  [1:0] v$C4_17134_out0;
wire  [1:0] v$C4_17135_out0;
wire  [1:0] v$C4_17136_out0;
wire  [1:0] v$C4_17137_out0;
wire  [1:0] v$C5_17520_out0;
wire  [1:0] v$C5_17522_out0;
wire  [1:0] v$C5_17524_out0;
wire  [1:0] v$C5_17526_out0;
wire  [1:0] v$C6_6771_out0;
wire  [1:0] v$C6_6772_out0;
wire  [1:0] v$C6_6773_out0;
wire  [1:0] v$C6_6774_out0;
wire  [1:0] v$C6_6775_out0;
wire  [1:0] v$C6_6776_out0;
wire  [1:0] v$C6_6777_out0;
wire  [1:0] v$C6_6778_out0;
wire  [1:0] v$END_12506_out0;
wire  [1:0] v$END_12724_out0;
wire  [1:0] v$END_407_out0;
wire  [1:0] v$END_408_out0;
wire  [1:0] v$FPU$OP_13331_out0;
wire  [1:0] v$FPU$OP_13332_out0;
wire  [1:0] v$FPU$OP_14679_out0;
wire  [1:0] v$FPU$OP_14680_out0;
wire  [1:0] v$FPU$OP_16334_out0;
wire  [1:0] v$FPU$OP_16335_out0;
wire  [1:0] v$INTERRUPTNUMBER_40_out0;
wire  [1:0] v$INTERRUPTNUMBER_41_out0;
wire  [1:0] v$IR1$D_15458_out0;
wire  [1:0] v$IR1$D_15459_out0;
wire  [1:0] v$IR1$D_4378_out0;
wire  [1:0] v$IR1$D_4379_out0;
wire  [1:0] v$IR1$FPU$OP$CODE_18922_out0;
wire  [1:0] v$IR1$FPU$OP$CODE_18923_out0;
wire  [1:0] v$IR1$FPU$OP_4019_out0;
wire  [1:0] v$IR1$FPU$OP_4020_out0;
wire  [1:0] v$IR1$M_13215_out0;
wire  [1:0] v$IR1$M_13216_out0;
wire  [1:0] v$IR1$M_13829_out0;
wire  [1:0] v$IR1$M_13830_out0;
wire  [1:0] v$IR1$RD$VIEWER_18976_out0;
wire  [1:0] v$IR1$RD$VIEWER_18977_out0;
wire  [1:0] v$IR1$RD_5731_out0;
wire  [1:0] v$IR1$RD_5732_out0;
wire  [1:0] v$IR1$RM$VIEWER_8237_out0;
wire  [1:0] v$IR1$RM$VIEWER_8238_out0;
wire  [1:0] v$IR1$RM_18905_out0;
wire  [1:0] v$IR1$RM_18906_out0;
wire  [1:0] v$IR1$RM_18_out0;
wire  [1:0] v$IR1$RM_19_out0;
wire  [1:0] v$IR2$D_15090_out0;
wire  [1:0] v$IR2$D_15091_out0;
wire  [1:0] v$IR2$D_5114_out0;
wire  [1:0] v$IR2$D_5115_out0;
wire  [1:0] v$IR2$FPU$OP_1845_out0;
wire  [1:0] v$IR2$FPU$OP_1846_out0;
wire  [1:0] v$IR2$FPU$OP_3088_out0;
wire  [1:0] v$IR2$FPU$OP_3089_out0;
wire  [1:0] v$IR2$FPU$OP_7868_out0;
wire  [1:0] v$IR2$FPU$OP_7869_out0;
wire  [1:0] v$IR2$M_13567_out0;
wire  [1:0] v$IR2$M_13568_out0;
wire  [1:0] v$IR2$M_9178_out0;
wire  [1:0] v$IR2$M_9179_out0;
wire  [1:0] v$IR2$RD$VIEWER_9452_out0;
wire  [1:0] v$IR2$RD$VIEWER_9453_out0;
wire  [1:0] v$IR2$RD_13875_out0;
wire  [1:0] v$IR2$RD_13876_out0;
wire  [1:0] v$IR2$RD_16976_out0;
wire  [1:0] v$IR2$RD_16977_out0;
wire  [1:0] v$MUX10_3816_out0;
wire  [1:0] v$MUX10_3817_out0;
wire  [1:0] v$MUX11_4657_out0;
wire  [1:0] v$MUX11_4658_out0;
wire  [1:0] v$MUX16_9038_out0;
wire  [1:0] v$MUX16_9039_out0;
wire  [1:0] v$MUX1_8649_out0;
wire  [1:0] v$MUX1_8650_out0;
wire  [1:0] v$MUX2_3090_out0;
wire  [1:0] v$MUX2_3091_out0;
wire  [1:0] v$MUX5_8281_out0;
wire  [1:0] v$MUX5_8282_out0;
wire  [1:0] v$MUX6_1472_out0;
wire  [1:0] v$MUX6_1473_out0;
wire  [1:0] v$MUX9_7977_out0;
wire  [1:0] v$MUX9_7978_out0;
wire  [1:0] v$NINTERRUPT_1752_out0;
wire  [1:0] v$NINTERRUPT_1753_out0;
wire  [1:0] v$NINT_3070_out0;
wire  [1:0] v$NINT_3071_out0;
wire  [1:0] v$OP_1485_out0;
wire  [1:0] v$OP_1486_out0;
wire  [1:0] v$RD$FPU_13518_out0;
wire  [1:0] v$RD$FPU_13519_out0;
wire  [1:0] v$RD$OUT_18500_out0;
wire  [1:0] v$RD$OUT_18501_out0;
wire  [1:0] v$RD_12364_out0;
wire  [1:0] v$RD_12365_out0;
wire  [1:0] v$S$REG_3653_out0;
wire  [1:0] v$S$REG_3654_out0;
wire  [1:0] v$SEL10_13393_out0;
wire  [1:0] v$SEL10_13394_out0;
wire  [1:0] v$SEL13_5054_out0;
wire  [1:0] v$SEL13_5055_out0;
wire  [1:0] v$SEL1_5457_out0;
wire  [1:0] v$SEL1_5458_out0;
wire  [1:0] v$SEL4_9817_out0;
wire  [1:0] v$SEL4_9818_out0;
wire  [1:0] v$SEL5_704_out0;
wire  [1:0] v$SEL5_705_out0;
wire  [1:0] v$SEL6_3219_out0;
wire  [1:0] v$SEL6_3220_out0;
wire  [1:0] v$SEL8_15723_out0;
wire  [1:0] v$SEL8_15724_out0;
wire  [1:0] v$SEL9_8299_out0;
wire  [1:0] v$SEL9_8300_out0;
wire  [1:0] v$SHIFT_7303_out0;
wire  [1:0] v$SHIFT_7304_out0;
wire  [1:0] v$SHIFT_8348_out0;
wire  [1:0] v$SHIFT_8349_out0;
wire  [1:0] v$SR_10350_out0;
wire  [1:0] v$SR_10351_out0;
wire  [1:0] v$SR_17424_out0;
wire  [1:0] v$SR_17425_out0;
wire  [1:0] v$SR_17426_out0;
wire  [1:0] v$SR_17427_out0;
wire  [1:0] v$SR_17428_out0;
wire  [1:0] v$SR_17429_out0;
wire  [1:0] v$SR_17430_out0;
wire  [1:0] v$SR_17431_out0;
wire  [1:0] v$SR_4532_out0;
wire  [1:0] v$SR_4533_out0;
wire  [1:0] v$SR_4534_out0;
wire  [1:0] v$SR_4535_out0;
wire  [1:0] v$SR_4536_out0;
wire  [1:0] v$SR_4537_out0;
wire  [1:0] v$SR_4538_out0;
wire  [1:0] v$SR_4539_out0;
wire  [1:0] v$XOR1_5225_out0;
wire  [1:0] v$XOR1_5226_out0;
wire  [1:0] v$XOR1_8639_out0;
wire  [1:0] v$XOR1_8640_out0;
wire  [1:0] v$XOR2_19103_out0;
wire  [1:0] v$XOR2_19104_out0;
wire  [1:0] v$XOR3_4194_out0;
wire  [1:0] v$XOR3_4195_out0;
wire  [1:0] v$Y_6731_out0;
wire  [1:0] v$Y_6732_out0;
wire  [1:0] v$Y_6733_out0;
wire  [1:0] v$Y_6734_out0;
wire  [1:0] v$Y_6735_out0;
wire  [1:0] v$Y_6736_out0;
wire  [1:0] v$Y_6737_out0;
wire  [1:0] v$Y_6738_out0;
wire  [1:0] v$Y_6739_out0;
wire  [1:0] v$Y_6740_out0;
wire  [1:0] v$Y_6741_out0;
wire  [1:0] v$Y_6742_out0;
wire  [1:0] v$Y_6743_out0;
wire  [1:0] v$Y_6744_out0;
wire  [1:0] v$Y_6745_out0;
wire  [1:0] v$Y_6746_out0;
wire  [1:0] v$Y_6747_out0;
wire  [1:0] v$Y_6748_out0;
wire  [1:0] v$Y_6749_out0;
wire  [1:0] v$Y_6750_out0;
wire  [1:0] v$Y_6751_out0;
wire  [1:0] v$Y_6752_out0;
wire  [1:0] v$Y_6753_out0;
wire  [1:0] v$Y_6754_out0;
wire  [1:0] v$Y_6755_out0;
wire  [1:0] v$Y_6756_out0;
wire  [1:0] v$Y_6757_out0;
wire  [1:0] v$Y_6758_out0;
wire  [1:0] v$Y_6759_out0;
wire  [1:0] v$Y_6760_out0;
wire  [1:0] v$Y_6761_out0;
wire  [1:0] v$Y_6762_out0;
wire  [1:0] v$Y_6763_out0;
wire  [1:0] v$Y_6764_out0;
wire  [1:0] v$Y_6765_out0;
wire  [1:0] v$Y_6766_out0;
wire  [1:0] v$_1012_out0;
wire  [1:0] v$_1013_out0;
wire  [1:0] v$_10333_out0;
wire  [1:0] v$_10334_out0;
wire  [1:0] v$_10339_out0;
wire  [1:0] v$_10340_out0;
wire  [1:0] v$_10689_out0;
wire  [1:0] v$_10690_out0;
wire  [1:0] v$_10691_out0;
wire  [1:0] v$_10692_out0;
wire  [1:0] v$_10693_out0;
wire  [1:0] v$_10694_out0;
wire  [1:0] v$_10898_out1;
wire  [1:0] v$_10899_out1;
wire  [1:0] v$_10900_out1;
wire  [1:0] v$_10901_out1;
wire  [1:0] v$_10902_out1;
wire  [1:0] v$_10903_out1;
wire  [1:0] v$_11264_out1;
wire  [1:0] v$_11265_out1;
wire  [1:0] v$_11266_out1;
wire  [1:0] v$_11267_out1;
wire  [1:0] v$_11268_out1;
wire  [1:0] v$_11269_out1;
wire  [1:0] v$_11286_out0;
wire  [1:0] v$_11287_out0;
wire  [1:0] v$_11306_out0;
wire  [1:0] v$_11306_out1;
wire  [1:0] v$_11307_out0;
wire  [1:0] v$_11307_out1;
wire  [1:0] v$_11413_out1;
wire  [1:0] v$_11414_out1;
wire  [1:0] v$_11415_out1;
wire  [1:0] v$_11416_out1;
wire  [1:0] v$_11417_out1;
wire  [1:0] v$_11418_out1;
wire  [1:0] v$_11463_out0;
wire  [1:0] v$_11464_out0;
wire  [1:0] v$_11465_out0;
wire  [1:0] v$_11466_out0;
wire  [1:0] v$_11467_out0;
wire  [1:0] v$_11468_out0;
wire  [1:0] v$_11481_out0;
wire  [1:0] v$_11482_out0;
wire  [1:0] v$_11596_out1;
wire  [1:0] v$_11597_out1;
wire  [1:0] v$_11598_out1;
wire  [1:0] v$_11599_out1;
wire  [1:0] v$_11600_out1;
wire  [1:0] v$_11601_out1;
wire  [1:0] v$_12388_out0;
wire  [1:0] v$_12388_out1;
wire  [1:0] v$_12389_out0;
wire  [1:0] v$_12389_out1;
wire  [1:0] v$_13411_out0;
wire  [1:0] v$_13411_out1;
wire  [1:0] v$_13412_out0;
wire  [1:0] v$_13412_out1;
wire  [1:0] v$_13413_out0;
wire  [1:0] v$_13413_out1;
wire  [1:0] v$_13414_out0;
wire  [1:0] v$_13414_out1;
wire  [1:0] v$_13415_out0;
wire  [1:0] v$_13415_out1;
wire  [1:0] v$_13416_out0;
wire  [1:0] v$_13416_out1;
wire  [1:0] v$_13417_out0;
wire  [1:0] v$_13417_out1;
wire  [1:0] v$_13418_out0;
wire  [1:0] v$_13418_out1;
wire  [1:0] v$_13419_out0;
wire  [1:0] v$_13419_out1;
wire  [1:0] v$_13420_out0;
wire  [1:0] v$_13420_out1;
wire  [1:0] v$_13421_out0;
wire  [1:0] v$_13421_out1;
wire  [1:0] v$_13422_out0;
wire  [1:0] v$_13422_out1;
wire  [1:0] v$_1347_out0;
wire  [1:0] v$_1348_out0;
wire  [1:0] v$_1349_out0;
wire  [1:0] v$_1350_out0;
wire  [1:0] v$_1351_out0;
wire  [1:0] v$_1352_out0;
wire  [1:0] v$_13641_out0;
wire  [1:0] v$_13642_out0;
wire  [1:0] v$_13729_out0;
wire  [1:0] v$_13729_out1;
wire  [1:0] v$_13730_out0;
wire  [1:0] v$_13730_out1;
wire  [1:0] v$_13803_out0;
wire  [1:0] v$_13804_out0;
wire  [1:0] v$_13839_out0;
wire  [1:0] v$_13839_out1;
wire  [1:0] v$_13840_out0;
wire  [1:0] v$_13840_out1;
wire  [1:0] v$_13867_out0;
wire  [1:0] v$_13867_out1;
wire  [1:0] v$_13868_out0;
wire  [1:0] v$_13868_out1;
wire  [1:0] v$_13873_out1;
wire  [1:0] v$_13874_out1;
wire  [1:0] v$_13877_out0;
wire  [1:0] v$_13878_out0;
wire  [1:0] v$_13879_out0;
wire  [1:0] v$_13880_out0;
wire  [1:0] v$_13881_out0;
wire  [1:0] v$_13882_out0;
wire  [1:0] v$_13995_out0;
wire  [1:0] v$_13996_out0;
wire  [1:0] v$_14021_out0;
wire  [1:0] v$_14022_out0;
wire  [1:0] v$_14023_out0;
wire  [1:0] v$_14024_out0;
wire  [1:0] v$_14025_out0;
wire  [1:0] v$_14026_out0;
wire  [1:0] v$_1429_out0;
wire  [1:0] v$_1430_out0;
wire  [1:0] v$_1462_out1;
wire  [1:0] v$_1463_out1;
wire  [1:0] v$_1464_out1;
wire  [1:0] v$_1465_out1;
wire  [1:0] v$_1466_out1;
wire  [1:0] v$_1467_out1;
wire  [1:0] v$_14777_out0;
wire  [1:0] v$_14778_out0;
wire  [1:0] v$_14779_out0;
wire  [1:0] v$_14780_out0;
wire  [1:0] v$_14814_out0;
wire  [1:0] v$_14815_out0;
wire  [1:0] v$_1515_out1;
wire  [1:0] v$_1516_out1;
wire  [1:0] v$_1517_out1;
wire  [1:0] v$_1518_out1;
wire  [1:0] v$_1519_out1;
wire  [1:0] v$_1520_out1;
wire  [1:0] v$_15215_out0;
wire  [1:0] v$_15216_out0;
wire  [1:0] v$_15382_out0;
wire  [1:0] v$_15383_out0;
wire  [1:0] v$_15446_out0;
wire  [1:0] v$_15447_out0;
wire  [1:0] v$_15448_out0;
wire  [1:0] v$_15449_out0;
wire  [1:0] v$_15450_out0;
wire  [1:0] v$_15451_out0;
wire  [1:0] v$_15509_out0;
wire  [1:0] v$_15510_out0;
wire  [1:0] v$_15614_out0;
wire  [1:0] v$_15615_out0;
wire  [1:0] v$_15616_out0;
wire  [1:0] v$_15617_out0;
wire  [1:0] v$_15618_out0;
wire  [1:0] v$_15619_out0;
wire  [1:0] v$_15630_out0;
wire  [1:0] v$_15631_out0;
wire  [1:0] v$_15632_out0;
wire  [1:0] v$_15633_out0;
wire  [1:0] v$_15634_out0;
wire  [1:0] v$_15635_out0;
wire  [1:0] v$_15636_out0;
wire  [1:0] v$_15636_out1;
wire  [1:0] v$_15637_out0;
wire  [1:0] v$_15637_out1;
wire  [1:0] v$_15758_out1;
wire  [1:0] v$_15759_out1;
wire  [1:0] v$_15760_out1;
wire  [1:0] v$_15761_out1;
wire  [1:0] v$_15762_out1;
wire  [1:0] v$_15763_out1;
wire  [1:0] v$_15881_out0;
wire  [1:0] v$_15882_out0;
wire  [1:0] v$_1625_out0;
wire  [1:0] v$_1625_out1;
wire  [1:0] v$_1626_out0;
wire  [1:0] v$_1626_out1;
wire  [1:0] v$_16303_out0;
wire  [1:0] v$_16304_out0;
wire  [1:0] v$_16305_out0;
wire  [1:0] v$_16306_out0;
wire  [1:0] v$_16307_out0;
wire  [1:0] v$_16308_out0;
wire  [1:0] v$_16528_out0;
wire  [1:0] v$_16529_out0;
wire  [1:0] v$_16562_out0;
wire  [1:0] v$_16563_out0;
wire  [1:0] v$_16610_out0;
wire  [1:0] v$_16611_out0;
wire  [1:0] v$_16742_out1;
wire  [1:0] v$_16743_out1;
wire  [1:0] v$_16744_out1;
wire  [1:0] v$_16745_out1;
wire  [1:0] v$_16746_out1;
wire  [1:0] v$_16747_out1;
wire  [1:0] v$_16748_out0;
wire  [1:0] v$_16749_out0;
wire  [1:0] v$_16841_out0;
wire  [1:0] v$_16841_out1;
wire  [1:0] v$_16842_out0;
wire  [1:0] v$_16842_out1;
wire  [1:0] v$_16876_out1;
wire  [1:0] v$_16877_out1;
wire  [1:0] v$_16878_out1;
wire  [1:0] v$_16879_out1;
wire  [1:0] v$_16880_out1;
wire  [1:0] v$_16881_out1;
wire  [1:0] v$_16924_out0;
wire  [1:0] v$_16925_out0;
wire  [1:0] v$_16926_out0;
wire  [1:0] v$_16927_out0;
wire  [1:0] v$_16928_out0;
wire  [1:0] v$_16929_out0;
wire  [1:0] v$_1733_out0;
wire  [1:0] v$_1734_out0;
wire  [1:0] v$_17358_out0;
wire  [1:0] v$_17359_out0;
wire  [1:0] v$_1735_out0;
wire  [1:0] v$_17361_out1;
wire  [1:0] v$_17362_out1;
wire  [1:0] v$_17363_out1;
wire  [1:0] v$_17364_out1;
wire  [1:0] v$_17365_out1;
wire  [1:0] v$_17366_out1;
wire  [1:0] v$_1736_out0;
wire  [1:0] v$_1737_out0;
wire  [1:0] v$_1738_out0;
wire  [1:0] v$_17395_out0;
wire  [1:0] v$_17396_out0;
wire  [1:0] v$_1761_out0;
wire  [1:0] v$_1761_out1;
wire  [1:0] v$_1762_out0;
wire  [1:0] v$_1762_out1;
wire  [1:0] v$_17652_out0;
wire  [1:0] v$_17653_out0;
wire  [1:0] v$_18098_out0;
wire  [1:0] v$_18099_out0;
wire  [1:0] v$_18100_out0;
wire  [1:0] v$_18101_out0;
wire  [1:0] v$_18102_out0;
wire  [1:0] v$_18103_out0;
wire  [1:0] v$_1855_out0;
wire  [1:0] v$_1855_out1;
wire  [1:0] v$_1856_out0;
wire  [1:0] v$_1856_out1;
wire  [1:0] v$_18585_out0;
wire  [1:0] v$_18586_out0;
wire  [1:0] v$_18787_out1;
wire  [1:0] v$_18788_out1;
wire  [1:0] v$_18789_out1;
wire  [1:0] v$_18790_out1;
wire  [1:0] v$_18791_out1;
wire  [1:0] v$_18792_out1;
wire  [1:0] v$_18901_out1;
wire  [1:0] v$_18902_out1;
wire  [1:0] v$_18932_out0;
wire  [1:0] v$_18933_out0;
wire  [1:0] v$_19017_out0;
wire  [1:0] v$_19018_out0;
wire  [1:0] v$_19129_out0;
wire  [1:0] v$_19130_out0;
wire  [1:0] v$_19177_out0;
wire  [1:0] v$_19178_out0;
wire  [1:0] v$_19274_out0;
wire  [1:0] v$_19275_out0;
wire  [1:0] v$_19276_out0;
wire  [1:0] v$_19277_out0;
wire  [1:0] v$_19278_out0;
wire  [1:0] v$_19279_out0;
wire  [1:0] v$_1954_out0;
wire  [1:0] v$_1955_out0;
wire  [1:0] v$_1956_out0;
wire  [1:0] v$_1957_out0;
wire  [1:0] v$_1958_out0;
wire  [1:0] v$_1959_out0;
wire  [1:0] v$_1989_out0;
wire  [1:0] v$_1990_out0;
wire  [1:0] v$_2014_out1;
wire  [1:0] v$_2015_out1;
wire  [1:0] v$_2016_out1;
wire  [1:0] v$_2017_out1;
wire  [1:0] v$_2018_out1;
wire  [1:0] v$_2019_out1;
wire  [1:0] v$_218_out0;
wire  [1:0] v$_218_out1;
wire  [1:0] v$_219_out0;
wire  [1:0] v$_219_out1;
wire  [1:0] v$_237_out0;
wire  [1:0] v$_237_out1;
wire  [1:0] v$_238_out0;
wire  [1:0] v$_238_out1;
wire  [1:0] v$_2471_out0;
wire  [1:0] v$_2472_out0;
wire  [1:0] v$_2493_out0;
wire  [1:0] v$_2493_out1;
wire  [1:0] v$_2494_out0;
wire  [1:0] v$_2494_out1;
wire  [1:0] v$_2613_out1;
wire  [1:0] v$_2646_out0;
wire  [1:0] v$_2647_out0;
wire  [1:0] v$_2648_out0;
wire  [1:0] v$_2649_out0;
wire  [1:0] v$_2650_out0;
wire  [1:0] v$_2651_out0;
wire  [1:0] v$_2810_out1;
wire  [1:0] v$_2866_out0;
wire  [1:0] v$_2867_out0;
wire  [1:0] v$_3064_out0;
wire  [1:0] v$_3065_out0;
wire  [1:0] v$_3066_out0;
wire  [1:0] v$_3067_out0;
wire  [1:0] v$_3068_out0;
wire  [1:0] v$_3069_out0;
wire  [1:0] v$_3129_out1;
wire  [1:0] v$_3130_out1;
wire  [1:0] v$_3131_out1;
wire  [1:0] v$_3132_out1;
wire  [1:0] v$_3133_out1;
wire  [1:0] v$_3134_out1;
wire  [1:0] v$_3363_out0;
wire  [1:0] v$_3364_out0;
wire  [1:0] v$_3826_out0;
wire  [1:0] v$_3827_out0;
wire  [1:0] v$_3828_out0;
wire  [1:0] v$_3829_out0;
wire  [1:0] v$_3830_out0;
wire  [1:0] v$_3831_out0;
wire  [1:0] v$_3881_out0;
wire  [1:0] v$_3881_out1;
wire  [1:0] v$_3882_out0;
wire  [1:0] v$_3882_out1;
wire  [1:0] v$_3967_out0;
wire  [1:0] v$_3968_out0;
wire  [1:0] v$_5301_out0;
wire  [1:0] v$_5302_out0;
wire  [1:0] v$_5360_out0;
wire  [1:0] v$_5360_out1;
wire  [1:0] v$_5361_out0;
wire  [1:0] v$_5361_out1;
wire  [1:0] v$_56_out0;
wire  [1:0] v$_56_out1;
wire  [1:0] v$_57_out0;
wire  [1:0] v$_57_out1;
wire  [1:0] v$_6173_out0;
wire  [1:0] v$_6174_out0;
wire  [1:0] v$_6175_out0;
wire  [1:0] v$_6176_out0;
wire  [1:0] v$_6177_out0;
wire  [1:0] v$_6178_out0;
wire  [1:0] v$_6352_out1;
wire  [1:0] v$_6353_out1;
wire  [1:0] v$_6443_out0;
wire  [1:0] v$_6444_out0;
wire  [1:0] v$_6532_out0;
wire  [1:0] v$_6533_out0;
wire  [1:0] v$_6534_out0;
wire  [1:0] v$_6535_out0;
wire  [1:0] v$_6536_out0;
wire  [1:0] v$_6537_out0;
wire  [1:0] v$_6538_out0;
wire  [1:0] v$_6539_out0;
wire  [1:0] v$_6540_out0;
wire  [1:0] v$_6541_out0;
wire  [1:0] v$_6542_out0;
wire  [1:0] v$_6543_out0;
wire  [1:0] v$_6544_out0;
wire  [1:0] v$_6545_out0;
wire  [1:0] v$_6546_out0;
wire  [1:0] v$_6547_out0;
wire  [1:0] v$_6548_out0;
wire  [1:0] v$_6549_out0;
wire  [1:0] v$_6550_out0;
wire  [1:0] v$_6551_out0;
wire  [1:0] v$_6552_out0;
wire  [1:0] v$_6553_out0;
wire  [1:0] v$_6554_out0;
wire  [1:0] v$_6555_out0;
wire  [1:0] v$_6556_out0;
wire  [1:0] v$_6557_out0;
wire  [1:0] v$_6558_out0;
wire  [1:0] v$_6559_out0;
wire  [1:0] v$_6560_out0;
wire  [1:0] v$_6561_out0;
wire  [1:0] v$_6562_out0;
wire  [1:0] v$_6563_out0;
wire  [1:0] v$_6564_out0;
wire  [1:0] v$_6565_out0;
wire  [1:0] v$_6566_out0;
wire  [1:0] v$_6567_out0;
wire  [1:0] v$_710_out0;
wire  [1:0] v$_711_out0;
wire  [1:0] v$_712_out0;
wire  [1:0] v$_713_out0;
wire  [1:0] v$_714_out0;
wire  [1:0] v$_715_out0;
wire  [1:0] v$_7355_out1;
wire  [1:0] v$_7356_out1;
wire  [1:0] v$_7357_out1;
wire  [1:0] v$_7358_out1;
wire  [1:0] v$_7359_out1;
wire  [1:0] v$_7360_out1;
wire  [1:0] v$_7687_out0;
wire  [1:0] v$_7687_out1;
wire  [1:0] v$_7688_out0;
wire  [1:0] v$_7688_out1;
wire  [1:0] v$_7786_out0;
wire  [1:0] v$_7786_out1;
wire  [1:0] v$_7787_out0;
wire  [1:0] v$_7787_out1;
wire  [1:0] v$_7874_out0;
wire  [1:0] v$_7875_out0;
wire  [1:0] v$_7876_out0;
wire  [1:0] v$_7877_out0;
wire  [1:0] v$_7878_out0;
wire  [1:0] v$_7879_out0;
wire  [1:0] v$_8051_out0;
wire  [1:0] v$_8052_out0;
wire  [1:0] v$_8088_out1;
wire  [1:0] v$_8089_out1;
wire  [1:0] v$_8090_out1;
wire  [1:0] v$_8091_out1;
wire  [1:0] v$_8092_out1;
wire  [1:0] v$_8093_out1;
wire  [1:0] v$_8193_out0;
wire  [1:0] v$_8194_out0;
wire  [1:0] v$_8195_out0;
wire  [1:0] v$_8196_out0;
wire  [1:0] v$_8197_out0;
wire  [1:0] v$_8198_out0;
wire  [1:0] v$_82_out0;
wire  [1:0] v$_83_out0;
wire  [1:0] v$_84_out0;
wire  [1:0] v$_8517_out0;
wire  [1:0] v$_8517_out1;
wire  [1:0] v$_8518_out0;
wire  [1:0] v$_8518_out1;
wire  [1:0] v$_85_out0;
wire  [1:0] v$_8641_out0;
wire  [1:0] v$_8642_out0;
wire  [1:0] v$_8643_out0;
wire  [1:0] v$_8644_out0;
wire  [1:0] v$_8645_out0;
wire  [1:0] v$_8646_out0;
wire  [1:0] v$_86_out0;
wire  [1:0] v$_8758_out0;
wire  [1:0] v$_8758_out1;
wire  [1:0] v$_8759_out0;
wire  [1:0] v$_8759_out1;
wire  [1:0] v$_8760_out0;
wire  [1:0] v$_8760_out1;
wire  [1:0] v$_8761_out0;
wire  [1:0] v$_8761_out1;
wire  [1:0] v$_8762_out0;
wire  [1:0] v$_8762_out1;
wire  [1:0] v$_8763_out0;
wire  [1:0] v$_8763_out1;
wire  [1:0] v$_8764_out0;
wire  [1:0] v$_8764_out1;
wire  [1:0] v$_8765_out0;
wire  [1:0] v$_8765_out1;
wire  [1:0] v$_8766_out0;
wire  [1:0] v$_8766_out1;
wire  [1:0] v$_8767_out0;
wire  [1:0] v$_8767_out1;
wire  [1:0] v$_8768_out0;
wire  [1:0] v$_8768_out1;
wire  [1:0] v$_8769_out0;
wire  [1:0] v$_8769_out1;
wire  [1:0] v$_87_out0;
wire  [1:0] v$_9235_out0;
wire  [1:0] v$_9236_out0;
wire  [1:0] v$_9237_out0;
wire  [1:0] v$_9238_out0;
wire  [1:0] v$_9239_out0;
wire  [1:0] v$_9240_out0;
wire  [1:0] v$_9389_out1;
wire  [1:0] v$_9390_out1;
wire  [1:0] v$_9391_out1;
wire  [1:0] v$_9392_out1;
wire  [1:0] v$_9393_out1;
wire  [1:0] v$_9394_out1;
wire  [1:0] v$_9795_out0;
wire  [1:0] v$_9795_out1;
wire  [1:0] v$_9796_out0;
wire  [1:0] v$_9796_out1;
wire  [1:0] v$_9811_out0;
wire  [1:0] v$_9812_out0;
wire  [1:0] v$_9831_out0;
wire  [1:0] v$_9832_out0;
wire  [21:0] v$SEL1_15978_out0;
wire  [21:0] v$SEL1_15983_out0;
wire  [21:0] v$SEL1_15988_out0;
wire  [21:0] v$SEL1_15993_out0;
wire  [21:0] v$SEL1_15998_out0;
wire  [21:0] v$SEL1_16003_out0;
wire  [21:0] v$SEL1_16009_out0;
wire  [21:0] v$SEL1_16014_out0;
wire  [21:0] v$SEL1_16019_out0;
wire  [21:0] v$SEL1_16024_out0;
wire  [21:0] v$SEL1_16029_out0;
wire  [21:0] v$SEL1_16034_out0;
wire  [21:0] v$SEL1_9050_out0;
wire  [21:0] v$SEL1_9055_out0;
wire  [21:0] v$SEL1_9060_out0;
wire  [21:0] v$SEL1_9065_out0;
wire  [21:0] v$SEL1_9070_out0;
wire  [21:0] v$SEL1_9075_out0;
wire  [21:0] v$SEL1_9081_out0;
wire  [21:0] v$SEL1_9086_out0;
wire  [21:0] v$SEL1_9091_out0;
wire  [21:0] v$SEL1_9096_out0;
wire  [21:0] v$SEL1_9101_out0;
wire  [21:0] v$SEL1_9106_out0;
wire  [22:0] v$A$MANTISA$MUL_2851_out0;
wire  [22:0] v$A$MANTISA$MUL_2852_out0;
wire  [22:0] v$A$MANTISA_12397_out0;
wire  [22:0] v$A$MANTISA_12398_out0;
wire  [22:0] v$A$MANTISA_15148_out0;
wire  [22:0] v$A$MANTISA_15149_out0;
wire  [22:0] v$A$MANTISA_18529_out0;
wire  [22:0] v$A$MANTISA_18530_out0;
wire  [22:0] v$B$MANTISA$MUL_8473_out0;
wire  [22:0] v$B$MANTISA$MUL_8474_out0;
wire  [22:0] v$B$MANTISA_3213_out0;
wire  [22:0] v$B$MANTISA_3214_out0;
wire  [22:0] v$B$MANTISA_4226_out0;
wire  [22:0] v$B$MANTISA_4227_out0;
wire  [22:0] v$B$MANTISA_5124_out0;
wire  [22:0] v$B$MANTISA_5125_out0;
wire  [22:0] v$C5_16212_out0;
wire  [22:0] v$C5_16213_out0;
wire  [22:0] v$MANTISA$ADDITION_13751_out0;
wire  [22:0] v$MANTISA$ADDITION_13752_out0;
wire  [22:0] v$MANTISA$RESULT$BEFORE$MERGE_19325_out0;
wire  [22:0] v$MANTISA$RESULT$BEFORE$MERGE_19326_out0;
wire  [22:0] v$MANTISA$RESULT$FPU$ADDER_12474_out0;
wire  [22:0] v$MANTISA$RESULT$FPU$ADDER_12475_out0;
wire  [22:0] v$MANTISA$RESULT_6779_out0;
wire  [22:0] v$MANTISA$RESULT_6780_out0;
wire  [22:0] v$MUX1_2096_out0;
wire  [22:0] v$MUX1_2097_out0;
wire  [22:0] v$MUX2_1765_out0;
wire  [22:0] v$MUX2_1766_out0;
wire  [22:0] v$MUX2_3183_out0;
wire  [22:0] v$MUX2_3184_out0;
wire  [22:0] v$MUX6_13339_out0;
wire  [22:0] v$MUX6_13340_out0;
wire  [22:0] v$MUX7_13312_out0;
wire  [22:0] v$MUX7_13313_out0;
wire  [22:0] v$MUX8_7366_out0;
wire  [22:0] v$MUX8_7367_out0;
wire  [22:0] v$OUT1_10858_out0;
wire  [22:0] v$OUT1_10859_out0;
wire  [22:0] v$SEL1_14967_out0;
wire  [22:0] v$SEL1_14968_out0;
wire  [22:0] v$SEL1_15976_out0;
wire  [22:0] v$SEL1_15981_out0;
wire  [22:0] v$SEL1_15986_out0;
wire  [22:0] v$SEL1_15989_out0;
wire  [22:0] v$SEL1_15996_out0;
wire  [22:0] v$SEL1_15999_out0;
wire  [22:0] v$SEL1_16004_out0;
wire  [22:0] v$SEL1_16007_out0;
wire  [22:0] v$SEL1_16012_out0;
wire  [22:0] v$SEL1_16017_out0;
wire  [22:0] v$SEL1_16020_out0;
wire  [22:0] v$SEL1_16027_out0;
wire  [22:0] v$SEL1_16030_out0;
wire  [22:0] v$SEL1_16035_out0;
wire  [22:0] v$SEL1_16347_out0;
wire  [22:0] v$SEL1_16348_out0;
wire  [22:0] v$SEL1_6308_out0;
wire  [22:0] v$SEL1_6309_out0;
wire  [22:0] v$SEL1_9048_out0;
wire  [22:0] v$SEL1_9053_out0;
wire  [22:0] v$SEL1_9058_out0;
wire  [22:0] v$SEL1_9061_out0;
wire  [22:0] v$SEL1_9068_out0;
wire  [22:0] v$SEL1_9071_out0;
wire  [22:0] v$SEL1_9076_out0;
wire  [22:0] v$SEL1_9079_out0;
wire  [22:0] v$SEL1_9084_out0;
wire  [22:0] v$SEL1_9089_out0;
wire  [22:0] v$SEL1_9092_out0;
wire  [22:0] v$SEL1_9099_out0;
wire  [22:0] v$SEL1_9102_out0;
wire  [22:0] v$SEL1_9107_out0;
wire  [22:0] v$SEL2_11519_out0;
wire  [22:0] v$SEL2_11520_out0;
wire  [22:0] v$SEL2_6314_out0;
wire  [22:0] v$SEL2_6315_out0;
wire  [22:0] v$SEL3_12468_out0;
wire  [22:0] v$SEL3_12469_out0;
wire  [22:0] v$SEL3_14851_out0;
wire  [22:0] v$SEL3_14852_out0;
wire  [22:0] v$SEL4_13548_out0;
wire  [22:0] v$SEL4_13549_out0;
wire  [22:0] v$SEL4_2485_out0;
wire  [22:0] v$SEL4_2486_out0;
wire  [22:0] v$SEL4_7880_out0;
wire  [22:0] v$SEL4_7881_out0;
wire  [22:0] v$SEL5_10785_out0;
wire  [22:0] v$SEL5_10786_out0;
wire  [22:0] v$SEL6_4609_out0;
wire  [22:0] v$SEL6_4610_out0;
wire  [22:0] v$SEL8_18134_out0;
wire  [22:0] v$SEL8_18135_out0;
wire  [22:0] v$SEL8_7593_out0;
wire  [22:0] v$SEL8_7594_out0;
wire  [22:0] v$_16853_out0;
wire  [22:0] v$_16854_out0;
wire  [22:0] v$_1843_out0;
wire  [22:0] v$_1844_out0;
wire  [22:0] v$_18695_out0;
wire  [22:0] v$_18696_out0;
wire  [22:0] v$_2436_out0;
wire  [22:0] v$_2437_out0;
wire  [23:0] v$A$MANTISA$COMPARATOR_7820_out0;
wire  [23:0] v$A$MANTISA$COMPARATOR_7821_out0;
wire  [23:0] v$A$MANTISA_3937_out0;
wire  [23:0] v$A$MANTISA_3938_out0;
wire  [23:0] v$A$MANTISSA_13764_out0;
wire  [23:0] v$A$MANTISSA_13765_out0;
wire  [23:0] v$A$VIEW_11537_out0;
wire  [23:0] v$A$VIEW_11538_out0;
wire  [23:0] v$A1_14170_out0;
wire  [23:0] v$A1_14171_out0;
wire  [23:0] v$A1_14172_out0;
wire  [23:0] v$A1_14173_out0;
wire  [23:0] v$A1_14174_out0;
wire  [23:0] v$A1_14175_out0;
wire  [23:0] v$ADDER$A_3875_out0;
wire  [23:0] v$ADDER$A_3876_out0;
wire  [23:0] v$ADDER$B_6686_out0;
wire  [23:0] v$ADDER$B_6687_out0;
wire  [23:0] v$A_14857_out0;
wire  [23:0] v$A_14858_out0;
wire  [23:0] v$A_3673_out0;
wire  [23:0] v$A_3674_out0;
wire  [23:0] v$B$MANTISA$COMPARATOR_16468_out0;
wire  [23:0] v$B$MANTISA$COMPARATOR_16469_out0;
wire  [23:0] v$B$MANTISA_16181_out0;
wire  [23:0] v$B$MANTISA_16182_out0;
wire  [23:0] v$B$MANTISSA_2870_out0;
wire  [23:0] v$B$MANTISSA_2871_out0;
wire  [23:0] v$B$SHIFTED_14379_out0;
wire  [23:0] v$B$SHIFTED_14380_out0;
wire  [23:0] v$B$VIEW_6013_out0;
wire  [23:0] v$B$VIEW_6014_out0;
wire  [23:0] v$B2_8720_out0;
wire  [23:0] v$B2_8721_out0;
wire  [23:0] v$B2_8722_out0;
wire  [23:0] v$B2_8723_out0;
wire  [23:0] v$B2_8724_out0;
wire  [23:0] v$B2_8725_out0;
wire  [23:0] v$B_14138_out0;
wire  [23:0] v$B_14139_out0;
wire  [23:0] v$B_80_out0;
wire  [23:0] v$B_81_out0;
wire  [23:0] v$C1_16843_out0;
wire  [23:0] v$C1_16844_out0;
wire  [23:0] v$C1_4623_out0;
wire  [23:0] v$C1_4624_out0;
wire  [23:0] v$C1_4625_out0;
wire  [23:0] v$C1_4626_out0;
wire  [23:0] v$C1_4627_out0;
wire  [23:0] v$C1_4628_out0;
wire  [23:0] v$C1_4629_out0;
wire  [23:0] v$C1_4630_out0;
wire  [23:0] v$C3_19045_out0;
wire  [23:0] v$C3_19046_out0;
wire  [23:0] v$C4_18589_out0;
wire  [23:0] v$C4_18590_out0;
wire  [23:0] v$C7_15247_out0;
wire  [23:0] v$C7_15248_out0;
wire  [23:0] v$C8_14199_out0;
wire  [23:0] v$C8_14200_out0;
wire  [23:0] v$C9_15847_out0;
wire  [23:0] v$C9_15848_out0;
wire  [23:0] v$END1_10352_out0;
wire  [23:0] v$END1_10353_out0;
wire  [23:0] v$END_2032_out0;
wire  [23:0] v$END_2033_out0;
wire  [23:0] v$FINAL$RESULT_2764_out0;
wire  [23:0] v$FINAL$RESULT_2765_out0;
wire  [23:0] v$IGNORE_13217_out0;
wire  [23:0] v$IGNORE_13218_out0;
wire  [23:0] v$IN_11584_out0;
wire  [23:0] v$IN_11585_out0;
wire  [23:0] v$IN_11586_out0;
wire  [23:0] v$IN_11587_out0;
wire  [23:0] v$IN_12204_out0;
wire  [23:0] v$IN_12205_out0;
wire  [23:0] v$IN_12206_out0;
wire  [23:0] v$IN_12207_out0;
wire  [23:0] v$IN_12352_out0;
wire  [23:0] v$IN_12353_out0;
wire  [23:0] v$IN_12354_out0;
wire  [23:0] v$IN_12355_out0;
wire  [23:0] v$IN_12356_out0;
wire  [23:0] v$IN_12357_out0;
wire  [23:0] v$IN_12358_out0;
wire  [23:0] v$IN_12359_out0;
wire  [23:0] v$IN_12360_out0;
wire  [23:0] v$IN_12361_out0;
wire  [23:0] v$IN_12362_out0;
wire  [23:0] v$IN_12363_out0;
wire  [23:0] v$IN_13743_out0;
wire  [23:0] v$IN_13744_out0;
wire  [23:0] v$IN_13745_out0;
wire  [23:0] v$IN_13746_out0;
wire  [23:0] v$IN_13747_out0;
wire  [23:0] v$IN_13748_out0;
wire  [23:0] v$IN_13749_out0;
wire  [23:0] v$IN_13750_out0;
wire  [23:0] v$IN_14140_out0;
wire  [23:0] v$IN_14142_out0;
wire  [23:0] v$IN_14144_out0;
wire  [23:0] v$IN_14146_out0;
wire  [23:0] v$IN_16196_out0;
wire  [23:0] v$IN_16197_out0;
wire  [23:0] v$IN_16198_out0;
wire  [23:0] v$IN_16199_out0;
wire  [23:0] v$IN_16200_out0;
wire  [23:0] v$IN_16201_out0;
wire  [23:0] v$IN_16202_out0;
wire  [23:0] v$IN_16203_out0;
wire  [23:0] v$IN_16204_out0;
wire  [23:0] v$IN_16205_out0;
wire  [23:0] v$IN_16206_out0;
wire  [23:0] v$IN_16207_out0;
wire  [23:0] v$IN_18605_out0;
wire  [23:0] v$IN_18606_out0;
wire  [23:0] v$IN_18864_out0;
wire  [23:0] v$IN_18865_out0;
wire  [23:0] v$IN_18866_out0;
wire  [23:0] v$IN_18867_out0;
wire  [23:0] v$IN_4036_out0;
wire  [23:0] v$IN_4037_out0;
wire  [23:0] v$IN_4038_out0;
wire  [23:0] v$IN_4039_out0;
wire  [23:0] v$IN_4040_out0;
wire  [23:0] v$IN_4041_out0;
wire  [23:0] v$IN_4042_out0;
wire  [23:0] v$IN_4043_out0;
wire  [23:0] v$IN_4044_out0;
wire  [23:0] v$IN_4045_out0;
wire  [23:0] v$IN_4046_out0;
wire  [23:0] v$IN_4047_out0;
wire  [23:0] v$IN_4048_out0;
wire  [23:0] v$IN_4049_out0;
wire  [23:0] v$IN_4050_out0;
wire  [23:0] v$IN_4051_out0;
wire  [23:0] v$IN_4052_out0;
wire  [23:0] v$IN_4053_out0;
wire  [23:0] v$IN_4348_out0;
wire  [23:0] v$IN_4349_out0;
wire  [23:0] v$IN_4350_out0;
wire  [23:0] v$IN_4351_out0;
wire  [23:0] v$IN_5233_out0;
wire  [23:0] v$IN_5234_out0;
wire  [23:0] v$IN_5235_out0;
wire  [23:0] v$IN_5236_out0;
wire  [23:0] v$IN_5237_out0;
wire  [23:0] v$IN_5238_out0;
wire  [23:0] v$IN_5239_out0;
wire  [23:0] v$IN_5240_out0;
wire  [23:0] v$IN_5241_out0;
wire  [23:0] v$IN_5242_out0;
wire  [23:0] v$IN_5243_out0;
wire  [23:0] v$IN_5244_out0;
wire  [23:0] v$IN_5245_out0;
wire  [23:0] v$IN_5246_out0;
wire  [23:0] v$IN_5247_out0;
wire  [23:0] v$IN_5248_out0;
wire  [23:0] v$IN_5249_out0;
wire  [23:0] v$IN_5250_out0;
wire  [23:0] v$IN_5251_out0;
wire  [23:0] v$IN_5252_out0;
wire  [23:0] v$IN_5365_out0;
wire  [23:0] v$IN_5366_out0;
wire  [23:0] v$IN_5367_out0;
wire  [23:0] v$IN_5368_out0;
wire  [23:0] v$IN_5369_out0;
wire  [23:0] v$IN_5370_out0;
wire  [23:0] v$IN_5371_out0;
wire  [23:0] v$IN_5372_out0;
wire  [23:0] v$IN_5373_out0;
wire  [23:0] v$IN_5374_out0;
wire  [23:0] v$IN_5375_out0;
wire  [23:0] v$IN_5376_out0;
wire  [23:0] v$IN_5377_out0;
wire  [23:0] v$IN_5378_out0;
wire  [23:0] v$IN_5379_out0;
wire  [23:0] v$IN_5380_out0;
wire  [23:0] v$IN_5381_out0;
wire  [23:0] v$IN_5382_out0;
wire  [23:0] v$IN_5383_out0;
wire  [23:0] v$IN_5384_out0;
wire  [23:0] v$IN_5385_out0;
wire  [23:0] v$IN_5386_out0;
wire  [23:0] v$IN_5387_out0;
wire  [23:0] v$IN_5388_out0;
wire  [23:0] v$IN_5389_out0;
wire  [23:0] v$IN_5390_out0;
wire  [23:0] v$IN_5391_out0;
wire  [23:0] v$IN_5392_out0;
wire  [23:0] v$IN_5393_out0;
wire  [23:0] v$IN_5394_out0;
wire  [23:0] v$IN_5395_out0;
wire  [23:0] v$IN_5396_out0;
wire  [23:0] v$IN_5397_out0;
wire  [23:0] v$IN_5398_out0;
wire  [23:0] v$IN_5399_out0;
wire  [23:0] v$IN_5400_out0;
wire  [23:0] v$IN_5401_out0;
wire  [23:0] v$IN_5402_out0;
wire  [23:0] v$IN_5403_out0;
wire  [23:0] v$IN_5404_out0;
wire  [23:0] v$IN_5405_out0;
wire  [23:0] v$IN_5406_out0;
wire  [23:0] v$IN_5407_out0;
wire  [23:0] v$IN_5408_out0;
wire  [23:0] v$IN_5409_out0;
wire  [23:0] v$IN_5410_out0;
wire  [23:0] v$IN_5411_out0;
wire  [23:0] v$IN_5412_out0;
wire  [23:0] v$IN_5413_out0;
wire  [23:0] v$IN_5414_out0;
wire  [23:0] v$IN_5415_out0;
wire  [23:0] v$IN_5416_out0;
wire  [23:0] v$IN_5417_out0;
wire  [23:0] v$IN_5418_out0;
wire  [23:0] v$IN_5419_out0;
wire  [23:0] v$IN_5420_out0;
wire  [23:0] v$IN_5421_out0;
wire  [23:0] v$IN_5422_out0;
wire  [23:0] v$IN_5423_out0;
wire  [23:0] v$IN_5424_out0;
wire  [23:0] v$IN_5425_out0;
wire  [23:0] v$IN_5426_out0;
wire  [23:0] v$IN_8605_out0;
wire  [23:0] v$IN_8606_out0;
wire  [23:0] v$IN_8607_out0;
wire  [23:0] v$IN_8608_out0;
wire  [23:0] v$LZD$INPUT_9184_out0;
wire  [23:0] v$LZD$INPUT_9185_out0;
wire  [23:0] v$MULTIPLIER$OUT_15586_out0;
wire  [23:0] v$MULTIPLIER$OUT_15587_out0;
wire  [23:0] v$MULTIPLIER$OUT_9712_out0;
wire  [23:0] v$MULTIPLIER$OUT_9713_out0;
wire  [23:0] v$MUX1_12191_out0;
wire  [23:0] v$MUX1_12192_out0;
wire  [23:0] v$MUX1_12193_out0;
wire  [23:0] v$MUX1_12194_out0;
wire  [23:0] v$MUX1_12195_out0;
wire  [23:0] v$MUX1_12196_out0;
wire  [23:0] v$MUX1_12197_out0;
wire  [23:0] v$MUX1_12198_out0;
wire  [23:0] v$MUX1_14796_out0;
wire  [23:0] v$MUX1_14797_out0;
wire  [23:0] v$MUX1_2543_out0;
wire  [23:0] v$MUX1_2544_out0;
wire  [23:0] v$MUX1_2545_out0;
wire  [23:0] v$MUX1_2546_out0;
wire  [23:0] v$MUX1_2547_out0;
wire  [23:0] v$MUX1_2548_out0;
wire  [23:0] v$MUX1_2549_out0;
wire  [23:0] v$MUX1_2550_out0;
wire  [23:0] v$MUX1_2551_out0;
wire  [23:0] v$MUX1_2552_out0;
wire  [23:0] v$MUX1_2553_out0;
wire  [23:0] v$MUX1_2554_out0;
wire  [23:0] v$MUX1_2555_out0;
wire  [23:0] v$MUX1_2556_out0;
wire  [23:0] v$MUX1_2557_out0;
wire  [23:0] v$MUX1_2558_out0;
wire  [23:0] v$MUX1_2559_out0;
wire  [23:0] v$MUX1_2560_out0;
wire  [23:0] v$MUX1_2561_out0;
wire  [23:0] v$MUX1_2562_out0;
wire  [23:0] v$MUX1_2563_out0;
wire  [23:0] v$MUX1_2564_out0;
wire  [23:0] v$MUX1_2565_out0;
wire  [23:0] v$MUX1_2566_out0;
wire  [23:0] v$MUX1_2567_out0;
wire  [23:0] v$MUX1_2568_out0;
wire  [23:0] v$MUX1_2569_out0;
wire  [23:0] v$MUX1_2570_out0;
wire  [23:0] v$MUX1_2571_out0;
wire  [23:0] v$MUX1_2572_out0;
wire  [23:0] v$MUX1_2573_out0;
wire  [23:0] v$MUX1_2574_out0;
wire  [23:0] v$MUX1_2575_out0;
wire  [23:0] v$MUX1_2576_out0;
wire  [23:0] v$MUX1_2577_out0;
wire  [23:0] v$MUX1_2578_out0;
wire  [23:0] v$MUX1_2579_out0;
wire  [23:0] v$MUX1_2580_out0;
wire  [23:0] v$MUX1_2581_out0;
wire  [23:0] v$MUX1_2582_out0;
wire  [23:0] v$MUX1_2583_out0;
wire  [23:0] v$MUX1_2584_out0;
wire  [23:0] v$MUX1_2585_out0;
wire  [23:0] v$MUX1_2586_out0;
wire  [23:0] v$MUX1_2587_out0;
wire  [23:0] v$MUX1_2588_out0;
wire  [23:0] v$MUX1_2589_out0;
wire  [23:0] v$MUX1_2590_out0;
wire  [23:0] v$MUX1_2591_out0;
wire  [23:0] v$MUX1_2592_out0;
wire  [23:0] v$MUX1_2593_out0;
wire  [23:0] v$MUX1_2594_out0;
wire  [23:0] v$MUX1_2595_out0;
wire  [23:0] v$MUX1_2596_out0;
wire  [23:0] v$MUX1_2597_out0;
wire  [23:0] v$MUX1_2598_out0;
wire  [23:0] v$MUX1_2599_out0;
wire  [23:0] v$MUX1_2600_out0;
wire  [23:0] v$MUX1_2601_out0;
wire  [23:0] v$MUX1_2602_out0;
wire  [23:0] v$MUX1_2603_out0;
wire  [23:0] v$MUX1_2604_out0;
wire  [23:0] v$MUX1_3094_out0;
wire  [23:0] v$MUX1_3095_out0;
wire  [23:0] v$MUX2_13050_out0;
wire  [23:0] v$MUX2_13051_out0;
wire  [23:0] v$MUX2_15434_out0;
wire  [23:0] v$MUX2_15435_out0;
wire  [23:0] v$MUX2_15436_out0;
wire  [23:0] v$MUX2_15437_out0;
wire  [23:0] v$MUX2_15438_out0;
wire  [23:0] v$MUX2_15439_out0;
wire  [23:0] v$MUX2_15817_out0;
wire  [23:0] v$MUX2_15818_out0;
wire  [23:0] v$MUX2_15819_out0;
wire  [23:0] v$MUX2_15820_out0;
wire  [23:0] v$MUX2_15821_out0;
wire  [23:0] v$MUX2_15822_out0;
wire  [23:0] v$MUX2_15823_out0;
wire  [23:0] v$MUX2_15824_out0;
wire  [23:0] v$MUX2_15825_out0;
wire  [23:0] v$MUX2_15826_out0;
wire  [23:0] v$MUX2_15827_out0;
wire  [23:0] v$MUX2_15828_out0;
wire  [23:0] v$MUX2_19185_out0;
wire  [23:0] v$MUX2_19186_out0;
wire  [23:0] v$MUX2_19187_out0;
wire  [23:0] v$MUX2_19188_out0;
wire  [23:0] v$MUX2_19189_out0;
wire  [23:0] v$MUX2_19190_out0;
wire  [23:0] v$MUX2_19191_out0;
wire  [23:0] v$MUX2_19192_out0;
wire  [23:0] v$MUX2_19193_out0;
wire  [23:0] v$MUX2_19194_out0;
wire  [23:0] v$MUX2_19195_out0;
wire  [23:0] v$MUX2_19196_out0;
wire  [23:0] v$MUX2_2670_out0;
wire  [23:0] v$MUX2_2671_out0;
wire  [23:0] v$MUX2_2672_out0;
wire  [23:0] v$MUX2_2673_out0;
wire  [23:0] v$MUX2_2674_out0;
wire  [23:0] v$MUX2_2675_out0;
wire  [23:0] v$MUX2_2676_out0;
wire  [23:0] v$MUX2_2677_out0;
wire  [23:0] v$MUX2_2678_out0;
wire  [23:0] v$MUX2_2679_out0;
wire  [23:0] v$MUX2_2680_out0;
wire  [23:0] v$MUX2_2681_out0;
wire  [23:0] v$MUX2_2688_out0;
wire  [23:0] v$MUX2_2689_out0;
wire  [23:0] v$MUX2_2690_out0;
wire  [23:0] v$MUX2_2691_out0;
wire  [23:0] v$MUX2_2692_out0;
wire  [23:0] v$MUX2_2693_out0;
wire  [23:0] v$MUX2_2694_out0;
wire  [23:0] v$MUX2_2695_out0;
wire  [23:0] v$MUX2_2696_out0;
wire  [23:0] v$MUX2_2697_out0;
wire  [23:0] v$MUX2_2698_out0;
wire  [23:0] v$MUX2_2699_out0;
wire  [23:0] v$MUX2_2700_out0;
wire  [23:0] v$MUX2_2701_out0;
wire  [23:0] v$MUX2_2702_out0;
wire  [23:0] v$MUX2_2703_out0;
wire  [23:0] v$MUX2_2704_out0;
wire  [23:0] v$MUX2_2705_out0;
wire  [23:0] v$MUX2_2706_out0;
wire  [23:0] v$MUX2_2707_out0;
wire  [23:0] v$MUX3_13369_out0;
wire  [23:0] v$MUX3_13370_out0;
wire  [23:0] v$MUX3_18515_out0;
wire  [23:0] v$MUX3_18516_out0;
wire  [23:0] v$MUX3_3320_out0;
wire  [23:0] v$MUX3_3321_out0;
wire  [23:0] v$MUX3_3953_out0;
wire  [23:0] v$MUX3_3954_out0;
wire  [23:0] v$MUX4_6167_out0;
wire  [23:0] v$MUX4_6168_out0;
wire  [23:0] v$MUX4_8416_out0;
wire  [23:0] v$MUX4_8417_out0;
wire  [23:0] v$MUX5_10765_out0;
wire  [23:0] v$MUX5_10766_out0;
wire  [23:0] v$MUX5_1767_out0;
wire  [23:0] v$MUX5_1768_out0;
wire  [23:0] v$MUX5_6486_out0;
wire  [23:0] v$MUX5_6487_out0;
wire  [23:0] v$MUX7_3505_out0;
wire  [23:0] v$MUX7_3506_out0;
wire  [23:0] v$MUX8_5638_out0;
wire  [23:0] v$MUX8_5639_out0;
wire  [23:0] v$MUX9_2652_out0;
wire  [23:0] v$MUX9_2653_out0;
wire  [23:0] v$OP1$MANTISA$ADDER_3834_out0;
wire  [23:0] v$OP1$MANTISA$ADDER_3835_out0;
wire  [23:0] v$OP1$MANTISA$MULTIPLY_12460_out0;
wire  [23:0] v$OP1$MANTISA$MULTIPLY_12461_out0;
wire  [23:0] v$OP1$MANTISA_12378_out0;
wire  [23:0] v$OP1$MANTISA_12379_out0;
wire  [23:0] v$OP1$MANTISA_3971_out0;
wire  [23:0] v$OP1$MANTISA_3972_out0;
wire  [23:0] v$OP1$MANTISA_9449_out0;
wire  [23:0] v$OP1$MANTISA_9450_out0;
wire  [23:0] v$OP1_4258_out0;
wire  [23:0] v$OP1_4259_out0;
wire  [23:0] v$OP2$MANTISA$ADDER_7808_out0;
wire  [23:0] v$OP2$MANTISA$ADDER_7809_out0;
wire  [23:0] v$OP2$MANTISA$MULTIPLY_2656_out0;
wire  [23:0] v$OP2$MANTISA$MULTIPLY_2657_out0;
wire  [23:0] v$OP2$MANTISA_2853_out0;
wire  [23:0] v$OP2$MANTISA_2854_out0;
wire  [23:0] v$OP2$MANTISA_3710_out0;
wire  [23:0] v$OP2$MANTISA_3711_out0;
wire  [23:0] v$OP2$MANTISA_9922_out0;
wire  [23:0] v$OP2$MANTISA_9923_out0;
wire  [23:0] v$OP2_13046_out0;
wire  [23:0] v$OP2_13047_out0;
wire  [23:0] v$OP2_4320_out0;
wire  [23:0] v$OP2_4321_out0;
wire  [23:0] v$OP2_5076_out0;
wire  [23:0] v$OP2_5077_out0;
wire  [23:0] v$OUT_10436_out0;
wire  [23:0] v$OUT_10437_out0;
wire  [23:0] v$OUT_10438_out0;
wire  [23:0] v$OUT_10439_out0;
wire  [23:0] v$OUT_10440_out0;
wire  [23:0] v$OUT_10441_out0;
wire  [23:0] v$OUT_10442_out0;
wire  [23:0] v$OUT_10443_out0;
wire  [23:0] v$OUT_15515_out0;
wire  [23:0] v$OUT_15516_out0;
wire  [23:0] v$OUT_15517_out0;
wire  [23:0] v$OUT_15518_out0;
wire  [23:0] v$OUT_15519_out0;
wire  [23:0] v$OUT_15520_out0;
wire  [23:0] v$OUT_15521_out0;
wire  [23:0] v$OUT_15522_out0;
wire  [23:0] v$OUT_15523_out0;
wire  [23:0] v$OUT_15524_out0;
wire  [23:0] v$OUT_15525_out0;
wire  [23:0] v$OUT_15526_out0;
wire  [23:0] v$OUT_15527_out0;
wire  [23:0] v$OUT_15528_out0;
wire  [23:0] v$OUT_15529_out0;
wire  [23:0] v$OUT_15530_out0;
wire  [23:0] v$OUT_15531_out0;
wire  [23:0] v$OUT_15532_out0;
wire  [23:0] v$OUT_15533_out0;
wire  [23:0] v$OUT_15534_out0;
wire  [23:0] v$OUT_15535_out0;
wire  [23:0] v$OUT_15536_out0;
wire  [23:0] v$OUT_15537_out0;
wire  [23:0] v$OUT_15538_out0;
wire  [23:0] v$OUT_15539_out0;
wire  [23:0] v$OUT_15540_out0;
wire  [23:0] v$OUT_15541_out0;
wire  [23:0] v$OUT_15542_out0;
wire  [23:0] v$OUT_15543_out0;
wire  [23:0] v$OUT_15544_out0;
wire  [23:0] v$OUT_15545_out0;
wire  [23:0] v$OUT_15546_out0;
wire  [23:0] v$OUT_15547_out0;
wire  [23:0] v$OUT_15548_out0;
wire  [23:0] v$OUT_15549_out0;
wire  [23:0] v$OUT_15550_out0;
wire  [23:0] v$OUT_15551_out0;
wire  [23:0] v$OUT_15552_out0;
wire  [23:0] v$OUT_15553_out0;
wire  [23:0] v$OUT_15554_out0;
wire  [23:0] v$OUT_15555_out0;
wire  [23:0] v$OUT_15556_out0;
wire  [23:0] v$OUT_15557_out0;
wire  [23:0] v$OUT_15558_out0;
wire  [23:0] v$OUT_15559_out0;
wire  [23:0] v$OUT_15560_out0;
wire  [23:0] v$OUT_15561_out0;
wire  [23:0] v$OUT_15562_out0;
wire  [23:0] v$OUT_15563_out0;
wire  [23:0] v$OUT_15564_out0;
wire  [23:0] v$OUT_15565_out0;
wire  [23:0] v$OUT_15566_out0;
wire  [23:0] v$OUT_15567_out0;
wire  [23:0] v$OUT_15568_out0;
wire  [23:0] v$OUT_15569_out0;
wire  [23:0] v$OUT_15570_out0;
wire  [23:0] v$OUT_15571_out0;
wire  [23:0] v$OUT_15572_out0;
wire  [23:0] v$OUT_15573_out0;
wire  [23:0] v$OUT_15574_out0;
wire  [23:0] v$OUT_15575_out0;
wire  [23:0] v$OUT_15576_out0;
wire  [23:0] v$OUT_5128_out0;
wire  [23:0] v$OUT_5129_out0;
wire  [23:0] v$OUT_5130_out0;
wire  [23:0] v$OUT_5131_out0;
wire  [23:0] v$RESULT_5279_out0;
wire  [23:0] v$RESULT_5280_out0;
wire  [23:0] v$SUM1_13397_out0;
wire  [23:0] v$SUM1_13398_out0;
wire  [23:0] v$SUM1_13399_out0;
wire  [23:0] v$SUM1_13400_out0;
wire  [23:0] v$SUM1_13401_out0;
wire  [23:0] v$SUM1_13402_out0;
wire  [23:0] v$SUM_2068_out0;
wire  [23:0] v$SUM_2069_out0;
wire  [23:0] v$SUM_9731_out0;
wire  [23:0] v$SUM_9732_out0;
wire  [23:0] v$SUM_9733_out0;
wire  [23:0] v$SUM_9734_out0;
wire  [23:0] v$SUM_9735_out0;
wire  [23:0] v$SUM_9736_out0;
wire  [23:0] v$XOR$IN_2450_out0;
wire  [23:0] v$XOR$IN_2451_out0;
wire  [23:0] v$XOR1_5640_out0;
wire  [23:0] v$XOR1_5641_out0;
wire  [23:0] v$XOR2_8172_out0;
wire  [23:0] v$XOR2_8173_out0;
wire  [23:0] v$_10327_out0;
wire  [23:0] v$_10328_out0;
wire  [23:0] v$_10329_out0;
wire  [23:0] v$_10330_out0;
wire  [23:0] v$_10331_out0;
wire  [23:0] v$_10332_out0;
wire  [23:0] v$_10464_out0;
wire  [23:0] v$_10465_out0;
wire  [23:0] v$_11523_out0;
wire  [23:0] v$_11524_out0;
wire  [23:0] v$_1303_out0;
wire  [23:0] v$_1304_out0;
wire  [23:0] v$_14703_out0;
wire  [23:0] v$_14704_out0;
wire  [23:0] v$_15937_out0;
wire  [23:0] v$_15938_out0;
wire  [23:0] v$_1665_out0;
wire  [23:0] v$_1666_out0;
wire  [23:0] v$_18382_out0;
wire  [23:0] v$_18383_out0;
wire  [23:0] v$_3939_out0;
wire  [23:0] v$_3940_out0;
wire  [23:0] v$_3941_out0;
wire  [23:0] v$_3942_out0;
wire  [23:0] v$_3943_out0;
wire  [23:0] v$_3944_out0;
wire  [23:0] v$_4406_out0;
wire  [23:0] v$_4407_out0;
wire  [23:0] v$_4408_out0;
wire  [23:0] v$_4409_out0;
wire  [23:0] v$_4410_out0;
wire  [23:0] v$_4411_out0;
wire  [23:0] v$_4412_out0;
wire  [23:0] v$_4413_out0;
wire  [23:0] v$_4414_out0;
wire  [23:0] v$_4415_out0;
wire  [23:0] v$_4416_out0;
wire  [23:0] v$_4417_out0;
wire  [23:0] v$_4418_out0;
wire  [23:0] v$_4419_out0;
wire  [23:0] v$_4420_out0;
wire  [23:0] v$_4421_out0;
wire  [23:0] v$_4422_out0;
wire  [23:0] v$_4423_out0;
wire  [23:0] v$_4424_out0;
wire  [23:0] v$_4425_out0;
wire  [23:0] v$_4426_out0;
wire  [23:0] v$_4427_out0;
wire  [23:0] v$_4428_out0;
wire  [23:0] v$_4429_out0;
wire  [23:0] v$_4430_out0;
wire  [23:0] v$_4431_out0;
wire  [23:0] v$_4432_out0;
wire  [23:0] v$_4433_out0;
wire  [23:0] v$_4434_out0;
wire  [23:0] v$_4435_out0;
wire  [23:0] v$_4436_out0;
wire  [23:0] v$_4437_out0;
wire  [23:0] v$_4438_out0;
wire  [23:0] v$_4439_out0;
wire  [23:0] v$_4440_out0;
wire  [23:0] v$_4441_out0;
wire  [23:0] v$_4442_out0;
wire  [23:0] v$_4443_out0;
wire  [23:0] v$_4444_out0;
wire  [23:0] v$_4445_out0;
wire  [23:0] v$_4446_out0;
wire  [23:0] v$_4447_out0;
wire  [23:0] v$_4448_out0;
wire  [23:0] v$_4449_out0;
wire  [23:0] v$_4450_out0;
wire  [23:0] v$_4451_out0;
wire  [23:0] v$_4452_out0;
wire  [23:0] v$_4453_out0;
wire  [23:0] v$_4454_out0;
wire  [23:0] v$_4455_out0;
wire  [23:0] v$_4456_out0;
wire  [23:0] v$_4457_out0;
wire  [23:0] v$_4458_out0;
wire  [23:0] v$_4459_out0;
wire  [23:0] v$_4460_out0;
wire  [23:0] v$_4461_out0;
wire  [23:0] v$_4462_out0;
wire  [23:0] v$_4463_out0;
wire  [23:0] v$_4464_out0;
wire  [23:0] v$_4465_out0;
wire  [23:0] v$_4466_out0;
wire  [23:0] v$_4467_out0;
wire  [23:0] v$_7693_out0;
wire  [23:0] v$_7694_out0;
wire  [23:0] v$_7735_out0;
wire  [23:0] v$_7736_out0;
wire  [23:0] v$_7943_out0;
wire  [23:0] v$_7944_out0;
wire  [23:0] v$_9307_out0;
wire  [23:0] v$_9308_out0;
wire  [23:0] v$_9309_out0;
wire  [23:0] v$_9310_out0;
wire  [23:0] v$_9311_out0;
wire  [23:0] v$_9312_out0;
wire  [23:0] v$_9313_out0;
wire  [23:0] v$_9314_out0;
wire  [23:0] v$_9315_out0;
wire  [23:0] v$_9316_out0;
wire  [23:0] v$_9317_out0;
wire  [23:0] v$_9318_out0;
wire  [23:0] v$_9319_out0;
wire  [23:0] v$_9320_out0;
wire  [23:0] v$_9321_out0;
wire  [23:0] v$_9322_out0;
wire  [23:0] v$_9323_out0;
wire  [23:0] v$_9324_out0;
wire  [23:0] v$_9325_out0;
wire  [23:0] v$_9326_out0;
wire  [23:0] v$_9327_out0;
wire  [23:0] v$_9328_out0;
wire  [23:0] v$_9329_out0;
wire  [23:0] v$_9330_out0;
wire  [23:0] v$_9331_out0;
wire  [23:0] v$_9332_out0;
wire  [23:0] v$_9333_out0;
wire  [23:0] v$_9334_out0;
wire  [23:0] v$_9335_out0;
wire  [23:0] v$_9336_out0;
wire  [23:0] v$_9337_out0;
wire  [23:0] v$_9338_out0;
wire  [23:0] v$_9339_out0;
wire  [23:0] v$_9340_out0;
wire  [23:0] v$_9341_out0;
wire  [23:0] v$_9342_out0;
wire  [23:0] v$_9343_out0;
wire  [23:0] v$_9344_out0;
wire  [23:0] v$_9345_out0;
wire  [23:0] v$_9346_out0;
wire  [23:0] v$_9347_out0;
wire  [23:0] v$_9348_out0;
wire  [23:0] v$_9349_out0;
wire  [23:0] v$_9350_out0;
wire  [23:0] v$_9351_out0;
wire  [23:0] v$_9352_out0;
wire  [23:0] v$_9353_out0;
wire  [23:0] v$_9354_out0;
wire  [23:0] v$_9355_out0;
wire  [23:0] v$_9356_out0;
wire  [23:0] v$_9357_out0;
wire  [23:0] v$_9358_out0;
wire  [23:0] v$_9359_out0;
wire  [23:0] v$_9360_out0;
wire  [23:0] v$_9361_out0;
wire  [23:0] v$_9362_out0;
wire  [23:0] v$_9363_out0;
wire  [23:0] v$_9364_out0;
wire  [23:0] v$_9365_out0;
wire  [23:0] v$_9366_out0;
wire  [23:0] v$_9367_out0;
wire  [23:0] v$_9368_out0;
wire  [27:0] v$_10354_out0;
wire  [27:0] v$_10355_out0;
wire  [2:0] v$9_14775_out0;
wire  [2:0] v$9_14776_out0;
wire  [2:0] v$ALU$OP_17437_out0;
wire  [2:0] v$ALU$OP_17438_out0;
wire  [2:0] v$C10_14117_out0;
wire  [2:0] v$C10_14118_out0;
wire  [2:0] v$C1_17454_out0;
wire  [2:0] v$C1_17455_out0;
wire  [2:0] v$C2_13910_out0;
wire  [2:0] v$C2_13911_out0;
wire  [2:0] v$C4_6859_out0;
wire  [2:0] v$C4_6860_out0;
wire  [2:0] v$IR1$OP_5761_out0;
wire  [2:0] v$IR1$OP_5762_out0;
wire  [2:0] v$IR2$OP_16464_out0;
wire  [2:0] v$IR2$OP_16465_out0;
wire  [2:0] v$IR2$OP_18625_out0;
wire  [2:0] v$IR2$OP_18626_out0;
wire  [2:0] v$MODE_1773_out0;
wire  [2:0] v$MODE_1774_out0;
wire  [2:0] v$MODE_9454_out0;
wire  [2:0] v$MODE_9455_out0;
wire  [2:0] v$MUX1_15297_out0;
wire  [2:0] v$MUX1_15298_out0;
wire  [2:0] v$MUX1_15299_out0;
wire  [2:0] v$MUX1_15300_out0;
wire  [2:0] v$MUX1_15301_out0;
wire  [2:0] v$MUX1_15302_out0;
wire  [2:0] v$MUX1_15303_out0;
wire  [2:0] v$MUX1_15304_out0;
wire  [2:0] v$MUX1_15305_out0;
wire  [2:0] v$MUX1_15306_out0;
wire  [2:0] v$Mode_11483_out0;
wire  [2:0] v$Mode_11484_out0;
wire  [2:0] v$Mode_13777_out0;
wire  [2:0] v$Mode_13778_out0;
wire  [2:0] v$NUPPER_18007_out0;
wire  [2:0] v$NUPPER_18008_out0;
wire  [2:0] v$NUPPER_18009_out0;
wire  [2:0] v$NUPPER_18010_out0;
wire  [2:0] v$OPCODE_8218_out0;
wire  [2:0] v$OPCODE_8219_out0;
wire  [2:0] v$OP_18253_out0;
wire  [2:0] v$OP_18254_out0;
wire  [2:0] v$OP_2034_out0;
wire  [2:0] v$OP_2035_out0;
wire  [2:0] v$SEL26_5050_out0;
wire  [2:0] v$SEL26_5051_out0;
wire  [2:0] v$SEL26_5052_out0;
wire  [2:0] v$SEL26_5053_out0;
wire  [2:0] v$Y_8074_out0;
wire  [2:0] v$Y_8075_out0;
wire  [2:0] v$Y_8076_out0;
wire  [2:0] v$Y_8077_out0;
wire  [2:0] v$Y_8078_out0;
wire  [2:0] v$Y_8079_out0;
wire  [2:0] v$Y_8080_out0;
wire  [2:0] v$Y_8081_out0;
wire  [2:0] v$Y_8082_out0;
wire  [2:0] v$Y_8083_out0;
wire  [2:0] v$_10356_out0;
wire  [2:0] v$_10356_out1;
wire  [2:0] v$_10357_out0;
wire  [2:0] v$_10357_out1;
wire  [2:0] v$_10358_out0;
wire  [2:0] v$_10358_out1;
wire  [2:0] v$_10359_out0;
wire  [2:0] v$_10359_out1;
wire  [2:0] v$_10360_out0;
wire  [2:0] v$_10360_out1;
wire  [2:0] v$_10361_out0;
wire  [2:0] v$_10361_out1;
wire  [2:0] v$_10474_out0;
wire  [2:0] v$_10474_out1;
wire  [2:0] v$_10475_out0;
wire  [2:0] v$_10475_out1;
wire  [2:0] v$_10476_out0;
wire  [2:0] v$_10476_out1;
wire  [2:0] v$_10477_out0;
wire  [2:0] v$_10477_out1;
wire  [2:0] v$_10478_out0;
wire  [2:0] v$_10478_out1;
wire  [2:0] v$_10479_out0;
wire  [2:0] v$_10479_out1;
wire  [2:0] v$_13561_out0;
wire  [2:0] v$_13561_out1;
wire  [2:0] v$_13562_out0;
wire  [2:0] v$_13562_out1;
wire  [2:0] v$_13563_out0;
wire  [2:0] v$_13563_out1;
wire  [2:0] v$_13564_out0;
wire  [2:0] v$_13564_out1;
wire  [2:0] v$_13565_out0;
wire  [2:0] v$_13565_out1;
wire  [2:0] v$_13566_out0;
wire  [2:0] v$_13566_out1;
wire  [2:0] v$_14324_out0;
wire  [2:0] v$_14324_out1;
wire  [2:0] v$_14325_out0;
wire  [2:0] v$_14325_out1;
wire  [2:0] v$_14326_out0;
wire  [2:0] v$_14326_out1;
wire  [2:0] v$_14327_out0;
wire  [2:0] v$_14327_out1;
wire  [2:0] v$_14328_out0;
wire  [2:0] v$_14328_out1;
wire  [2:0] v$_14329_out0;
wire  [2:0] v$_14329_out1;
wire  [2:0] v$_14355_out0;
wire  [2:0] v$_14355_out1;
wire  [2:0] v$_14356_out0;
wire  [2:0] v$_14356_out1;
wire  [2:0] v$_14357_out0;
wire  [2:0] v$_14357_out1;
wire  [2:0] v$_14358_out0;
wire  [2:0] v$_14358_out1;
wire  [2:0] v$_14359_out0;
wire  [2:0] v$_14359_out1;
wire  [2:0] v$_14360_out0;
wire  [2:0] v$_14360_out1;
wire  [2:0] v$_17304_out0;
wire  [2:0] v$_17305_out0;
wire  [2:0] v$_18340_out0;
wire  [2:0] v$_18340_out1;
wire  [2:0] v$_18341_out0;
wire  [2:0] v$_18341_out1;
wire  [2:0] v$_18342_out0;
wire  [2:0] v$_18342_out1;
wire  [2:0] v$_18343_out0;
wire  [2:0] v$_18343_out1;
wire  [2:0] v$_18344_out0;
wire  [2:0] v$_18344_out1;
wire  [2:0] v$_18345_out0;
wire  [2:0] v$_18345_out1;
wire  [2:0] v$_19027_out0;
wire  [2:0] v$_19027_out1;
wire  [2:0] v$_19028_out0;
wire  [2:0] v$_19028_out1;
wire  [2:0] v$_19029_out0;
wire  [2:0] v$_19029_out1;
wire  [2:0] v$_19030_out0;
wire  [2:0] v$_19030_out1;
wire  [2:0] v$_19031_out0;
wire  [2:0] v$_19031_out1;
wire  [2:0] v$_19032_out0;
wire  [2:0] v$_19032_out1;
wire  [2:0] v$_19155_out0;
wire  [2:0] v$_19156_out0;
wire  [2:0] v$_2024_out0;
wire  [2:0] v$_2024_out1;
wire  [2:0] v$_2025_out0;
wire  [2:0] v$_2025_out1;
wire  [2:0] v$_2026_out0;
wire  [2:0] v$_2026_out1;
wire  [2:0] v$_2027_out0;
wire  [2:0] v$_2027_out1;
wire  [2:0] v$_2028_out0;
wire  [2:0] v$_2028_out1;
wire  [2:0] v$_2029_out0;
wire  [2:0] v$_2029_out1;
wire  [2:0] v$_5112_out0;
wire  [2:0] v$_5113_out0;
wire  [2:0] v$_5212_out0;
wire  [2:0] v$_5213_out0;
wire  [2:0] v$_5705_out0;
wire  [2:0] v$_5706_out0;
wire  [2:0] v$_5707_out0;
wire  [2:0] v$_5708_out0;
wire  [2:0] v$_5709_out0;
wire  [2:0] v$_5710_out0;
wire  [2:0] v$_5711_out0;
wire  [2:0] v$_5712_out0;
wire  [2:0] v$_5713_out0;
wire  [2:0] v$_5714_out0;
wire  [2:0] v$_8414_out0;
wire  [2:0] v$_8415_out0;
wire  [2:0] v$_8453_out0;
wire  [2:0] v$_8454_out0;
wire  [2:0] v$_8455_out0;
wire  [2:0] v$_8456_out0;
wire  [2:0] v$_8457_out0;
wire  [2:0] v$_8458_out0;
wire  [2:0] v$_8459_out0;
wire  [2:0] v$_8460_out0;
wire  [2:0] v$_8461_out0;
wire  [2:0] v$_8462_out0;
wire  [30:0] v$C4_8567_out0;
wire  [30:0] v$C4_8569_out0;
wire  [30:0] v$MUX12_15750_out0;
wire  [30:0] v$MUX12_15751_out0;
wire  [30:0] v$MUX2_14209_out0;
wire  [30:0] v$MUX2_14211_out0;
wire  [30:0] v$MUX6_18078_out0;
wire  [30:0] v$MUX6_18079_out0;
wire  [30:0] v$SINGLE$MERGE_12686_out0;
wire  [30:0] v$SINGLE$MERGE_12687_out0;
wire  [30:0] v$_12403_out0;
wire  [30:0] v$_12404_out0;
wire  [30:0] v$_15939_out0;
wire  [30:0] v$_15940_out0;
wire  [30:0] v$_16451_out0;
wire  [30:0] v$_16453_out0;
wire  [30:0] v$_58_out0;
wire  [30:0] v$_59_out0;
wire  [30:0] v$_7305_out0;
wire  [30:0] v$_7306_out0;
wire  [31:0] v$A$32$BIT$MUL_3965_out0;
wire  [31:0] v$A$32$BIT$MUL_3966_out0;
wire  [31:0] v$A$32$BIT_17442_out0;
wire  [31:0] v$A$32$BIT_17443_out0;
wire  [31:0] v$A$32BIT_3201_out0;
wire  [31:0] v$A$32BIT_3202_out0;
wire  [31:0] v$A$FPU$ADDER$32$BIT_16490_out0;
wire  [31:0] v$A$FPU$ADDER$32$BIT_16491_out0;
wire  [31:0] v$A_14400_out0;
wire  [31:0] v$A_14402_out0;
wire  [31:0] v$A_14404_out0;
wire  [31:0] v$A_14406_out0;
wire  [31:0] v$B$32$BIT$FPU$ADDER_10641_out0;
wire  [31:0] v$B$32$BIT$FPU$ADDER_10642_out0;
wire  [31:0] v$B$32$BIT_18291_out0;
wire  [31:0] v$B$32$BIT_18292_out0;
wire  [31:0] v$B$32$MUL_13837_out0;
wire  [31:0] v$B$32$MUL_13838_out0;
wire  [31:0] v$B$32BIT_19081_out0;
wire  [31:0] v$B$32BIT_19082_out0;
wire  [31:0] v$B_5039_out0;
wire  [31:0] v$B_5041_out0;
wire  [31:0] v$B_5043_out0;
wire  [31:0] v$B_5045_out0;
wire  [31:0] v$C1_15809_out0;
wire  [31:0] v$C1_15810_out0;
wire  [31:0] v$C4_14636_out0;
wire  [31:0] v$C4_14637_out0;
wire  [31:0] v$C5_4269_out0;
wire  [31:0] v$C5_4270_out0;
wire  [31:0] v$FPU$ADDER$OUT_4166_out0;
wire  [31:0] v$FPU$ADDER$OUT_4167_out0;
wire  [31:0] v$FPU$ADDER$OUT_6072_out0;
wire  [31:0] v$FPU$ADDER$OUT_6073_out0;
wire  [31:0] v$FPU$MULTIPLIER$OUT_11425_out0;
wire  [31:0] v$FPU$MULTIPLIER$OUT_11426_out0;
wire  [31:0] v$HALF$PRECISION$32$BIT_15410_out0;
wire  [31:0] v$HALF$PRECISION$32$BIT_15411_out0;
wire  [31:0] v$HALF$PRECISION_10767_out0;
wire  [31:0] v$HALF$PRECISION_10768_out0;
wire  [31:0] v$MUX12_17418_out0;
wire  [31:0] v$MUX12_17419_out0;
wire  [31:0] v$MUX13_11226_out0;
wire  [31:0] v$MUX13_11227_out0;
wire  [31:0] v$MUX14_1335_out0;
wire  [31:0] v$MUX14_1336_out0;
wire  [31:0] v$MUX1_14132_out0;
wire  [31:0] v$MUX1_14133_out0;
wire  [31:0] v$MUX2_16839_out0;
wire  [31:0] v$MUX2_16840_out0;
wire  [31:0] v$MUX3_9291_out0;
wire  [31:0] v$MUX3_9292_out0;
wire  [31:0] v$MUX4_1411_out0;
wire  [31:0] v$MUX4_1412_out0;
wire  [31:0] v$MUX7_5078_out0;
wire  [31:0] v$MUX7_5079_out0;
wire  [31:0] v$OUT1_18415_out0;
wire  [31:0] v$OUT1_18416_out0;
wire  [31:0] v$OUT_13073_out0;
wire  [31:0] v$OUT_13075_out0;
wire  [31:0] v$OUT_3588_out0;
wire  [31:0] v$OUT_3589_out0;
wire  [31:0] v$SINGLE$PRECISION$32$BITS_14286_out0;
wire  [31:0] v$SINGLE$PRECISION$32$BITS_14287_out0;
wire  [31:0] v$SINGLE$PRECISION_8227_out0;
wire  [31:0] v$SINGLE$PRECISION_8228_out0;
wire  [31:0] v$_13118_out0;
wire  [31:0] v$_13119_out0;
wire  [31:0] v$_16430_out0;
wire  [31:0] v$_16431_out0;
wire  [31:0] v$_17132_out0;
wire  [31:0] v$_17133_out0;
wire  [31:0] v$_17422_out0;
wire  [31:0] v$_17423_out0;
wire  [31:0] v$_17630_out0;
wire  [31:0] v$_17631_out0;
wire  [31:0] v$_18862_out0;
wire  [31:0] v$_18863_out0;
wire  [31:0] v$_19024_out0;
wire  [31:0] v$_19026_out0;
wire  [31:0] v$_2012_out0;
wire  [31:0] v$_2013_out0;
wire  [3:0] v$3_13980_out0;
wire  [3:0] v$3_13981_out0;
wire  [3:0] v$9_14918_out0;
wire  [3:0] v$9_14919_out0;
wire  [3:0] v$ADDRMSB_15646_out0;
wire  [3:0] v$ADDRMSB_15647_out0;
wire  [3:0] v$A_11856_out0;
wire  [3:0] v$A_11858_out0;
wire  [3:0] v$A_11859_out0;
wire  [3:0] v$A_11860_out0;
wire  [3:0] v$A_11862_out0;
wire  [3:0] v$A_11863_out0;
wire  [3:0] v$A_11866_out0;
wire  [3:0] v$A_11867_out0;
wire  [3:0] v$A_11870_out0;
wire  [3:0] v$A_11871_out0;
wire  [3:0] v$A_11872_out0;
wire  [3:0] v$A_11874_out0;
wire  [3:0] v$A_11875_out0;
wire  [3:0] v$A_11876_out0;
wire  [3:0] v$A_11878_out0;
wire  [3:0] v$A_11879_out0;
wire  [3:0] v$A_11882_out0;
wire  [3:0] v$A_11883_out0;
wire  [3:0] v$A_11886_out0;
wire  [3:0] v$A_11887_out0;
wire  [3:0] v$B_13793_out0;
wire  [3:0] v$B_13794_out0;
wire  [3:0] v$B_15028_out0;
wire  [3:0] v$B_15030_out0;
wire  [3:0] v$B_15031_out0;
wire  [3:0] v$B_15032_out0;
wire  [3:0] v$B_15034_out0;
wire  [3:0] v$B_15035_out0;
wire  [3:0] v$B_15038_out0;
wire  [3:0] v$B_15039_out0;
wire  [3:0] v$B_15042_out0;
wire  [3:0] v$B_15043_out0;
wire  [3:0] v$B_15044_out0;
wire  [3:0] v$B_15046_out0;
wire  [3:0] v$B_15047_out0;
wire  [3:0] v$B_15048_out0;
wire  [3:0] v$B_15050_out0;
wire  [3:0] v$B_15051_out0;
wire  [3:0] v$B_15054_out0;
wire  [3:0] v$B_15055_out0;
wire  [3:0] v$B_15058_out0;
wire  [3:0] v$B_15059_out0;
wire  [3:0] v$B_15227_out0;
wire  [3:0] v$B_15228_out0;
wire  [3:0] v$B_3885_out0;
wire  [3:0] v$B_3886_out0;
wire  [3:0] v$B_8628_out0;
wire  [3:0] v$B_8629_out0;
wire  [3:0] v$C0_208_out0;
wire  [3:0] v$C0_209_out0;
wire  [3:0] v$C12_3507_out0;
wire  [3:0] v$C12_3508_out0;
wire  [3:0] v$C1_13395_out0;
wire  [3:0] v$C1_13396_out0;
wire  [3:0] v$C1_5654_out0;
wire  [3:0] v$C1_5655_out0;
wire  [3:0] v$C1_6245_out0;
wire  [3:0] v$C1_6250_out0;
wire  [3:0] v$C1_6255_out0;
wire  [3:0] v$C1_6259_out0;
wire  [3:0] v$C1_6265_out0;
wire  [3:0] v$C1_6269_out0;
wire  [3:0] v$C1_6276_out0;
wire  [3:0] v$C1_6281_out0;
wire  [3:0] v$C1_6286_out0;
wire  [3:0] v$C1_6290_out0;
wire  [3:0] v$C1_6296_out0;
wire  [3:0] v$C1_6300_out0;
wire  [3:0] v$C1_8289_out0;
wire  [3:0] v$C1_8293_out0;
wire  [3:0] v$C2_107_out0;
wire  [3:0] v$C2_112_out0;
wire  [3:0] v$C2_117_out0;
wire  [3:0] v$C2_121_out0;
wire  [3:0] v$C2_127_out0;
wire  [3:0] v$C2_131_out0;
wire  [3:0] v$C2_138_out0;
wire  [3:0] v$C2_143_out0;
wire  [3:0] v$C2_148_out0;
wire  [3:0] v$C2_152_out0;
wire  [3:0] v$C2_158_out0;
wire  [3:0] v$C2_162_out0;
wire  [3:0] v$C4_11272_out0;
wire  [3:0] v$C4_11273_out0;
wire  [3:0] v$C8_7599_out0;
wire  [3:0] v$C8_7600_out0;
wire  [3:0] v$C8_8637_out0;
wire  [3:0] v$C8_8638_out0;
wire  [3:0] v$IN_15677_out0;
wire  [3:0] v$IN_15678_out0;
wire  [3:0] v$IN_15679_out0;
wire  [3:0] v$IN_15680_out0;
wire  [3:0] v$IN_15681_out0;
wire  [3:0] v$IN_15682_out0;
wire  [3:0] v$IN_15683_out0;
wire  [3:0] v$IN_15684_out0;
wire  [3:0] v$IN_15685_out0;
wire  [3:0] v$IN_15686_out0;
wire  [3:0] v$IN_15687_out0;
wire  [3:0] v$IN_15688_out0;
wire  [3:0] v$IN_15689_out0;
wire  [3:0] v$IN_15690_out0;
wire  [3:0] v$IN_15691_out0;
wire  [3:0] v$IN_15692_out0;
wire  [3:0] v$IN_15693_out0;
wire  [3:0] v$IN_15694_out0;
wire  [3:0] v$IN_15695_out0;
wire  [3:0] v$IN_15696_out0;
wire  [3:0] v$IN_15697_out0;
wire  [3:0] v$IN_15698_out0;
wire  [3:0] v$IN_15699_out0;
wire  [3:0] v$IN_15700_out0;
wire  [3:0] v$IN_15701_out0;
wire  [3:0] v$IN_15702_out0;
wire  [3:0] v$IN_15703_out0;
wire  [3:0] v$IN_15704_out0;
wire  [3:0] v$IN_15705_out0;
wire  [3:0] v$IN_15706_out0;
wire  [3:0] v$IN_15707_out0;
wire  [3:0] v$IN_15708_out0;
wire  [3:0] v$IN_15709_out0;
wire  [3:0] v$IN_15710_out0;
wire  [3:0] v$IN_15711_out0;
wire  [3:0] v$IN_15712_out0;
wire  [3:0] v$IR1$FULL$OP$CODE_17650_out0;
wire  [3:0] v$IR1$FULL$OP$CODE_17651_out0;
wire  [3:0] v$IR1$N_16365_out0;
wire  [3:0] v$IR1$N_16366_out0;
wire  [3:0] v$IR1$OPCODE_3102_out0;
wire  [3:0] v$IR1$OPCODE_3103_out0;
wire  [3:0] v$IR1$OPCODE_9944_out0;
wire  [3:0] v$IR1$OPCODE_9945_out0;
wire  [3:0] v$IR2$FULL$OP$CODE_12392_out0;
wire  [3:0] v$IR2$FULL$OP$CODE_12393_out0;
wire  [3:0] v$IR2$N_3195_out0;
wire  [3:0] v$IR2$N_3196_out0;
wire  [3:0] v$IR2$OPCODE_2761_out0;
wire  [3:0] v$IR2$OPCODE_2762_out0;
wire  [3:0] v$LSBS_15901_out0;
wire  [3:0] v$LSBS_15902_out0;
wire  [3:0] v$MUX3_18114_out0;
wire  [3:0] v$MUX3_18115_out0;
wire  [3:0] v$MUX3_18116_out0;
wire  [3:0] v$MUX3_18117_out0;
wire  [3:0] v$MUX4_3084_out0;
wire  [3:0] v$MUX4_3085_out0;
wire  [3:0] v$MUX4_3086_out0;
wire  [3:0] v$MUX4_3087_out0;
wire  [3:0] v$MUX5_15088_out0;
wire  [3:0] v$MUX5_15089_out0;
wire  [3:0] v$MUX5_4213_out0;
wire  [3:0] v$MUX5_4215_out0;
wire  [3:0] v$MUX5_4217_out0;
wire  [3:0] v$MUX5_4219_out0;
wire  [3:0] v$MUX6_3072_out0;
wire  [3:0] v$MUX6_3073_out0;
wire  [3:0] v$OPCODE_18655_out0;
wire  [3:0] v$OPCODE_18656_out0;
wire  [3:0] v$OP_11500_out0;
wire  [3:0] v$OP_11501_out0;
wire  [3:0] v$OP_15388_out0;
wire  [3:0] v$OP_15389_out0;
wire  [3:0] v$OP_18409_out0;
wire  [3:0] v$OP_18410_out0;
wire  [3:0] v$OP_3869_out0;
wire  [3:0] v$OP_3870_out0;
wire  [3:0] v$OP_5253_out0;
wire  [3:0] v$OP_5254_out0;
wire  [3:0] v$OUT_9282_out0;
wire  [3:0] v$OUT_9284_out0;
wire  [3:0] v$OUT_9286_out0;
wire  [3:0] v$OUT_9288_out0;
wire  [3:0] v$QP_19149_out0;
wire  [3:0] v$QP_19150_out0;
wire  [3:0] v$Q_13552_out0;
wire  [3:0] v$Q_13553_out0;
wire  [3:0] v$Q_6418_out0;
wire  [3:0] v$Q_6419_out0;
wire  [3:0] v$RXFSMQP_10456_out0;
wire  [3:0] v$RXFSMQP_10457_out0;
wire  [3:0] v$RXFSMQ_11310_out0;
wire  [3:0] v$RXFSMQ_11311_out0;
wire  [3:0] v$SEL12_13371_out0;
wire  [3:0] v$SEL12_13372_out0;
wire  [3:0] v$SEL1_10745_out0;
wire  [3:0] v$SEL1_10746_out0;
wire  [3:0] v$SEL1_10747_out0;
wire  [3:0] v$SEL1_10748_out0;
wire  [3:0] v$SEL1_10749_out0;
wire  [3:0] v$SEL1_10750_out0;
wire  [3:0] v$SEL1_10751_out0;
wire  [3:0] v$SEL1_10752_out0;
wire  [3:0] v$SEL1_17079_out0;
wire  [3:0] v$SEL1_17080_out0;
wire  [3:0] v$SEL1_17081_out0;
wire  [3:0] v$SEL1_17082_out0;
wire  [3:0] v$SEL1_17083_out0;
wire  [3:0] v$SEL1_17084_out0;
wire  [3:0] v$SEL1_17085_out0;
wire  [3:0] v$SEL1_17086_out0;
wire  [3:0] v$SEL1_17087_out0;
wire  [3:0] v$SEL1_17088_out0;
wire  [3:0] v$SEL1_17307_out0;
wire  [3:0] v$SEL1_17309_out0;
wire  [3:0] v$SEL1_17311_out0;
wire  [3:0] v$SEL1_17313_out0;
wire  [3:0] v$SEL1_18848_out0;
wire  [3:0] v$SEL1_18849_out0;
wire  [3:0] v$SEL1_9141_out0;
wire  [3:0] v$SEL1_9142_out0;
wire  [3:0] v$SEL2_14439_out0;
wire  [3:0] v$SEL2_14440_out0;
wire  [3:0] v$SEL2_14441_out0;
wire  [3:0] v$SEL2_14442_out0;
wire  [3:0] v$SEL2_18082_out0;
wire  [3:0] v$SEL2_18083_out0;
wire  [3:0] v$SEL2_18084_out0;
wire  [3:0] v$SEL2_18085_out0;
wire  [3:0] v$SEL2_18086_out0;
wire  [3:0] v$SEL2_18087_out0;
wire  [3:0] v$SEL2_18088_out0;
wire  [3:0] v$SEL2_18089_out0;
wire  [3:0] v$SEL2_2628_out0;
wire  [3:0] v$SEL2_2629_out0;
wire  [3:0] v$SEL2_3235_out0;
wire  [3:0] v$SEL2_3236_out0;
wire  [3:0] v$SEL2_3237_out0;
wire  [3:0] v$SEL2_3238_out0;
wire  [3:0] v$SEL2_3239_out0;
wire  [3:0] v$SEL2_3240_out0;
wire  [3:0] v$SEL2_3241_out0;
wire  [3:0] v$SEL2_3242_out0;
wire  [3:0] v$SEL2_3243_out0;
wire  [3:0] v$SEL2_3244_out0;
wire  [3:0] v$SEL3_17270_out0;
wire  [3:0] v$SEL3_17271_out0;
wire  [3:0] v$SEL3_19229_out0;
wire  [3:0] v$SEL3_19230_out0;
wire  [3:0] v$SEL3_19231_out0;
wire  [3:0] v$SEL3_19232_out0;
wire  [3:0] v$SEL3_7683_out0;
wire  [3:0] v$SEL3_7684_out0;
wire  [3:0] v$SEL3_7685_out0;
wire  [3:0] v$SEL3_7686_out0;
wire  [3:0] v$SEL3_9373_out0;
wire  [3:0] v$SEL3_9374_out0;
wire  [3:0] v$SEL3_9375_out0;
wire  [3:0] v$SEL3_9376_out0;
wire  [3:0] v$SEL3_9377_out0;
wire  [3:0] v$SEL3_9378_out0;
wire  [3:0] v$SEL3_9379_out0;
wire  [3:0] v$SEL3_9380_out0;
wire  [3:0] v$SEL4_17971_out0;
wire  [3:0] v$SEL4_17972_out0;
wire  [3:0] v$SEL4_17973_out0;
wire  [3:0] v$SEL4_17974_out0;
wire  [3:0] v$SEL4_17975_out0;
wire  [3:0] v$SEL4_17976_out0;
wire  [3:0] v$SEL4_17977_out0;
wire  [3:0] v$SEL4_17978_out0;
wire  [3:0] v$SEL4_3592_out0;
wire  [3:0] v$SEL4_3593_out0;
wire  [3:0] v$SEL4_3594_out0;
wire  [3:0] v$SEL4_3595_out0;
wire  [3:0] v$SEL4_9954_out0;
wire  [3:0] v$SEL4_9955_out0;
wire  [3:0] v$SEL4_9956_out0;
wire  [3:0] v$SEL4_9957_out0;
wire  [3:0] v$TXFSMQP_9121_out0;
wire  [3:0] v$TXFSMQP_9122_out0;
wire  [3:0] v$TXFSMQ_6469_out0;
wire  [3:0] v$TXFSMQ_6470_out0;
wire  [3:0] v$USELESS_16072_out0;
wire  [3:0] v$_10703_out0;
wire  [3:0] v$_10704_out0;
wire  [3:0] v$_10811_out0;
wire  [3:0] v$_10812_out0;
wire  [3:0] v$_10813_out0;
wire  [3:0] v$_10814_out0;
wire  [3:0] v$_10815_out0;
wire  [3:0] v$_10816_out0;
wire  [3:0] v$_10817_out0;
wire  [3:0] v$_10818_out0;
wire  [3:0] v$_10819_out0;
wire  [3:0] v$_10820_out0;
wire  [3:0] v$_10821_out0;
wire  [3:0] v$_10822_out0;
wire  [3:0] v$_13431_out0;
wire  [3:0] v$_13431_out1;
wire  [3:0] v$_13432_out0;
wire  [3:0] v$_13432_out1;
wire  [3:0] v$_13433_out0;
wire  [3:0] v$_13433_out1;
wire  [3:0] v$_13434_out0;
wire  [3:0] v$_13434_out1;
wire  [3:0] v$_13435_out0;
wire  [3:0] v$_13435_out1;
wire  [3:0] v$_13436_out0;
wire  [3:0] v$_13436_out1;
wire  [3:0] v$_13437_out0;
wire  [3:0] v$_13437_out1;
wire  [3:0] v$_13438_out0;
wire  [3:0] v$_13438_out1;
wire  [3:0] v$_13439_out0;
wire  [3:0] v$_13439_out1;
wire  [3:0] v$_13440_out0;
wire  [3:0] v$_13440_out1;
wire  [3:0] v$_13441_out0;
wire  [3:0] v$_13441_out1;
wire  [3:0] v$_13442_out0;
wire  [3:0] v$_13442_out1;
wire  [3:0] v$_13473_out0;
wire  [3:0] v$_13474_out0;
wire  [3:0] v$_13589_out0;
wire  [3:0] v$_13590_out0;
wire  [3:0] v$_1382_out0;
wire  [3:0] v$_1383_out0;
wire  [3:0] v$_13854_out0;
wire  [3:0] v$_13857_out0;
wire  [3:0] v$_1395_out0;
wire  [3:0] v$_1396_out0;
wire  [3:0] v$_1397_out0;
wire  [3:0] v$_1398_out0;
wire  [3:0] v$_1399_out0;
wire  [3:0] v$_1400_out0;
wire  [3:0] v$_14314_out0;
wire  [3:0] v$_14315_out0;
wire  [3:0] v$_14316_out0;
wire  [3:0] v$_14317_out0;
wire  [3:0] v$_14318_out0;
wire  [3:0] v$_14319_out0;
wire  [3:0] v$_14634_out1;
wire  [3:0] v$_14635_out1;
wire  [3:0] v$_14896_out0;
wire  [3:0] v$_14897_out0;
wire  [3:0] v$_14898_out0;
wire  [3:0] v$_14899_out0;
wire  [3:0] v$_14900_out0;
wire  [3:0] v$_14901_out0;
wire  [3:0] v$_16655_out0;
wire  [3:0] v$_16656_out0;
wire  [3:0] v$_16740_out0;
wire  [3:0] v$_16741_out0;
wire  [3:0] v$_16866_out0;
wire  [3:0] v$_16867_out0;
wire  [3:0] v$_16868_out0;
wire  [3:0] v$_16869_out0;
wire  [3:0] v$_16870_out0;
wire  [3:0] v$_16871_out0;
wire  [3:0] v$_1713_out0;
wire  [3:0] v$_1714_out0;
wire  [3:0] v$_1715_out0;
wire  [3:0] v$_1716_out0;
wire  [3:0] v$_1717_out0;
wire  [3:0] v$_1718_out0;
wire  [3:0] v$_17497_out0;
wire  [3:0] v$_17498_out0;
wire  [3:0] v$_18052_out0;
wire  [3:0] v$_18053_out0;
wire  [3:0] v$_18579_out0;
wire  [3:0] v$_18580_out0;
wire  [3:0] v$_18581_out0;
wire  [3:0] v$_18582_out0;
wire  [3:0] v$_18583_out0;
wire  [3:0] v$_18584_out0;
wire  [3:0] v$_18850_out0;
wire  [3:0] v$_18851_out0;
wire  [3:0] v$_18907_out0;
wire  [3:0] v$_18908_out0;
wire  [3:0] v$_18909_out0;
wire  [3:0] v$_18910_out0;
wire  [3:0] v$_18911_out0;
wire  [3:0] v$_18912_out0;
wire  [3:0] v$_19069_out0;
wire  [3:0] v$_19069_out1;
wire  [3:0] v$_19070_out0;
wire  [3:0] v$_19070_out1;
wire  [3:0] v$_19217_out0;
wire  [3:0] v$_19218_out0;
wire  [3:0] v$_1999_out0;
wire  [3:0] v$_2000_out0;
wire  [3:0] v$_2539_out0;
wire  [3:0] v$_2539_out1;
wire  [3:0] v$_2540_out0;
wire  [3:0] v$_2540_out1;
wire  [3:0] v$_267_out0;
wire  [3:0] v$_268_out0;
wire  [3:0] v$_3104_out0;
wire  [3:0] v$_3104_out1;
wire  [3:0] v$_3105_out0;
wire  [3:0] v$_3105_out1;
wire  [3:0] v$_316_out0;
wire  [3:0] v$_317_out0;
wire  [3:0] v$_3887_out0;
wire  [3:0] v$_3888_out0;
wire  [3:0] v$_3981_out0;
wire  [3:0] v$_3982_out0;
wire  [3:0] v$_4136_out0;
wire  [3:0] v$_4137_out0;
wire  [3:0] v$_4138_out0;
wire  [3:0] v$_4139_out0;
wire  [3:0] v$_4322_out0;
wire  [3:0] v$_4323_out0;
wire  [3:0] v$_5310_out0;
wire  [3:0] v$_5312_out0;
wire  [3:0] v$_5314_out0;
wire  [3:0] v$_5316_out0;
wire  [3:0] v$_5447_out0;
wire  [3:0] v$_5448_out0;
wire  [3:0] v$_5715_out0;
wire  [3:0] v$_5716_out0;
wire  [3:0] v$_5759_out0;
wire  [3:0] v$_5760_out0;
wire  [3:0] v$_6594_out0;
wire  [3:0] v$_6595_out0;
wire  [3:0] v$_6707_out0;
wire  [3:0] v$_6707_out1;
wire  [3:0] v$_6708_out0;
wire  [3:0] v$_6708_out1;
wire  [3:0] v$_7272_out0;
wire  [3:0] v$_7273_out0;
wire  [3:0] v$_7307_out0;
wire  [3:0] v$_7308_out0;
wire  [3:0] v$_746_out0;
wire  [3:0] v$_747_out0;
wire  [3:0] v$_7568_out0;
wire  [3:0] v$_7569_out0;
wire  [3:0] v$_7570_out0;
wire  [3:0] v$_7571_out0;
wire  [3:0] v$_7572_out0;
wire  [3:0] v$_7573_out0;
wire  [3:0] v$_7595_out0;
wire  [3:0] v$_7691_out0;
wire  [3:0] v$_7692_out0;
wire  [3:0] v$_7719_out0;
wire  [3:0] v$_7720_out0;
wire  [3:0] v$_7721_out0;
wire  [3:0] v$_7722_out0;
wire  [3:0] v$_7723_out0;
wire  [3:0] v$_7724_out0;
wire  [3:0] v$_7872_out0;
wire  [3:0] v$_7873_out0;
wire  [3:0] v$_8521_out0;
wire  [3:0] v$_8521_out1;
wire  [3:0] v$_8522_out0;
wire  [3:0] v$_8522_out1;
wire  [3:0] v$_8712_out0;
wire  [3:0] v$_8712_out1;
wire  [3:0] v$_8713_out0;
wire  [3:0] v$_8713_out1;
wire  [3:0] v$_9042_out0;
wire  [3:0] v$_9043_out0;
wire  [3:0] v$_9130_out0;
wire  [3:0] v$_9132_out0;
wire  [3:0] v$_9134_out0;
wire  [3:0] v$_9136_out0;
wire  [3:0] v$_9231_out0;
wire  [3:0] v$_9232_out0;
wire  [3:0] v$_9233_out0;
wire  [3:0] v$_9234_out0;
wire  [3:0] v$_9265_out0;
wire  [3:0] v$_9266_out0;
wire  [3:0] v$_9807_out0;
wire  [3:0] v$_9808_out0;
wire  [3:0] v$_9865_out0;
wire  [3:0] v$_9866_out0;
wire  [3:0] v$_9867_out0;
wire  [3:0] v$_9868_out0;
wire  [3:0] v$_9869_out0;
wire  [3:0] v$_9870_out0;
wire  [43:0] v$AROM1_16768_out0;
wire  [43:0] v$AROM1_16769_out0;
wire  [4:0] v$A$EXP_296_out0;
wire  [4:0] v$A$EXP_298_out0;
wire  [4:0] v$A$EXP_300_out0;
wire  [4:0] v$A$EXP_302_out0;
wire  [4:0] v$A1_12374_out0;
wire  [4:0] v$A1_12375_out0;
wire  [4:0] v$A1_2859_out0;
wire  [4:0] v$A1_2861_out0;
wire  [4:0] v$A1_3146_out0;
wire  [4:0] v$A1_3147_out0;
wire  [4:0] v$A1_6076_out0;
wire  [4:0] v$A1_6078_out0;
wire  [4:0] v$A1_6080_out0;
wire  [4:0] v$A1_6082_out0;
wire  [4:0] v$A1_8047_out0;
wire  [4:0] v$A1_8048_out0;
wire  [4:0] v$A2_10470_out0;
wire  [4:0] v$A2_10472_out0;
wire  [4:0] v$AMOUNT$OF$SHIFT_9833_out0;
wire  [4:0] v$AMOUNT$OF$SHIFT_9834_out0;
wire  [4:0] v$AMOUNT$OF$SHIFT_9835_out0;
wire  [4:0] v$AMOUNT$OF$SHIFT_9836_out0;
wire  [4:0] v$A_11864_out0;
wire  [4:0] v$A_11868_out0;
wire  [4:0] v$A_11880_out0;
wire  [4:0] v$A_11884_out0;
wire  [4:0] v$B$EXP_17294_out0;
wire  [4:0] v$B$EXP_17296_out0;
wire  [4:0] v$B$EXP_17298_out0;
wire  [4:0] v$B$EXP_17300_out0;
wire  [4:0] v$B_15036_out0;
wire  [4:0] v$B_15040_out0;
wire  [4:0] v$B_15052_out0;
wire  [4:0] v$B_15056_out0;
wire  [4:0] v$C1_14148_out0;
wire  [4:0] v$C1_14150_out0;
wire  [4:0] v$C1_14152_out0;
wire  [4:0] v$C1_14154_out0;
wire  [4:0] v$C1_16272_out0;
wire  [4:0] v$C1_16273_out0;
wire  [4:0] v$C1_16332_out0;
wire  [4:0] v$C1_16333_out0;
wire  [4:0] v$C1_5455_out0;
wire  [4:0] v$C1_5456_out0;
wire  [4:0] v$C1_6236_out0;
wire  [4:0] v$C1_6238_out0;
wire  [4:0] v$C1_7742_out0;
wire  [4:0] v$C1_7743_out0;
wire  [4:0] v$C3_7297_out0;
wire  [4:0] v$C3_7298_out0;
wire  [4:0] v$C4_15259_out0;
wire  [4:0] v$C4_15260_out0;
wire  [4:0] v$DIFF_9414_out0;
wire  [4:0] v$DIFF_9416_out0;
wire  [4:0] v$DIFF_9418_out0;
wire  [4:0] v$DIFF_9420_out0;
wire  [4:0] v$D_6009_out0;
wire  [4:0] v$D_6010_out0;
wire  [4:0] v$EXPONENT_16622_out0;
wire  [4:0] v$EXPONENT_16623_out0;
wire  [4:0] v$EXPONENT_17014_out0;
wire  [4:0] v$EXPONENT_17015_out0;
wire  [4:0] v$EXPONENT_18683_out0;
wire  [4:0] v$EXPONENT_18684_out0;
wire  [4:0] v$HALF$PRECISION$EXPONENT$DENORM_6394_out0;
wire  [4:0] v$HALF$PRECISION$EXPONENT$DENORM_6395_out0;
wire  [4:0] v$HALF$PRECISION$EXPONENT_15275_out0;
wire  [4:0] v$HALF$PRECISION$EXPONENT_15276_out0;
wire  [4:0] v$HALF$PRECISION$EXPONENT_6622_out0;
wire  [4:0] v$HALF$PRECISION$EXPONENT_6623_out0;
wire  [4:0] v$HALF$PRECISSION$ADDITION$IN_1291_out0;
wire  [4:0] v$HALF$PRECISSION$ADDITION$IN_1292_out0;
wire  [4:0] v$K_313_out0;
wire  [4:0] v$K_314_out0;
wire  [4:0] v$LARGER$EXP_10729_out0;
wire  [4:0] v$LARGER$EXP_10731_out0;
wire  [4:0] v$MUX1_15871_out0;
wire  [4:0] v$MUX1_15872_out0;
wire  [4:0] v$MUX1_18537_out0;
wire  [4:0] v$MUX1_18539_out0;
wire  [4:0] v$MUX1_18541_out0;
wire  [4:0] v$MUX1_18543_out0;
wire  [4:0] v$MUX1_19207_out0;
wire  [4:0] v$MUX1_19208_out0;
wire  [4:0] v$MUX1_5354_out0;
wire  [4:0] v$MUX1_5355_out0;
wire  [4:0] v$MUX2_14121_out0;
wire  [4:0] v$MUX2_14122_out0;
wire  [4:0] v$MUX3_3599_out0;
wire  [4:0] v$MUX3_3601_out0;
wire  [4:0] v$MUX3_3603_out0;
wire  [4:0] v$MUX3_3605_out0;
wire  [4:0] v$MUX5_4212_out0;
wire  [4:0] v$MUX5_4214_out0;
wire  [4:0] v$MUX5_4216_out0;
wire  [4:0] v$MUX5_4218_out0;
wire  [4:0] v$NORMALIZATION$SHIFT_1985_out0;
wire  [4:0] v$NORMALIZATION$SHIFT_1986_out0;
wire  [4:0] v$NORMALIZATION$SHIFT_4562_out0;
wire  [4:0] v$NORMALIZATION$SHIFT_4563_out0;
wire  [4:0] v$N_16856_out0;
wire  [4:0] v$N_16857_out0;
wire  [4:0] v$N_16858_out0;
wire  [4:0] v$N_16859_out0;
wire  [4:0] v$OUT_170_out0;
wire  [4:0] v$OUT_171_out0;
wire  [4:0] v$OUT_5217_out0;
wire  [4:0] v$OUT_5218_out0;
wire  [4:0] v$OUT_6454_out0;
wire  [4:0] v$OUT_6455_out0;
wire  [4:0] v$OUT_9253_out0;
wire  [4:0] v$OUT_9254_out0;
wire  [4:0] v$OUT_9281_out0;
wire  [4:0] v$OUT_9283_out0;
wire  [4:0] v$OUT_9285_out0;
wire  [4:0] v$OUT_9287_out0;
wire  [4:0] v$SEL10_3221_out0;
wire  [4:0] v$SEL10_3222_out0;
wire  [4:0] v$SEL14_9427_out0;
wire  [4:0] v$SEL14_9428_out0;
wire  [4:0] v$SEL18_18852_out0;
wire  [4:0] v$SEL18_18853_out0;
wire  [4:0] v$SEL1_7850_out0;
wire  [4:0] v$SEL1_7852_out0;
wire  [4:0] v$SEL1_7854_out0;
wire  [4:0] v$SEL1_7856_out0;
wire  [4:0] v$SEL1_9839_out0;
wire  [4:0] v$SEL1_9840_out0;
wire  [4:0] v$SEL25_14039_out0;
wire  [4:0] v$SEL25_14040_out0;
wire  [4:0] v$SEL25_14041_out0;
wire  [4:0] v$SEL25_14042_out0;
wire  [4:0] v$SEL2_7250_out0;
wire  [4:0] v$SEL2_7252_out0;
wire  [4:0] v$SEL2_7254_out0;
wire  [4:0] v$SEL2_7256_out0;
wire  [4:0] v$SEL9_3955_out0;
wire  [4:0] v$SEL9_3956_out0;
wire  [4:0] v$SMALLER$EXP_3150_out0;
wire  [4:0] v$SMALLER$EXP_3152_out0;
wire  [4:0] v$XOR1_11435_out0;
wire  [4:0] v$XOR1_11436_out0;
wire  [4:0] v$XOR1_4124_out0;
wire  [4:0] v$XOR1_4125_out0;
wire  [4:0] v$XOR1_7916_out0;
wire  [4:0] v$XOR1_7918_out0;
wire  [4:0] v$XOR1_7920_out0;
wire  [4:0] v$XOR1_7922_out0;
wire  [4:0] v$_1487_out0;
wire  [4:0] v$_1488_out0;
wire  [4:0] v$_2872_out0;
wire  [4:0] v$_2873_out0;
wire  [4:0] v$_3551_out0;
wire  [4:0] v$_3552_out0;
wire  [4:0] v$_5309_out0;
wire  [4:0] v$_5311_out0;
wire  [4:0] v$_5313_out0;
wire  [4:0] v$_5315_out0;
wire  [4:0] v$_6592_out0;
wire  [4:0] v$_6593_out0;
wire  [4:0] v$_7591_out0;
wire  [4:0] v$_7592_out0;
wire  [4:0] v$_9129_out0;
wire  [4:0] v$_9131_out0;
wire  [4:0] v$_9133_out0;
wire  [4:0] v$_9135_out0;
wire  [5:0] v$A1_4168_out0;
wire  [5:0] v$A1_4169_out0;
wire  [5:0] v$A2_15432_out0;
wire  [5:0] v$A2_15433_out0;
wire  [5:0] v$ADDRESS_15181_out0;
wire  [5:0] v$ADDRESS_15182_out0;
wire  [5:0] v$C2_16596_out0;
wire  [5:0] v$C2_16597_out0;
wire  [5:0] v$C3_13741_out0;
wire  [5:0] v$C3_13742_out0;
wire  [5:0] v$C6_8360_out0;
wire  [5:0] v$C6_8361_out0;
wire  [5:0] v$MUX1_10337_out0;
wire  [5:0] v$MUX1_10338_out0;
wire  [5:0] v$_1369_out0;
wire  [5:0] v$_1369_out1;
wire  [5:0] v$_1370_out0;
wire  [5:0] v$_1370_out1;
wire  [5:0] v$_1371_out0;
wire  [5:0] v$_1371_out1;
wire  [5:0] v$_1372_out0;
wire  [5:0] v$_1372_out1;
wire  [5:0] v$_1373_out0;
wire  [5:0] v$_1373_out1;
wire  [5:0] v$_1374_out0;
wire  [5:0] v$_1374_out1;
wire  [5:0] v$_16723_out0;
wire  [5:0] v$_16723_out1;
wire  [5:0] v$_16724_out0;
wire  [5:0] v$_16724_out1;
wire  [5:0] v$_16725_out0;
wire  [5:0] v$_16725_out1;
wire  [5:0] v$_16726_out0;
wire  [5:0] v$_16726_out1;
wire  [5:0] v$_16727_out0;
wire  [5:0] v$_16727_out1;
wire  [5:0] v$_16728_out0;
wire  [5:0] v$_16728_out1;
wire  [5:0] v$_1677_out0;
wire  [5:0] v$_1677_out1;
wire  [5:0] v$_1678_out0;
wire  [5:0] v$_1678_out1;
wire  [5:0] v$_1679_out0;
wire  [5:0] v$_1679_out1;
wire  [5:0] v$_1680_out0;
wire  [5:0] v$_1680_out1;
wire  [5:0] v$_1681_out0;
wire  [5:0] v$_1681_out1;
wire  [5:0] v$_1682_out0;
wire  [5:0] v$_1682_out1;
wire  [5:0] v$_17622_out0;
wire  [5:0] v$_17622_out1;
wire  [5:0] v$_17623_out0;
wire  [5:0] v$_17623_out1;
wire  [5:0] v$_17624_out0;
wire  [5:0] v$_17624_out1;
wire  [5:0] v$_17625_out0;
wire  [5:0] v$_17625_out1;
wire  [5:0] v$_17626_out0;
wire  [5:0] v$_17626_out1;
wire  [5:0] v$_17627_out0;
wire  [5:0] v$_17627_out1;
wire  [7:0] v$8LSB_7934_out0;
wire  [7:0] v$8LSB_7935_out0;
wire  [7:0] v$A$EXP_297_out0;
wire  [7:0] v$A$EXP_299_out0;
wire  [7:0] v$A$EXP_301_out0;
wire  [7:0] v$A$EXP_303_out0;
wire  [7:0] v$A1_16363_out0;
wire  [7:0] v$A1_16364_out0;
wire  [7:0] v$A1_2860_out0;
wire  [7:0] v$A1_2862_out0;
wire  [7:0] v$A1_6077_out0;
wire  [7:0] v$A1_6079_out0;
wire  [7:0] v$A1_6081_out0;
wire  [7:0] v$A1_6083_out0;
wire  [7:0] v$A1_698_out0;
wire  [7:0] v$A1_699_out0;
wire  [7:0] v$A2_10471_out0;
wire  [7:0] v$A2_10473_out0;
wire  [7:0] v$A_11857_out0;
wire  [7:0] v$A_11861_out0;
wire  [7:0] v$A_11865_out0;
wire  [7:0] v$A_11869_out0;
wire  [7:0] v$A_11873_out0;
wire  [7:0] v$A_11877_out0;
wire  [7:0] v$A_11881_out0;
wire  [7:0] v$A_11885_out0;
wire  [7:0] v$B$EXP_17295_out0;
wire  [7:0] v$B$EXP_17297_out0;
wire  [7:0] v$B$EXP_17299_out0;
wire  [7:0] v$B$EXP_17301_out0;
wire  [7:0] v$B_15029_out0;
wire  [7:0] v$B_15033_out0;
wire  [7:0] v$B_15037_out0;
wire  [7:0] v$B_15041_out0;
wire  [7:0] v$B_15045_out0;
wire  [7:0] v$B_15049_out0;
wire  [7:0] v$B_15053_out0;
wire  [7:0] v$B_15057_out0;
wire  [7:0] v$C1_14033_out0;
wire  [7:0] v$C1_14034_out0;
wire  [7:0] v$C1_14149_out0;
wire  [7:0] v$C1_14151_out0;
wire  [7:0] v$C1_14153_out0;
wire  [7:0] v$C1_14155_out0;
wire  [7:0] v$C1_14599_out0;
wire  [7:0] v$C1_14600_out0;
wire  [7:0] v$C1_15419_out0;
wire  [7:0] v$C1_15420_out0;
wire  [7:0] v$C1_1711_out0;
wire  [7:0] v$C1_1712_out0;
wire  [7:0] v$C1_6237_out0;
wire  [7:0] v$C1_6239_out0;
wire  [7:0] v$C1_6243_out0;
wire  [7:0] v$C1_6248_out0;
wire  [7:0] v$C1_6253_out0;
wire  [7:0] v$C1_6258_out0;
wire  [7:0] v$C1_6263_out0;
wire  [7:0] v$C1_6268_out0;
wire  [7:0] v$C1_6274_out0;
wire  [7:0] v$C1_6279_out0;
wire  [7:0] v$C1_6284_out0;
wire  [7:0] v$C1_6289_out0;
wire  [7:0] v$C1_6294_out0;
wire  [7:0] v$C1_6299_out0;
wire  [7:0] v$C1_8290_out0;
wire  [7:0] v$C1_8294_out0;
wire  [7:0] v$C2_105_out0;
wire  [7:0] v$C2_110_out0;
wire  [7:0] v$C2_115_out0;
wire  [7:0] v$C2_120_out0;
wire  [7:0] v$C2_125_out0;
wire  [7:0] v$C2_130_out0;
wire  [7:0] v$C2_136_out0;
wire  [7:0] v$C2_141_out0;
wire  [7:0] v$C2_146_out0;
wire  [7:0] v$C2_151_out0;
wire  [7:0] v$C2_156_out0;
wire  [7:0] v$C2_161_out0;
wire  [7:0] v$DIFF$VIEW$MANTISA$ADDER_13293_out0;
wire  [7:0] v$DIFF$VIEW$MANTISA$ADDER_13294_out0;
wire  [7:0] v$DIFF_13242_out0;
wire  [7:0] v$DIFF_13243_out0;
wire  [7:0] v$DIFF_16536_out0;
wire  [7:0] v$DIFF_16537_out0;
wire  [7:0] v$DIFF_18144_out0;
wire  [7:0] v$DIFF_18145_out0;
wire  [7:0] v$DIFF_18146_out0;
wire  [7:0] v$DIFF_18147_out0;
wire  [7:0] v$DIFF_3044_out0;
wire  [7:0] v$DIFF_3045_out0;
wire  [7:0] v$DIFF_304_out0;
wire  [7:0] v$DIFF_305_out0;
wire  [7:0] v$DIFF_9415_out0;
wire  [7:0] v$DIFF_9417_out0;
wire  [7:0] v$DIFF_9419_out0;
wire  [7:0] v$DIFF_9421_out0;
wire  [7:0] v$EDGEMODE_3092_out0;
wire  [7:0] v$EDGEMODE_3093_out0;
wire  [7:0] v$END_13282_out0;
wire  [7:0] v$END_13283_out0;
wire  [7:0] v$EXP$DIFF_13064_out0;
wire  [7:0] v$EXP$DIFF_13065_out0;
wire  [7:0] v$EXP$DIFF_14375_out0;
wire  [7:0] v$EXP$DIFF_14376_out0;
wire  [7:0] v$EXP$DIFF_14934_out0;
wire  [7:0] v$EXP$DIFF_14935_out0;
wire  [7:0] v$EXP$DIFF_18281_out0;
wire  [7:0] v$EXP$DIFF_18282_out0;
wire  [7:0] v$EXPONENT_14267_out0;
wire  [7:0] v$EXPONENT_14268_out0;
wire  [7:0] v$EXPONENT_1521_out0;
wire  [7:0] v$EXPONENT_1522_out0;
wire  [7:0] v$IN_15465_out0;
wire  [7:0] v$IN_15466_out0;
wire  [7:0] v$IN_15467_out0;
wire  [7:0] v$IN_15468_out0;
wire  [7:0] v$IN_15469_out0;
wire  [7:0] v$IN_15470_out0;
wire  [7:0] v$IN_15471_out0;
wire  [7:0] v$IN_15472_out0;
wire  [7:0] v$IN_15473_out0;
wire  [7:0] v$IN_15474_out0;
wire  [7:0] v$LARGER$EXP_10730_out0;
wire  [7:0] v$LARGER$EXP_10732_out0;
wire  [7:0] v$LSBS_8263_out0;
wire  [7:0] v$LSBS_8264_out0;
wire  [7:0] v$MODEIN_6068_out0;
wire  [7:0] v$MODEIN_6069_out0;
wire  [7:0] v$MODE_11296_out0;
wire  [7:0] v$MODE_11297_out0;
wire  [7:0] v$MODE_18452_out0;
wire  [7:0] v$MODE_18453_out0;
wire  [7:0] v$MODE_50_out0;
wire  [7:0] v$MODE_51_out0;
wire  [7:0] v$MUX13_10825_out0;
wire  [7:0] v$MUX13_10826_out0;
wire  [7:0] v$MUX1_18538_out0;
wire  [7:0] v$MUX1_18540_out0;
wire  [7:0] v$MUX1_18542_out0;
wire  [7:0] v$MUX1_18544_out0;
wire  [7:0] v$MUX2_18372_out0;
wire  [7:0] v$MUX2_18373_out0;
wire  [7:0] v$MUX3_3600_out0;
wire  [7:0] v$MUX3_3602_out0;
wire  [7:0] v$MUX3_3604_out0;
wire  [7:0] v$MUX3_3606_out0;
wire  [7:0] v$MUX5_13753_out0;
wire  [7:0] v$MUX5_13754_out0;
wire  [7:0] v$MUX6_14288_out0;
wire  [7:0] v$MUX6_14289_out0;
wire  [7:0] v$MUX6_8275_out0;
wire  [7:0] v$MUX6_8276_out0;
wire  [7:0] v$NORMALIZATION$SHIFT$WHOLE_6909_out0;
wire  [7:0] v$NORMALIZATION$SHIFT$WHOLE_6910_out0;
wire  [7:0] v$NORMALIZATION$SHIFT_11230_out0;
wire  [7:0] v$NORMALIZATION$SHIFT_11231_out0;
wire  [7:0] v$NORMALIZATION$SHIFT_1311_out0;
wire  [7:0] v$NORMALIZATION$SHIFT_1312_out0;
wire  [7:0] v$NORMALIZATION$SHIFT_19233_out0;
wire  [7:0] v$NORMALIZATION$SHIFT_19234_out0;
wire  [7:0] v$NORMALIZATION$SHIFT_3477_out0;
wire  [7:0] v$NORMALIZATION$SHIFT_3478_out0;
wire  [7:0] v$N_14681_out0;
wire  [7:0] v$N_14682_out0;
wire  [7:0] v$N_14683_out0;
wire  [7:0] v$N_14684_out0;
wire  [7:0] v$OUT_15386_out0;
wire  [7:0] v$OUT_15387_out0;
wire  [7:0] v$OUT_16707_out0;
wire  [7:0] v$OUT_16708_out0;
wire  [7:0] v$PIN_6869_out0;
wire  [7:0] v$PIN_6870_out0;
wire  [7:0] v$PIN_6871_out0;
wire  [7:0] v$PIN_6872_out0;
wire  [7:0] v$PIN_6873_out0;
wire  [7:0] v$PIN_6874_out0;
wire  [7:0] v$PIN_6875_out0;
wire  [7:0] v$PIN_6876_out0;
wire  [7:0] v$PIN_6877_out0;
wire  [7:0] v$PIN_6878_out0;
wire  [7:0] v$PIN_6879_out0;
wire  [7:0] v$PIN_6880_out0;
wire  [7:0] v$POUT_10823_out0;
wire  [7:0] v$POUT_10824_out0;
wire  [7:0] v$POut_14269_out0;
wire  [7:0] v$POut_14270_out0;
wire  [7:0] v$RXBYTE_10010_out0;
wire  [7:0] v$RXBYTE_10011_out0;
wire  [7:0] v$RXBYTE_18996_out0;
wire  [7:0] v$RXBYTE_18997_out0;
wire  [7:0] v$SEL17_5630_out0;
wire  [7:0] v$SEL17_5631_out0;
wire  [7:0] v$SEL1_15974_out0;
wire  [7:0] v$SEL1_15979_out0;
wire  [7:0] v$SEL1_15984_out0;
wire  [7:0] v$SEL1_15992_out0;
wire  [7:0] v$SEL1_15994_out0;
wire  [7:0] v$SEL1_16002_out0;
wire  [7:0] v$SEL1_16005_out0;
wire  [7:0] v$SEL1_16010_out0;
wire  [7:0] v$SEL1_16015_out0;
wire  [7:0] v$SEL1_16023_out0;
wire  [7:0] v$SEL1_16025_out0;
wire  [7:0] v$SEL1_16033_out0;
wire  [7:0] v$SEL1_17306_out0;
wire  [7:0] v$SEL1_17308_out0;
wire  [7:0] v$SEL1_17310_out0;
wire  [7:0] v$SEL1_17312_out0;
wire  [7:0] v$SEL1_18066_out0;
wire  [7:0] v$SEL1_18067_out0;
wire  [7:0] v$SEL1_368_out0;
wire  [7:0] v$SEL1_369_out0;
wire  [7:0] v$SEL1_7851_out0;
wire  [7:0] v$SEL1_7853_out0;
wire  [7:0] v$SEL1_7855_out0;
wire  [7:0] v$SEL1_7857_out0;
wire  [7:0] v$SEL1_8397_out0;
wire  [7:0] v$SEL1_8398_out0;
wire  [7:0] v$SEL1_8399_out0;
wire  [7:0] v$SEL1_8400_out0;
wire  [7:0] v$SEL1_9046_out0;
wire  [7:0] v$SEL1_9051_out0;
wire  [7:0] v$SEL1_9056_out0;
wire  [7:0] v$SEL1_9064_out0;
wire  [7:0] v$SEL1_9066_out0;
wire  [7:0] v$SEL1_9074_out0;
wire  [7:0] v$SEL1_9077_out0;
wire  [7:0] v$SEL1_9082_out0;
wire  [7:0] v$SEL1_9087_out0;
wire  [7:0] v$SEL1_9095_out0;
wire  [7:0] v$SEL1_9097_out0;
wire  [7:0] v$SEL1_9105_out0;
wire  [7:0] v$SEL2_18013_out0;
wire  [7:0] v$SEL2_18014_out0;
wire  [7:0] v$SEL2_18152_out0;
wire  [7:0] v$SEL2_18153_out0;
wire  [7:0] v$SEL2_18154_out0;
wire  [7:0] v$SEL2_18155_out0;
wire  [7:0] v$SEL2_7251_out0;
wire  [7:0] v$SEL2_7253_out0;
wire  [7:0] v$SEL2_7255_out0;
wire  [7:0] v$SEL2_7257_out0;
wire  [7:0] v$SEL3_18385_out0;
wire  [7:0] v$SEL3_18386_out0;
wire  [7:0] v$SEL3_18423_out0;
wire  [7:0] v$SEL3_18424_out0;
wire  [7:0] v$SEL4_12427_out0;
wire  [7:0] v$SEL4_12428_out0;
wire  [7:0] v$SEL4_12764_out0;
wire  [7:0] v$SEL4_12765_out0;
wire  [7:0] v$SHIFT$AMOUNT_7702_out0;
wire  [7:0] v$SHIFT$AMOUNT_7703_out0;
wire  [7:0] v$SHIFT$AMOUNT_7704_out0;
wire  [7:0] v$SHIFT$AMOUNT_7705_out0;
wire  [7:0] v$SHIFT$AMOUNT_7706_out0;
wire  [7:0] v$SHIFT$AMOUNT_7707_out0;
wire  [7:0] v$SHIFT$AMOUNT_7708_out0;
wire  [7:0] v$SHIFT$AMOUNT_7709_out0;
wire  [7:0] v$SINGLE$EXPONENT_7376_out0;
wire  [7:0] v$SINGLE$EXPONENT_7377_out0;
wire  [7:0] v$SINGLE$PRECISION$EXPONENT_11558_out0;
wire  [7:0] v$SINGLE$PRECISION$EXPONENT_11559_out0;
wire  [7:0] v$SMALLER$EXP_3151_out0;
wire  [7:0] v$SMALLER$EXP_3153_out0;
wire  [7:0] v$STATUS_32_out0;
wire  [7:0] v$STATUS_33_out0;
wire  [7:0] v$STATUS_9155_out0;
wire  [7:0] v$STATUS_9156_out0;
wire  [7:0] v$Status_3973_out0;
wire  [7:0] v$Status_3974_out0;
wire  [7:0] v$XOR1_15146_out0;
wire  [7:0] v$XOR1_15147_out0;
wire  [7:0] v$XOR1_7917_out0;
wire  [7:0] v$XOR1_7919_out0;
wire  [7:0] v$XOR1_7921_out0;
wire  [7:0] v$XOR1_7923_out0;
wire  [7:0] v$_10833_out0;
wire  [7:0] v$_10834_out0;
wire  [7:0] v$_1319_out0;
wire  [7:0] v$_1320_out0;
wire  [7:0] v$_1321_out0;
wire  [7:0] v$_1322_out0;
wire  [7:0] v$_1323_out0;
wire  [7:0] v$_1324_out0;
wire  [7:0] v$_13473_out1;
wire  [7:0] v$_13474_out1;
wire  [7:0] v$_13855_out0;
wire  [7:0] v$_13858_out0;
wire  [7:0] v$_14705_out0;
wire  [7:0] v$_14706_out0;
wire  [7:0] v$_14916_out0;
wire  [7:0] v$_14917_out0;
wire  [7:0] v$_15204_out0;
wire  [7:0] v$_15208_out0;
wire  [7:0] v$_15240_out0;
wire  [7:0] v$_15244_out0;
wire  [7:0] v$_15255_out0;
wire  [7:0] v$_15256_out0;
wire  [7:0] v$_16264_out0;
wire  [7:0] v$_16265_out0;
wire  [7:0] v$_16778_out0;
wire  [7:0] v$_16779_out0;
wire  [7:0] v$_1683_out0;
wire  [7:0] v$_1683_out1;
wire  [7:0] v$_1684_out0;
wire  [7:0] v$_1684_out1;
wire  [7:0] v$_17371_out0;
wire  [7:0] v$_17375_out0;
wire  [7:0] v$_17381_out0;
wire  [7:0] v$_17381_out1;
wire  [7:0] v$_17382_out0;
wire  [7:0] v$_17382_out1;
wire  [7:0] v$_17995_out0;
wire  [7:0] v$_17996_out0;
wire  [7:0] v$_17997_out0;
wire  [7:0] v$_17998_out0;
wire  [7:0] v$_17999_out0;
wire  [7:0] v$_18000_out0;
wire  [7:0] v$_18048_out0;
wire  [7:0] v$_18049_out0;
wire  [7:0] v$_1827_out0;
wire  [7:0] v$_1828_out0;
wire  [7:0] v$_1829_out0;
wire  [7:0] v$_1829_out1;
wire  [7:0] v$_1830_out0;
wire  [7:0] v$_1830_out1;
wire  [7:0] v$_18358_out0;
wire  [7:0] v$_18359_out0;
wire  [7:0] v$_18360_out0;
wire  [7:0] v$_18361_out0;
wire  [7:0] v$_18362_out0;
wire  [7:0] v$_18363_out0;
wire  [7:0] v$_3866_out0;
wire  [7:0] v$_3867_out0;
wire  [7:0] v$_4248_out0;
wire  [7:0] v$_4249_out0;
wire  [7:0] v$_4250_out0;
wire  [7:0] v$_4251_out0;
wire  [7:0] v$_4252_out0;
wire  [7:0] v$_4253_out0;
wire  [7:0] v$_5016_out0;
wire  [7:0] v$_5020_out0;
wire  [7:0] v$_6893_out0;
wire  [7:0] v$_6894_out0;
wire  [7:0] v$_6895_out0;
wire  [7:0] v$_6896_out0;
wire  [7:0] v$_6897_out0;
wire  [7:0] v$_6898_out0;
wire  [7:0] v$_7595_out1;
wire  [7:0] v$_7938_out0;
wire  [7:0] v$_7939_out0;
wire  [7:0] v$_8112_out0;
wire  [7:0] v$_8113_out0;
wire  [7:0] v$_8114_out0;
wire  [7:0] v$_8115_out0;
wire  [7:0] v$_8116_out0;
wire  [7:0] v$_8117_out0;
wire  [7:0] v$_8229_out0;
wire  [7:0] v$_8229_out1;
wire  [7:0] v$_8230_out0;
wire  [7:0] v$_8230_out1;
wire  [7:0] v$_9303_out0;
wire  [7:0] v$_9303_out1;
wire  [7:0] v$_9304_out0;
wire  [7:0] v$_9304_out1;
wire  [7:0] v$_9369_out0;
wire  [7:0] v$_9370_out0;
wire  [9:0] v$HALF$PRECISION$MANTISA$DENORM_15096_out0;
wire  [9:0] v$HALF$PRECISION$MANTISA$DENORM_15097_out0;
wire  [9:0] v$SEL10_3429_out0;
wire  [9:0] v$SEL10_3430_out0;
wire  [9:0] v$SEL12_16_out0;
wire  [9:0] v$SEL12_17_out0;
wire  [9:0] v$SEL2_8412_out0;
wire  [9:0] v$SEL2_8413_out0;
wire  [9:0] v$SEL5_8136_out0;
wire  [9:0] v$SEL5_8137_out0;
wire  [9:0] v$SEL7_13070_out0;
wire  [9:0] v$SEL7_13071_out0;
wire  [9:0] v$SEL7_3499_out0;
wire  [9:0] v$SEL7_3500_out0;
wire  [9:0] v$SEL9_10394_out0;
wire  [9:0] v$SEL9_10395_out0;
wire  [9:0] v$_2613_out0;
wire  [9:0] v$_2810_out0;
wire v$1_1687_out0;
wire v$1_1688_out0;
wire v$2StopBits_3683_out0;
wire v$2StopBits_3684_out0;
wire v$32$BIT$INPUT_206_out0;
wire v$32$BIT$INPUT_207_out0;
wire v$32$BIT$VIEWER$IN$FPU_4548_out0;
wire v$32$BIT$VIEWER$IN$FPU_4549_out0;
wire v$32BIT_11437_out0;
wire v$32BIT_11438_out0;
wire v$32BIT_16476_out0;
wire v$32BIT_16477_out0;
wire v$4_15776_out0;
wire v$4_15777_out0;
wire v$5_12857_out0;
wire v$5_12858_out0;
wire v$6_10287_out0;
wire v$6_10288_out0;
wire v$6_2112_out0;
wire v$6_2113_out0;
wire v$7_15947_out0;
wire v$7_15948_out0;
wire v$8_16131_out0;
wire v$8_16132_out0;
wire v$A$EXP$LARGER_18122_out0;
wire v$A$EXP$LARGER_18123_out0;
wire v$A$EXP$LARGER_18846_out0;
wire v$A$EXP$LARGER_18847_out0;
wire v$A$EXP$LARGER_9815_out0;
wire v$A$EXP$LARGER_9816_out0;
wire v$A$IS$OP1_5221_out0;
wire v$A$IS$OP1_5222_out0;
wire v$A$MANTISA$LARGER_15319_out0;
wire v$A$MANTISA$LARGER_15320_out0;
wire v$A$MANTISA$LARGER_16641_out0;
wire v$A$MANTISA$LARGER_16642_out0;
wire v$A0$COMP$B0_8303_out0;
wire v$A0$COMP$B0_8304_out0;
wire v$A0$COMP$B0_8305_out0;
wire v$A0$COMP$B0_8306_out0;
wire v$A0$COMP$B0_8307_out0;
wire v$A0$COMP$B0_8308_out0;
wire v$A0$COMP$B0_8309_out0;
wire v$A0$COMP$B0_8310_out0;
wire v$A0$COMP$B0_8311_out0;
wire v$A0$COMP$B0_8312_out0;
wire v$A0$COMP$B0_8313_out0;
wire v$A0$COMP$B0_8314_out0;
wire v$A0$COMP$B0_8315_out0;
wire v$A0$COMP$B0_8316_out0;
wire v$A0$COMP$B0_8317_out0;
wire v$A0$COMP$B0_8318_out0;
wire v$A0$COMP$B0_8319_out0;
wire v$A0$COMP$B0_8320_out0;
wire v$A0$COMP$B0_8321_out0;
wire v$A0$COMP$B0_8322_out0;
wire v$A0$COMP$B0_8323_out0;
wire v$A0$COMP$B0_8324_out0;
wire v$A0$COMP$B0_8325_out0;
wire v$A0$COMP$B0_8326_out0;
wire v$A0XNORB0_1583_out0;
wire v$A0XNORB0_1584_out0;
wire v$A0XNORB0_1585_out0;
wire v$A0XNORB0_1586_out0;
wire v$A0XNORB0_1587_out0;
wire v$A0XNORB0_1588_out0;
wire v$A0XNORB0_1589_out0;
wire v$A0XNORB0_1590_out0;
wire v$A0XNORB0_1591_out0;
wire v$A0XNORB0_1592_out0;
wire v$A0XNORB0_1593_out0;
wire v$A0XNORB0_1594_out0;
wire v$A0XNORB0_1595_out0;
wire v$A0XNORB0_1596_out0;
wire v$A0XNORB0_1597_out0;
wire v$A0XNORB0_1598_out0;
wire v$A0XNORB0_1599_out0;
wire v$A0XNORB0_1600_out0;
wire v$A0XNORB0_1601_out0;
wire v$A0XNORB0_1602_out0;
wire v$A0XNORB0_1603_out0;
wire v$A0XNORB0_1604_out0;
wire v$A0XNORB0_1605_out0;
wire v$A0XNORB0_1606_out0;
wire v$A0_1885_out0;
wire v$A0_1886_out0;
wire v$A0_1887_out0;
wire v$A0_1888_out0;
wire v$A0_1889_out0;
wire v$A0_1890_out0;
wire v$A0_1891_out0;
wire v$A0_1892_out0;
wire v$A0_1893_out0;
wire v$A0_1894_out0;
wire v$A0_1895_out0;
wire v$A0_1896_out0;
wire v$A0_1897_out0;
wire v$A0_1898_out0;
wire v$A0_1899_out0;
wire v$A0_1900_out0;
wire v$A0_1901_out0;
wire v$A0_1902_out0;
wire v$A0_1903_out0;
wire v$A0_1904_out0;
wire v$A0_1905_out0;
wire v$A0_1906_out0;
wire v$A0_1907_out0;
wire v$A0_1908_out0;
wire v$A0_4468_out0;
wire v$A0_4469_out0;
wire v$A0_4470_out0;
wire v$A0_4471_out0;
wire v$A0_4472_out0;
wire v$A0_4473_out0;
wire v$A1$COMP$B1_13080_out0;
wire v$A1$COMP$B1_13081_out0;
wire v$A1$COMP$B1_13082_out0;
wire v$A1$COMP$B1_13083_out0;
wire v$A1$COMP$B1_13084_out0;
wire v$A1$COMP$B1_13085_out0;
wire v$A1$COMP$B1_13086_out0;
wire v$A1$COMP$B1_13087_out0;
wire v$A1$COMP$B1_13088_out0;
wire v$A1$COMP$B1_13089_out0;
wire v$A1$COMP$B1_13090_out0;
wire v$A1$COMP$B1_13091_out0;
wire v$A1$COMP$B1_13092_out0;
wire v$A1$COMP$B1_13093_out0;
wire v$A1$COMP$B1_13094_out0;
wire v$A1$COMP$B1_13095_out0;
wire v$A1$COMP$B1_13096_out0;
wire v$A1$COMP$B1_13097_out0;
wire v$A1$COMP$B1_13098_out0;
wire v$A1$COMP$B1_13099_out0;
wire v$A1$COMP$B1_13100_out0;
wire v$A1$COMP$B1_13101_out0;
wire v$A1$COMP$B1_13102_out0;
wire v$A1$COMP$B1_13103_out0;
wire v$A10A_16612_out0;
wire v$A10A_16612_out1;
wire v$A10A_16613_out0;
wire v$A10A_16613_out1;
wire v$A10A_16614_out0;
wire v$A10A_16614_out1;
wire v$A10A_16615_out0;
wire v$A10A_16615_out1;
wire v$A10A_16616_out0;
wire v$A10A_16616_out1;
wire v$A10A_16617_out0;
wire v$A10A_16617_out1;
wire v$A10_1703_out0;
wire v$A10_1704_out0;
wire v$A10_1705_out0;
wire v$A10_1706_out0;
wire v$A10_1707_out0;
wire v$A10_1708_out0;
wire v$A11_10386_out0;
wire v$A11_10387_out0;
wire v$A11_10388_out0;
wire v$A11_10389_out0;
wire v$A11_10390_out0;
wire v$A11_10391_out0;
wire v$A11_18484_out0;
wire v$A11_18484_out1;
wire v$A11_18485_out0;
wire v$A11_18485_out1;
wire v$A11_18486_out0;
wire v$A11_18486_out1;
wire v$A11_18487_out0;
wire v$A11_18487_out1;
wire v$A11_18488_out0;
wire v$A11_18488_out1;
wire v$A11_18489_out0;
wire v$A11_18489_out1;
wire v$A12A_4613_out0;
wire v$A12A_4613_out1;
wire v$A12A_4614_out0;
wire v$A12A_4614_out1;
wire v$A12A_4615_out0;
wire v$A12A_4615_out1;
wire v$A12A_4616_out0;
wire v$A12A_4616_out1;
wire v$A12A_4617_out0;
wire v$A12A_4617_out1;
wire v$A12A_4618_out0;
wire v$A12A_4618_out1;
wire v$A12_3355_out0;
wire v$A12_3356_out0;
wire v$A12_3357_out0;
wire v$A12_3358_out0;
wire v$A12_3359_out0;
wire v$A12_3360_out0;
wire v$A13_14445_out0;
wire v$A13_14446_out0;
wire v$A13_14447_out0;
wire v$A13_14448_out0;
wire v$A13_14449_out0;
wire v$A13_14450_out0;
wire v$A13_7554_out0;
wire v$A13_7554_out1;
wire v$A13_7555_out0;
wire v$A13_7555_out1;
wire v$A13_7556_out0;
wire v$A13_7556_out1;
wire v$A13_7557_out0;
wire v$A13_7557_out1;
wire v$A13_7558_out0;
wire v$A13_7558_out1;
wire v$A13_7559_out0;
wire v$A13_7559_out1;
wire v$A14_15941_out0;
wire v$A14_15941_out1;
wire v$A14_15942_out0;
wire v$A14_15942_out1;
wire v$A14_15943_out0;
wire v$A14_15943_out1;
wire v$A14_15944_out0;
wire v$A14_15944_out1;
wire v$A14_15945_out0;
wire v$A14_15945_out1;
wire v$A14_15946_out0;
wire v$A14_15946_out1;
wire v$A14_738_out0;
wire v$A14_739_out0;
wire v$A14_740_out0;
wire v$A14_741_out0;
wire v$A14_742_out0;
wire v$A14_743_out0;
wire v$A15_13797_out0;
wire v$A15_13797_out1;
wire v$A15_13798_out0;
wire v$A15_13798_out1;
wire v$A15_13799_out0;
wire v$A15_13799_out1;
wire v$A15_13800_out0;
wire v$A15_13800_out1;
wire v$A15_13801_out0;
wire v$A15_13801_out1;
wire v$A15_13802_out0;
wire v$A15_13802_out1;
wire v$A15_17957_out0;
wire v$A15_17958_out0;
wire v$A15_17959_out0;
wire v$A15_17960_out0;
wire v$A15_17961_out0;
wire v$A15_17962_out0;
wire v$A16A_15158_out0;
wire v$A16A_15158_out1;
wire v$A16A_15159_out0;
wire v$A16A_15159_out1;
wire v$A16A_15160_out0;
wire v$A16A_15160_out1;
wire v$A16A_15161_out0;
wire v$A16A_15161_out1;
wire v$A16A_15162_out0;
wire v$A16A_15162_out1;
wire v$A16A_15163_out0;
wire v$A16A_15163_out1;
wire v$A16_14191_out0;
wire v$A16_14192_out0;
wire v$A16_14193_out0;
wire v$A16_14194_out0;
wire v$A16_14195_out0;
wire v$A16_14196_out0;
wire v$A17A_2682_out0;
wire v$A17A_2682_out1;
wire v$A17A_2683_out0;
wire v$A17A_2683_out1;
wire v$A17A_2684_out0;
wire v$A17A_2684_out1;
wire v$A17A_2685_out0;
wire v$A17A_2685_out1;
wire v$A17A_2686_out0;
wire v$A17A_2686_out1;
wire v$A17A_2687_out0;
wire v$A17A_2687_out1;
wire v$A17_17342_out0;
wire v$A17_17343_out0;
wire v$A17_17344_out0;
wire v$A17_17345_out0;
wire v$A17_17346_out0;
wire v$A17_17347_out0;
wire v$A18_10458_out0;
wire v$A18_10458_out1;
wire v$A18_10459_out0;
wire v$A18_10459_out1;
wire v$A18_10460_out0;
wire v$A18_10460_out1;
wire v$A18_10461_out0;
wire v$A18_10461_out1;
wire v$A18_10462_out0;
wire v$A18_10462_out1;
wire v$A18_10463_out0;
wire v$A18_10463_out1;
wire v$A18_18300_out0;
wire v$A18_18301_out0;
wire v$A18_18302_out0;
wire v$A18_18303_out0;
wire v$A18_18304_out0;
wire v$A18_18305_out0;
wire v$A19_1363_out0;
wire v$A19_1364_out0;
wire v$A19_1365_out0;
wire v$A19_1366_out0;
wire v$A19_1367_out0;
wire v$A19_1368_out0;
wire v$A19_16511_out0;
wire v$A19_16511_out1;
wire v$A19_16512_out0;
wire v$A19_16512_out1;
wire v$A19_16513_out0;
wire v$A19_16513_out1;
wire v$A19_16514_out0;
wire v$A19_16514_out1;
wire v$A19_16515_out0;
wire v$A19_16515_out1;
wire v$A19_16516_out0;
wire v$A19_16516_out1;
wire v$A1A_12224_out0;
wire v$A1A_12224_out1;
wire v$A1A_12225_out0;
wire v$A1A_12225_out1;
wire v$A1A_12226_out0;
wire v$A1A_12226_out1;
wire v$A1A_12227_out0;
wire v$A1A_12227_out1;
wire v$A1A_12228_out0;
wire v$A1A_12228_out1;
wire v$A1A_12229_out0;
wire v$A1A_12229_out1;
wire v$A1XNORB1_16659_out0;
wire v$A1XNORB1_16660_out0;
wire v$A1XNORB1_16661_out0;
wire v$A1XNORB1_16662_out0;
wire v$A1XNORB1_16663_out0;
wire v$A1XNORB1_16664_out0;
wire v$A1XNORB1_16665_out0;
wire v$A1XNORB1_16666_out0;
wire v$A1XNORB1_16667_out0;
wire v$A1XNORB1_16668_out0;
wire v$A1XNORB1_16669_out0;
wire v$A1XNORB1_16670_out0;
wire v$A1XNORB1_16671_out0;
wire v$A1XNORB1_16672_out0;
wire v$A1XNORB1_16673_out0;
wire v$A1XNORB1_16674_out0;
wire v$A1XNORB1_16675_out0;
wire v$A1XNORB1_16676_out0;
wire v$A1XNORB1_16677_out0;
wire v$A1XNORB1_16678_out0;
wire v$A1XNORB1_16679_out0;
wire v$A1XNORB1_16680_out0;
wire v$A1XNORB1_16681_out0;
wire v$A1XNORB1_16682_out0;
wire v$A1_12374_out1;
wire v$A1_12375_out1;
wire v$A1_14282_out1;
wire v$A1_14283_out1;
wire v$A1_14943_out0;
wire v$A1_14944_out0;
wire v$A1_14945_out0;
wire v$A1_14946_out0;
wire v$A1_14947_out0;
wire v$A1_14948_out0;
wire v$A1_14949_out0;
wire v$A1_14950_out0;
wire v$A1_14951_out0;
wire v$A1_14952_out0;
wire v$A1_14953_out0;
wire v$A1_14954_out0;
wire v$A1_14955_out0;
wire v$A1_14956_out0;
wire v$A1_14957_out0;
wire v$A1_14958_out0;
wire v$A1_14959_out0;
wire v$A1_14960_out0;
wire v$A1_14961_out0;
wire v$A1_14962_out0;
wire v$A1_14963_out0;
wire v$A1_14964_out0;
wire v$A1_14965_out0;
wire v$A1_14966_out0;
wire v$A1_15427_out1;
wire v$A1_15428_out1;
wire v$A1_16363_out1;
wire v$A1_16364_out1;
wire v$A1_1869_out0;
wire v$A1_1870_out0;
wire v$A1_1871_out0;
wire v$A1_1872_out0;
wire v$A1_1873_out0;
wire v$A1_1874_out0;
wire v$A1_2859_out1;
wire v$A1_2860_out1;
wire v$A1_2861_out1;
wire v$A1_2862_out1;
wire v$A1_3146_out1;
wire v$A1_3147_out1;
wire v$A1_4168_out1;
wire v$A1_4169_out1;
wire v$A1_6076_out1;
wire v$A1_6077_out1;
wire v$A1_6078_out1;
wire v$A1_6079_out1;
wire v$A1_6080_out1;
wire v$A1_6081_out1;
wire v$A1_6082_out1;
wire v$A1_6083_out1;
wire v$A1_6652_out1;
wire v$A1_6653_out1;
wire v$A1_698_out1;
wire v$A1_699_out1;
wire v$A1_8047_out1;
wire v$A1_8048_out1;
wire v$A1_9805_out1;
wire v$A1_9806_out1;
wire v$A2$COMP$B2_2135_out0;
wire v$A2$COMP$B2_2136_out0;
wire v$A2$COMP$B2_2137_out0;
wire v$A2$COMP$B2_2138_out0;
wire v$A2$COMP$B2_2139_out0;
wire v$A2$COMP$B2_2140_out0;
wire v$A2$COMP$B2_2141_out0;
wire v$A2$COMP$B2_2142_out0;
wire v$A2$COMP$B2_2143_out0;
wire v$A2$COMP$B2_2144_out0;
wire v$A2$COMP$B2_2145_out0;
wire v$A2$COMP$B2_2146_out0;
wire v$A2$COMP$B2_2147_out0;
wire v$A2$COMP$B2_2148_out0;
wire v$A2$COMP$B2_2149_out0;
wire v$A2$COMP$B2_2150_out0;
wire v$A2$COMP$B2_2151_out0;
wire v$A2$COMP$B2_2152_out0;
wire v$A2$COMP$B2_2153_out0;
wire v$A2$COMP$B2_2154_out0;
wire v$A2$COMP$B2_2155_out0;
wire v$A2$COMP$B2_2156_out0;
wire v$A2$COMP$B2_2157_out0;
wire v$A2$COMP$B2_2158_out0;
wire v$A20_16992_out0;
wire v$A20_16992_out1;
wire v$A20_16993_out0;
wire v$A20_16993_out1;
wire v$A20_16994_out0;
wire v$A20_16994_out1;
wire v$A20_16995_out0;
wire v$A20_16995_out1;
wire v$A20_16996_out0;
wire v$A20_16996_out1;
wire v$A20_16997_out0;
wire v$A20_16997_out1;
wire v$A20_4603_out0;
wire v$A20_4604_out0;
wire v$A20_4605_out0;
wire v$A20_4606_out0;
wire v$A20_4607_out0;
wire v$A20_4608_out0;
wire v$A21_19179_out0;
wire v$A21_19179_out1;
wire v$A21_19180_out0;
wire v$A21_19180_out1;
wire v$A21_19181_out0;
wire v$A21_19181_out1;
wire v$A21_19182_out0;
wire v$A21_19182_out1;
wire v$A21_19183_out0;
wire v$A21_19183_out1;
wire v$A21_19184_out0;
wire v$A21_19184_out1;
wire v$A21_2792_out0;
wire v$A21_2793_out0;
wire v$A21_2794_out0;
wire v$A21_2795_out0;
wire v$A21_2796_out0;
wire v$A21_2797_out0;
wire v$A22_18127_out0;
wire v$A22_18127_out1;
wire v$A22_18128_out0;
wire v$A22_18128_out1;
wire v$A22_18129_out0;
wire v$A22_18129_out1;
wire v$A22_18130_out0;
wire v$A22_18130_out1;
wire v$A22_18131_out0;
wire v$A22_18131_out1;
wire v$A22_18132_out0;
wire v$A22_18132_out1;
wire v$A22_4590_out0;
wire v$A22_4591_out0;
wire v$A22_4592_out0;
wire v$A22_4593_out0;
wire v$A22_4594_out0;
wire v$A22_4595_out0;
wire v$A23_5281_out0;
wire v$A23_5282_out0;
wire v$A23_5283_out0;
wire v$A23_5284_out0;
wire v$A23_5285_out0;
wire v$A23_5286_out0;
wire v$A23_9924_out0;
wire v$A23_9924_out1;
wire v$A23_9925_out0;
wire v$A23_9925_out1;
wire v$A23_9926_out0;
wire v$A23_9926_out1;
wire v$A23_9927_out0;
wire v$A23_9927_out1;
wire v$A23_9928_out0;
wire v$A23_9928_out1;
wire v$A23_9929_out0;
wire v$A23_9929_out1;
wire v$A24_17569_out0;
wire v$A24_17569_out1;
wire v$A24_17570_out0;
wire v$A24_17570_out1;
wire v$A24_17571_out0;
wire v$A24_17571_out1;
wire v$A24_17572_out0;
wire v$A24_17572_out1;
wire v$A24_17573_out0;
wire v$A24_17573_out1;
wire v$A24_17574_out0;
wire v$A24_17574_out1;
wire v$A2A_1788_out0;
wire v$A2A_1788_out1;
wire v$A2A_1789_out0;
wire v$A2A_1789_out1;
wire v$A2A_1790_out0;
wire v$A2A_1790_out1;
wire v$A2A_1791_out0;
wire v$A2A_1791_out1;
wire v$A2A_1792_out0;
wire v$A2A_1792_out1;
wire v$A2A_1793_out0;
wire v$A2A_1793_out1;
wire v$A2XNORB2_4659_out0;
wire v$A2XNORB2_4660_out0;
wire v$A2XNORB2_4661_out0;
wire v$A2XNORB2_4662_out0;
wire v$A2XNORB2_4663_out0;
wire v$A2XNORB2_4664_out0;
wire v$A2XNORB2_4665_out0;
wire v$A2XNORB2_4666_out0;
wire v$A2XNORB2_4667_out0;
wire v$A2XNORB2_4668_out0;
wire v$A2XNORB2_4669_out0;
wire v$A2XNORB2_4670_out0;
wire v$A2XNORB2_4671_out0;
wire v$A2XNORB2_4672_out0;
wire v$A2XNORB2_4673_out0;
wire v$A2XNORB2_4674_out0;
wire v$A2XNORB2_4675_out0;
wire v$A2XNORB2_4676_out0;
wire v$A2XNORB2_4677_out0;
wire v$A2XNORB2_4678_out0;
wire v$A2XNORB2_4679_out0;
wire v$A2XNORB2_4680_out0;
wire v$A2XNORB2_4681_out0;
wire v$A2XNORB2_4682_out0;
wire v$A2_10470_out1;
wire v$A2_10471_out1;
wire v$A2_10472_out1;
wire v$A2_10473_out1;
wire v$A2_15432_out1;
wire v$A2_15433_out1;
wire v$A2_18868_out0;
wire v$A2_18869_out0;
wire v$A2_18870_out0;
wire v$A2_18871_out0;
wire v$A2_18872_out0;
wire v$A2_18873_out0;
wire v$A2_8371_out0;
wire v$A2_8372_out0;
wire v$A2_8373_out0;
wire v$A2_8374_out0;
wire v$A2_8375_out0;
wire v$A2_8376_out0;
wire v$A2_8377_out0;
wire v$A2_8378_out0;
wire v$A2_8379_out0;
wire v$A2_8380_out0;
wire v$A2_8381_out0;
wire v$A2_8382_out0;
wire v$A2_8383_out0;
wire v$A2_8384_out0;
wire v$A2_8385_out0;
wire v$A2_8386_out0;
wire v$A2_8387_out0;
wire v$A2_8388_out0;
wire v$A2_8389_out0;
wire v$A2_8390_out0;
wire v$A2_8391_out0;
wire v$A2_8392_out0;
wire v$A2_8393_out0;
wire v$A2_8394_out0;
wire v$A3$COMP$B3_5160_out0;
wire v$A3$COMP$B3_5161_out0;
wire v$A3$COMP$B3_5162_out0;
wire v$A3$COMP$B3_5163_out0;
wire v$A3$COMP$B3_5164_out0;
wire v$A3$COMP$B3_5165_out0;
wire v$A3$COMP$B3_5166_out0;
wire v$A3$COMP$B3_5167_out0;
wire v$A3$COMP$B3_5168_out0;
wire v$A3$COMP$B3_5169_out0;
wire v$A3$COMP$B3_5170_out0;
wire v$A3$COMP$B3_5171_out0;
wire v$A3$COMP$B3_5172_out0;
wire v$A3$COMP$B3_5173_out0;
wire v$A3$COMP$B3_5174_out0;
wire v$A3$COMP$B3_5175_out0;
wire v$A3$COMP$B3_5176_out0;
wire v$A3$COMP$B3_5177_out0;
wire v$A3$COMP$B3_5178_out0;
wire v$A3$COMP$B3_5179_out0;
wire v$A3$COMP$B3_5180_out0;
wire v$A3$COMP$B3_5181_out0;
wire v$A3$COMP$B3_5182_out0;
wire v$A3$COMP$B3_5183_out0;
wire v$A3A_12525_out0;
wire v$A3A_12525_out1;
wire v$A3A_12526_out0;
wire v$A3A_12526_out1;
wire v$A3A_12527_out0;
wire v$A3A_12527_out1;
wire v$A3A_12528_out0;
wire v$A3A_12528_out1;
wire v$A3A_12529_out0;
wire v$A3A_12529_out1;
wire v$A3A_12530_out0;
wire v$A3A_12530_out1;
wire v$A3XNORB3_15323_out0;
wire v$A3XNORB3_15324_out0;
wire v$A3XNORB3_15325_out0;
wire v$A3XNORB3_15326_out0;
wire v$A3XNORB3_15327_out0;
wire v$A3XNORB3_15328_out0;
wire v$A3XNORB3_15329_out0;
wire v$A3XNORB3_15330_out0;
wire v$A3XNORB3_15331_out0;
wire v$A3XNORB3_15332_out0;
wire v$A3XNORB3_15333_out0;
wire v$A3XNORB3_15334_out0;
wire v$A3XNORB3_15335_out0;
wire v$A3XNORB3_15336_out0;
wire v$A3XNORB3_15337_out0;
wire v$A3XNORB3_15338_out0;
wire v$A3XNORB3_15339_out0;
wire v$A3XNORB3_15340_out0;
wire v$A3XNORB3_15341_out0;
wire v$A3XNORB3_15342_out0;
wire v$A3XNORB3_15343_out0;
wire v$A3XNORB3_15344_out0;
wire v$A3XNORB3_15345_out0;
wire v$A3XNORB3_15346_out0;
wire v$A3_11200_out0;
wire v$A3_11201_out0;
wire v$A3_11202_out0;
wire v$A3_11203_out0;
wire v$A3_11204_out0;
wire v$A3_11205_out0;
wire v$A3_11206_out0;
wire v$A3_11207_out0;
wire v$A3_11208_out0;
wire v$A3_11209_out0;
wire v$A3_11210_out0;
wire v$A3_11211_out0;
wire v$A3_11212_out0;
wire v$A3_11213_out0;
wire v$A3_11214_out0;
wire v$A3_11215_out0;
wire v$A3_11216_out0;
wire v$A3_11217_out0;
wire v$A3_11218_out0;
wire v$A3_11219_out0;
wire v$A3_11220_out0;
wire v$A3_11221_out0;
wire v$A3_11222_out0;
wire v$A3_11223_out0;
wire v$A3_15209_out0;
wire v$A3_15210_out0;
wire v$A3_15211_out0;
wire v$A3_15212_out0;
wire v$A3_15213_out0;
wire v$A3_15214_out0;
wire v$A4$COMP$B4_7725_out0;
wire v$A4$COMP$B4_7726_out0;
wire v$A4$COMP$B4_7727_out0;
wire v$A4$COMP$B4_7728_out0;
wire v$A4A_13731_out0;
wire v$A4A_13731_out1;
wire v$A4A_13732_out0;
wire v$A4A_13732_out1;
wire v$A4A_13733_out0;
wire v$A4A_13733_out1;
wire v$A4A_13734_out0;
wire v$A4A_13734_out1;
wire v$A4A_13735_out0;
wire v$A4A_13735_out1;
wire v$A4A_13736_out0;
wire v$A4A_13736_out1;
wire v$A4XNORB4_1535_out0;
wire v$A4XNORB4_1536_out0;
wire v$A4XNORB4_1537_out0;
wire v$A4XNORB4_1538_out0;
wire v$A4_15624_out0;
wire v$A4_15625_out0;
wire v$A4_15626_out0;
wire v$A4_15627_out0;
wire v$A4_18138_out0;
wire v$A4_18139_out0;
wire v$A4_18140_out0;
wire v$A4_18141_out0;
wire v$A4_18142_out0;
wire v$A4_18143_out0;
wire v$A5A_16709_out0;
wire v$A5A_16709_out1;
wire v$A5A_16710_out0;
wire v$A5A_16710_out1;
wire v$A5A_16711_out0;
wire v$A5A_16711_out1;
wire v$A5A_16712_out0;
wire v$A5A_16712_out1;
wire v$A5A_16713_out0;
wire v$A5A_16713_out1;
wire v$A5A_16714_out0;
wire v$A5A_16714_out1;
wire v$A5_6901_out0;
wire v$A5_6902_out0;
wire v$A5_6903_out0;
wire v$A5_6904_out0;
wire v$A5_6905_out0;
wire v$A5_6906_out0;
wire v$A6A_3334_out0;
wire v$A6A_3334_out1;
wire v$A6A_3335_out0;
wire v$A6A_3335_out1;
wire v$A6A_3336_out0;
wire v$A6A_3336_out1;
wire v$A6A_3337_out0;
wire v$A6A_3337_out1;
wire v$A6A_3338_out0;
wire v$A6A_3338_out1;
wire v$A6A_3339_out0;
wire v$A6A_3339_out1;
wire v$A6_320_out0;
wire v$A6_321_out0;
wire v$A6_322_out0;
wire v$A6_323_out0;
wire v$A6_324_out0;
wire v$A6_325_out0;
wire v$A7A_1815_out0;
wire v$A7A_1815_out1;
wire v$A7A_1816_out0;
wire v$A7A_1816_out1;
wire v$A7A_1817_out0;
wire v$A7A_1817_out1;
wire v$A7A_1818_out0;
wire v$A7A_1818_out1;
wire v$A7A_1819_out0;
wire v$A7A_1819_out1;
wire v$A7A_1820_out0;
wire v$A7A_1820_out1;
wire v$A7_15891_out0;
wire v$A7_15892_out0;
wire v$A7_15893_out0;
wire v$A7_15894_out0;
wire v$A7_15895_out0;
wire v$A7_15896_out0;
wire v$A8A_1659_out0;
wire v$A8A_1659_out1;
wire v$A8A_1660_out0;
wire v$A8A_1660_out1;
wire v$A8A_1661_out0;
wire v$A8A_1661_out1;
wire v$A8A_1662_out0;
wire v$A8A_1662_out1;
wire v$A8A_1663_out0;
wire v$A8A_1663_out1;
wire v$A8A_1664_out0;
wire v$A8A_1664_out1;
wire v$A8_18697_out0;
wire v$A8_18698_out0;
wire v$A8_18699_out0;
wire v$A8_18700_out0;
wire v$A8_18701_out0;
wire v$A8_18702_out0;
wire v$A9A_10862_out0;
wire v$A9A_10862_out1;
wire v$A9A_10863_out0;
wire v$A9A_10863_out1;
wire v$A9A_10864_out0;
wire v$A9A_10864_out1;
wire v$A9A_10865_out0;
wire v$A9A_10865_out1;
wire v$A9A_10866_out0;
wire v$A9A_10866_out1;
wire v$A9A_10867_out0;
wire v$A9A_10867_out1;
wire v$A9_3643_out0;
wire v$A9_3644_out0;
wire v$A9_3645_out0;
wire v$A9_3646_out0;
wire v$A9_3647_out0;
wire v$A9_3648_out0;
wire v$AD3$EQUALS$AD2_15156_out0;
wire v$AD3$EQUALS$AD2_15157_out0;
wire v$ADD_8527_out0;
wire v$ADD_8528_out0;
wire v$ARBHALT0_3114_out0;
wire v$ARBHALT1_5693_out0;
wire v$ARR0_11485_out0;
wire v$ARR1_9395_out0;
wire v$AUTODISABLE_18814_out0;
wire v$AUTODISABLE_18815_out0;
wire v$AWR0_1960_out0;
wire v$AWR1_16492_out0;
wire v$A_7391_out0;
wire v$A_7392_out0;
wire v$A_7393_out0;
wire v$A_7394_out0;
wire v$A_7395_out0;
wire v$A_7396_out0;
wire v$A_7397_out0;
wire v$A_7398_out0;
wire v$A_7399_out0;
wire v$A_7400_out0;
wire v$A_7401_out0;
wire v$A_7402_out0;
wire v$A_7403_out0;
wire v$A_7404_out0;
wire v$A_7405_out0;
wire v$A_7406_out0;
wire v$A_7407_out0;
wire v$A_7408_out0;
wire v$A_7409_out0;
wire v$A_7410_out0;
wire v$A_7411_out0;
wire v$A_7412_out0;
wire v$A_7413_out0;
wire v$A_7414_out0;
wire v$A_7415_out0;
wire v$A_7416_out0;
wire v$A_7417_out0;
wire v$A_7418_out0;
wire v$A_7419_out0;
wire v$A_7420_out0;
wire v$A_7421_out0;
wire v$A_7422_out0;
wire v$A_7423_out0;
wire v$A_7424_out0;
wire v$A_7425_out0;
wire v$A_7426_out0;
wire v$A_7427_out0;
wire v$A_7428_out0;
wire v$A_7429_out0;
wire v$A_7430_out0;
wire v$A_7431_out0;
wire v$A_7432_out0;
wire v$A_7433_out0;
wire v$A_7434_out0;
wire v$A_7435_out0;
wire v$A_7436_out0;
wire v$A_7437_out0;
wire v$A_7438_out0;
wire v$A_7439_out0;
wire v$A_7440_out0;
wire v$A_7441_out0;
wire v$A_7442_out0;
wire v$A_7443_out0;
wire v$A_7444_out0;
wire v$A_7445_out0;
wire v$A_7446_out0;
wire v$A_7447_out0;
wire v$A_7448_out0;
wire v$A_7449_out0;
wire v$A_7450_out0;
wire v$A_7451_out0;
wire v$A_7452_out0;
wire v$A_7453_out0;
wire v$A_7454_out0;
wire v$A_7455_out0;
wire v$A_7456_out0;
wire v$A_7457_out0;
wire v$A_7458_out0;
wire v$A_7459_out0;
wire v$A_7460_out0;
wire v$A_7461_out0;
wire v$A_7462_out0;
wire v$A_7463_out0;
wire v$A_7464_out0;
wire v$A_7465_out0;
wire v$A_7466_out0;
wire v$A_7467_out0;
wire v$A_7468_out0;
wire v$A_7469_out0;
wire v$A_7470_out0;
wire v$A_7471_out0;
wire v$A_7472_out0;
wire v$A_7473_out0;
wire v$A_7474_out0;
wire v$A_7475_out0;
wire v$A_7476_out0;
wire v$A_7477_out0;
wire v$A_7478_out0;
wire v$A_7479_out0;
wire v$A_7480_out0;
wire v$A_7481_out0;
wire v$A_7482_out0;
wire v$A_7483_out0;
wire v$A_7484_out0;
wire v$A_7485_out0;
wire v$A_7486_out0;
wire v$A_7487_out0;
wire v$A_7488_out0;
wire v$A_7489_out0;
wire v$A_7490_out0;
wire v$A_7491_out0;
wire v$A_7492_out0;
wire v$A_7493_out0;
wire v$A_7494_out0;
wire v$A_7495_out0;
wire v$A_7496_out0;
wire v$A_7497_out0;
wire v$A_7498_out0;
wire v$A_7499_out0;
wire v$A_7500_out0;
wire v$A_7501_out0;
wire v$A_7502_out0;
wire v$A_7503_out0;
wire v$A_7504_out0;
wire v$A_7505_out0;
wire v$A_7506_out0;
wire v$A_7507_out0;
wire v$A_7508_out0;
wire v$A_7509_out0;
wire v$A_7510_out0;
wire v$A_7511_out0;
wire v$A_7512_out0;
wire v$A_7513_out0;
wire v$A_7514_out0;
wire v$A_7515_out0;
wire v$A_7516_out0;
wire v$A_7517_out0;
wire v$A_7518_out0;
wire v$A_7519_out0;
wire v$A_7520_out0;
wire v$A_7521_out0;
wire v$A_7522_out0;
wire v$A_7523_out0;
wire v$A_7524_out0;
wire v$A_7525_out0;
wire v$A_7526_out0;
wire v$A_7527_out0;
wire v$A_7528_out0;
wire v$A_7529_out0;
wire v$A_7530_out0;
wire v$A_7531_out0;
wire v$A_7532_out0;
wire v$A_7533_out0;
wire v$A_7534_out0;
wire v$B$IS$RD_14695_out0;
wire v$B$IS$RD_14696_out0;
wire v$B0_3421_out0;
wire v$B0_3422_out0;
wire v$B0_3423_out0;
wire v$B0_3424_out0;
wire v$B0_3425_out0;
wire v$B0_3426_out0;
wire v$B0_3836_out0;
wire v$B0_3837_out0;
wire v$B0_3838_out0;
wire v$B0_3839_out0;
wire v$B0_3840_out0;
wire v$B0_3841_out0;
wire v$B0_3842_out0;
wire v$B0_3843_out0;
wire v$B0_3844_out0;
wire v$B0_3845_out0;
wire v$B0_3846_out0;
wire v$B0_3847_out0;
wire v$B0_3848_out0;
wire v$B0_3849_out0;
wire v$B0_3850_out0;
wire v$B0_3851_out0;
wire v$B0_3852_out0;
wire v$B0_3853_out0;
wire v$B0_3854_out0;
wire v$B0_3855_out0;
wire v$B0_3856_out0;
wire v$B0_3857_out0;
wire v$B0_3858_out0;
wire v$B0_3859_out0;
wire v$B10_10297_out0;
wire v$B10_10298_out0;
wire v$B10_10299_out0;
wire v$B10_10300_out0;
wire v$B10_10301_out0;
wire v$B10_10302_out0;
wire v$B11_9443_out0;
wire v$B11_9444_out0;
wire v$B11_9445_out0;
wire v$B11_9446_out0;
wire v$B11_9447_out0;
wire v$B11_9448_out0;
wire v$B12_2114_out0;
wire v$B12_2115_out0;
wire v$B12_2116_out0;
wire v$B12_2117_out0;
wire v$B12_2118_out0;
wire v$B12_2119_out0;
wire v$B13_9022_out0;
wire v$B13_9023_out0;
wire v$B13_9024_out0;
wire v$B13_9025_out0;
wire v$B13_9026_out0;
wire v$B13_9027_out0;
wire v$B14_4158_out0;
wire v$B14_4159_out0;
wire v$B14_4160_out0;
wire v$B14_4161_out0;
wire v$B14_4162_out0;
wire v$B14_4163_out0;
wire v$B15_10446_out0;
wire v$B15_10447_out0;
wire v$B15_10448_out0;
wire v$B15_10449_out0;
wire v$B15_10450_out0;
wire v$B15_10451_out0;
wire v$B16_17034_out0;
wire v$B16_17035_out0;
wire v$B16_17036_out0;
wire v$B16_17037_out0;
wire v$B16_17038_out0;
wire v$B16_17039_out0;
wire v$B17_16125_out0;
wire v$B17_16126_out0;
wire v$B17_16127_out0;
wire v$B17_16128_out0;
wire v$B17_16129_out0;
wire v$B17_16130_out0;
wire v$B18_11368_out0;
wire v$B18_11369_out0;
wire v$B18_11370_out0;
wire v$B18_11371_out0;
wire v$B18_11372_out0;
wire v$B18_11373_out0;
wire v$B19_17410_out0;
wire v$B19_17411_out0;
wire v$B19_17412_out0;
wire v$B19_17413_out0;
wire v$B19_17414_out0;
wire v$B19_17415_out0;
wire v$B1_14822_out0;
wire v$B1_14823_out0;
wire v$B1_14824_out0;
wire v$B1_14825_out0;
wire v$B1_14826_out0;
wire v$B1_14827_out0;
wire v$B1_14828_out0;
wire v$B1_14829_out0;
wire v$B1_14830_out0;
wire v$B1_14831_out0;
wire v$B1_14832_out0;
wire v$B1_14833_out0;
wire v$B1_14834_out0;
wire v$B1_14835_out0;
wire v$B1_14836_out0;
wire v$B1_14837_out0;
wire v$B1_14838_out0;
wire v$B1_14839_out0;
wire v$B1_14840_out0;
wire v$B1_14841_out0;
wire v$B1_14842_out0;
wire v$B1_14843_out0;
wire v$B1_14844_out0;
wire v$B1_14845_out0;
wire v$B1_8426_out0;
wire v$B1_8427_out0;
wire v$B1_8428_out0;
wire v$B1_8429_out0;
wire v$B1_8430_out0;
wire v$B1_8431_out0;
wire v$B20_4112_out0;
wire v$B20_4113_out0;
wire v$B20_4114_out0;
wire v$B20_4115_out0;
wire v$B20_4116_out0;
wire v$B20_4117_out0;
wire v$B21_18689_out0;
wire v$B21_18690_out0;
wire v$B21_18691_out0;
wire v$B21_18692_out0;
wire v$B21_18693_out0;
wire v$B21_18694_out0;
wire v$B22_11300_out0;
wire v$B22_11301_out0;
wire v$B22_11302_out0;
wire v$B22_11303_out0;
wire v$B22_11304_out0;
wire v$B22_11305_out0;
wire v$B23_1441_out0;
wire v$B23_1442_out0;
wire v$B23_1443_out0;
wire v$B23_1444_out0;
wire v$B23_1445_out0;
wire v$B23_1446_out0;
wire v$B2_17244_out0;
wire v$B2_17245_out0;
wire v$B2_17246_out0;
wire v$B2_17247_out0;
wire v$B2_17248_out0;
wire v$B2_17249_out0;
wire v$B2_17250_out0;
wire v$B2_17251_out0;
wire v$B2_17252_out0;
wire v$B2_17253_out0;
wire v$B2_17254_out0;
wire v$B2_17255_out0;
wire v$B2_17256_out0;
wire v$B2_17257_out0;
wire v$B2_17258_out0;
wire v$B2_17259_out0;
wire v$B2_17260_out0;
wire v$B2_17261_out0;
wire v$B2_17262_out0;
wire v$B2_17263_out0;
wire v$B2_17264_out0;
wire v$B2_17265_out0;
wire v$B2_17266_out0;
wire v$B2_17267_out0;
wire v$B2_3326_out0;
wire v$B2_3327_out0;
wire v$B2_3328_out0;
wire v$B2_3329_out0;
wire v$B2_3330_out0;
wire v$B2_3331_out0;
wire v$B3_18460_out0;
wire v$B3_18461_out0;
wire v$B3_18462_out0;
wire v$B3_18463_out0;
wire v$B3_18464_out0;
wire v$B3_18465_out0;
wire v$B3_18466_out0;
wire v$B3_18467_out0;
wire v$B3_18468_out0;
wire v$B3_18469_out0;
wire v$B3_18470_out0;
wire v$B3_18471_out0;
wire v$B3_18472_out0;
wire v$B3_18473_out0;
wire v$B3_18474_out0;
wire v$B3_18475_out0;
wire v$B3_18476_out0;
wire v$B3_18477_out0;
wire v$B3_18478_out0;
wire v$B3_18479_out0;
wire v$B3_18480_out0;
wire v$B3_18481_out0;
wire v$B3_18482_out0;
wire v$B3_18483_out0;
wire v$B3_9845_out0;
wire v$B3_9846_out0;
wire v$B3_9847_out0;
wire v$B3_9848_out0;
wire v$B3_9849_out0;
wire v$B3_9850_out0;
wire v$B4_15266_out0;
wire v$B4_15267_out0;
wire v$B4_15268_out0;
wire v$B4_15269_out0;
wire v$B4_15270_out0;
wire v$B4_15271_out0;
wire v$B4_17533_out0;
wire v$B4_17534_out0;
wire v$B4_17535_out0;
wire v$B4_17536_out0;
wire v$B5_18978_out0;
wire v$B5_18979_out0;
wire v$B5_18980_out0;
wire v$B5_18981_out0;
wire v$B5_18982_out0;
wire v$B5_18983_out0;
wire v$B6_13883_out0;
wire v$B6_13884_out0;
wire v$B6_13885_out0;
wire v$B6_13886_out0;
wire v$B6_13887_out0;
wire v$B6_13888_out0;
wire v$B7_17634_out0;
wire v$B7_17635_out0;
wire v$B7_17636_out0;
wire v$B7_17637_out0;
wire v$B7_17638_out0;
wire v$B7_17639_out0;
wire v$B8_13715_out0;
wire v$B8_13716_out0;
wire v$B8_13717_out0;
wire v$B8_13718_out0;
wire v$B8_13719_out0;
wire v$B8_13720_out0;
wire v$B9_4220_out0;
wire v$B9_4221_out0;
wire v$B9_4222_out0;
wire v$B9_4223_out0;
wire v$B9_4224_out0;
wire v$B9_4225_out0;
wire v$B_2896_out0;
wire v$B_2897_out0;
wire v$B_2898_out0;
wire v$B_2899_out0;
wire v$B_2900_out0;
wire v$B_2901_out0;
wire v$B_2902_out0;
wire v$B_2903_out0;
wire v$B_2904_out0;
wire v$B_2905_out0;
wire v$B_2906_out0;
wire v$B_2907_out0;
wire v$B_2908_out0;
wire v$B_2909_out0;
wire v$B_2910_out0;
wire v$B_2911_out0;
wire v$B_2912_out0;
wire v$B_2913_out0;
wire v$B_2914_out0;
wire v$B_2915_out0;
wire v$B_2916_out0;
wire v$B_2917_out0;
wire v$B_2918_out0;
wire v$B_2919_out0;
wire v$B_2920_out0;
wire v$B_2921_out0;
wire v$B_2922_out0;
wire v$B_2923_out0;
wire v$B_2924_out0;
wire v$B_2925_out0;
wire v$B_2926_out0;
wire v$B_2927_out0;
wire v$B_2928_out0;
wire v$B_2929_out0;
wire v$B_2930_out0;
wire v$B_2931_out0;
wire v$B_2932_out0;
wire v$B_2933_out0;
wire v$B_2934_out0;
wire v$B_2935_out0;
wire v$B_2936_out0;
wire v$B_2937_out0;
wire v$B_2938_out0;
wire v$B_2939_out0;
wire v$B_2940_out0;
wire v$B_2941_out0;
wire v$B_2942_out0;
wire v$B_2943_out0;
wire v$B_2944_out0;
wire v$B_2945_out0;
wire v$B_2946_out0;
wire v$B_2947_out0;
wire v$B_2948_out0;
wire v$B_2949_out0;
wire v$B_2950_out0;
wire v$B_2951_out0;
wire v$B_2952_out0;
wire v$B_2953_out0;
wire v$B_2954_out0;
wire v$B_2955_out0;
wire v$B_2956_out0;
wire v$B_2957_out0;
wire v$B_2958_out0;
wire v$B_2959_out0;
wire v$B_2960_out0;
wire v$B_2961_out0;
wire v$B_2962_out0;
wire v$B_2963_out0;
wire v$B_2964_out0;
wire v$B_2965_out0;
wire v$B_2966_out0;
wire v$B_2967_out0;
wire v$B_2968_out0;
wire v$B_2969_out0;
wire v$B_2970_out0;
wire v$B_2971_out0;
wire v$B_2972_out0;
wire v$B_2973_out0;
wire v$B_2974_out0;
wire v$B_2975_out0;
wire v$B_2976_out0;
wire v$B_2977_out0;
wire v$B_2978_out0;
wire v$B_2979_out0;
wire v$B_2980_out0;
wire v$B_2981_out0;
wire v$B_2982_out0;
wire v$B_2983_out0;
wire v$B_2984_out0;
wire v$B_2985_out0;
wire v$B_2986_out0;
wire v$B_2987_out0;
wire v$B_2988_out0;
wire v$B_2989_out0;
wire v$B_2990_out0;
wire v$B_2991_out0;
wire v$B_2992_out0;
wire v$B_2993_out0;
wire v$B_2994_out0;
wire v$B_2995_out0;
wire v$B_2996_out0;
wire v$B_2997_out0;
wire v$B_2998_out0;
wire v$B_2999_out0;
wire v$B_3000_out0;
wire v$B_3001_out0;
wire v$B_3002_out0;
wire v$B_3003_out0;
wire v$B_3004_out0;
wire v$B_3005_out0;
wire v$B_3006_out0;
wire v$B_3007_out0;
wire v$B_3008_out0;
wire v$B_3009_out0;
wire v$B_3010_out0;
wire v$B_3011_out0;
wire v$B_3012_out0;
wire v$B_3013_out0;
wire v$B_3014_out0;
wire v$B_3015_out0;
wire v$B_3016_out0;
wire v$B_3017_out0;
wire v$B_3018_out0;
wire v$B_3019_out0;
wire v$B_3020_out0;
wire v$B_3021_out0;
wire v$B_3022_out0;
wire v$B_3023_out0;
wire v$B_3024_out0;
wire v$B_3025_out0;
wire v$B_3026_out0;
wire v$B_3027_out0;
wire v$B_3028_out0;
wire v$B_3029_out0;
wire v$B_3030_out0;
wire v$B_3031_out0;
wire v$B_3032_out0;
wire v$B_3033_out0;
wire v$B_3034_out0;
wire v$B_3035_out0;
wire v$B_3036_out0;
wire v$B_3037_out0;
wire v$B_3038_out0;
wire v$B_3039_out0;
wire v$C0_11188_out0;
wire v$C0_11189_out0;
wire v$C0_11190_out0;
wire v$C0_11191_out0;
wire v$C0_11192_out0;
wire v$C0_11193_out0;
wire v$C0_9745_out0;
wire v$C0_9746_out0;
wire v$C0_9747_out0;
wire v$C0_9748_out0;
wire v$C0_9749_out0;
wire v$C0_9750_out0;
wire v$C10_13301_out0;
wire v$C10_13302_out0;
wire v$C10_13303_out0;
wire v$C10_13304_out0;
wire v$C10_13305_out0;
wire v$C10_13306_out0;
wire v$C10_2103_out0;
wire v$C10_2104_out0;
wire v$C10_2105_out0;
wire v$C10_2106_out0;
wire v$C10_2107_out0;
wire v$C10_2108_out0;
wire v$C11_15404_out0;
wire v$C11_15405_out0;
wire v$C11_15406_out0;
wire v$C11_15407_out0;
wire v$C11_15408_out0;
wire v$C11_15409_out0;
wire v$C11_3822_out0;
wire v$C11_3823_out0;
wire v$C11_9887_out0;
wire v$C11_9888_out0;
wire v$C11_9889_out0;
wire v$C11_9890_out0;
wire v$C11_9891_out0;
wire v$C11_9892_out0;
wire v$C12_14094_out0;
wire v$C12_14095_out0;
wire v$C12_14096_out0;
wire v$C12_14097_out0;
wire v$C12_14098_out0;
wire v$C12_14099_out0;
wire v$C12_9767_out0;
wire v$C12_9768_out0;
wire v$C12_9769_out0;
wire v$C12_9770_out0;
wire v$C12_9771_out0;
wire v$C12_9772_out0;
wire v$C13_12346_out0;
wire v$C13_12347_out0;
wire v$C13_12348_out0;
wire v$C13_12349_out0;
wire v$C13_12350_out0;
wire v$C13_12351_out0;
wire v$C13_19197_out0;
wire v$C13_19198_out0;
wire v$C13_19199_out0;
wire v$C13_19200_out0;
wire v$C13_19201_out0;
wire v$C13_19202_out0;
wire v$C14_290_out0;
wire v$C14_291_out0;
wire v$C14_292_out0;
wire v$C14_293_out0;
wire v$C14_294_out0;
wire v$C14_295_out0;
wire v$C14_340_out0;
wire v$C14_341_out0;
wire v$C14_342_out0;
wire v$C14_343_out0;
wire v$C14_344_out0;
wire v$C14_345_out0;
wire v$C15_13707_out0;
wire v$C15_13708_out0;
wire v$C15_13709_out0;
wire v$C15_13710_out0;
wire v$C15_13711_out0;
wire v$C15_13712_out0;
wire v$C15_8447_out0;
wire v$C15_8448_out0;
wire v$C15_8449_out0;
wire v$C15_8450_out0;
wire v$C15_8451_out0;
wire v$C15_8452_out0;
wire v$C16_1423_out0;
wire v$C16_1424_out0;
wire v$C16_1425_out0;
wire v$C16_1426_out0;
wire v$C16_1427_out0;
wire v$C16_1428_out0;
wire v$C16_15768_out0;
wire v$C16_15769_out0;
wire v$C16_15770_out0;
wire v$C16_15771_out0;
wire v$C16_15772_out0;
wire v$C16_15773_out0;
wire v$C17_2716_out0;
wire v$C17_2717_out0;
wire v$C17_2718_out0;
wire v$C17_2719_out0;
wire v$C17_2720_out0;
wire v$C17_2721_out0;
wire v$C17_6342_out0;
wire v$C17_6343_out0;
wire v$C17_6344_out0;
wire v$C17_6345_out0;
wire v$C17_6346_out0;
wire v$C17_6347_out0;
wire v$C18_16902_out0;
wire v$C18_16903_out0;
wire v$C18_16904_out0;
wire v$C18_16905_out0;
wire v$C18_16906_out0;
wire v$C18_16907_out0;
wire v$C18_18609_out0;
wire v$C18_18610_out0;
wire v$C18_18611_out0;
wire v$C18_18612_out0;
wire v$C18_18613_out0;
wire v$C18_18614_out0;
wire v$C19_14421_out0;
wire v$C19_14422_out0;
wire v$C19_14423_out0;
wire v$C19_14424_out0;
wire v$C19_14425_out0;
wire v$C19_14426_out0;
wire v$C19_8467_out0;
wire v$C19_8468_out0;
wire v$C19_8469_out0;
wire v$C19_8470_out0;
wire v$C19_8471_out0;
wire v$C19_8472_out0;
wire v$C1_12421_out0;
wire v$C1_12422_out0;
wire v$C1_12423_out0;
wire v$C1_12424_out0;
wire v$C1_12425_out0;
wire v$C1_12426_out0;
wire v$C1_13423_out0;
wire v$C1_13424_out0;
wire v$C1_14639_out0;
wire v$C1_14640_out0;
wire v$C1_1623_out0;
wire v$C1_1624_out0;
wire v$C1_16317_out0;
wire v$C1_16318_out0;
wire v$C1_16319_out0;
wire v$C1_16320_out0;
wire v$C1_16526_out0;
wire v$C1_16527_out0;
wire v$C1_1669_out0;
wire v$C1_1670_out0;
wire v$C1_17401_out0;
wire v$C1_17402_out0;
wire v$C1_17403_out0;
wire v$C1_17404_out0;
wire v$C1_17405_out0;
wire v$C1_17406_out0;
wire v$C1_17979_out0;
wire v$C1_17980_out0;
wire v$C1_17981_out0;
wire v$C1_17982_out0;
wire v$C1_18266_out0;
wire v$C1_18267_out0;
wire v$C1_18268_out0;
wire v$C1_18269_out0;
wire v$C1_18270_out0;
wire v$C1_18271_out0;
wire v$C1_18272_out0;
wire v$C1_18273_out0;
wire v$C1_18274_out0;
wire v$C1_18275_out0;
wire v$C1_2830_out0;
wire v$C1_2831_out0;
wire v$C1_2832_out0;
wire v$C1_2833_out0;
wire v$C1_2834_out0;
wire v$C1_2835_out0;
wire v$C1_2836_out0;
wire v$C1_2837_out0;
wire v$C1_2838_out0;
wire v$C1_2839_out0;
wire v$C1_2840_out0;
wire v$C1_2841_out0;
wire v$C1_4520_out0;
wire v$C1_4521_out0;
wire v$C1_4633_out0;
wire v$C1_4634_out0;
wire v$C1_4635_out0;
wire v$C1_4636_out0;
wire v$C1_4637_out0;
wire v$C1_4638_out0;
wire v$C1_5674_out0;
wire v$C1_5675_out0;
wire v$C1_6244_out0;
wire v$C1_6249_out0;
wire v$C1_6254_out0;
wire v$C1_6257_out0;
wire v$C1_6264_out0;
wire v$C1_6267_out0;
wire v$C1_6272_out0;
wire v$C1_6275_out0;
wire v$C1_6280_out0;
wire v$C1_6285_out0;
wire v$C1_6288_out0;
wire v$C1_6295_out0;
wire v$C1_6298_out0;
wire v$C1_6303_out0;
wire v$C1_6703_out0;
wire v$C1_6704_out0;
wire v$C1_8287_out0;
wire v$C1_8291_out0;
wire v$C20_15592_out0;
wire v$C20_15593_out0;
wire v$C20_15594_out0;
wire v$C20_15595_out0;
wire v$C20_15596_out0;
wire v$C20_15597_out0;
wire v$C20_16079_out0;
wire v$C20_16080_out0;
wire v$C20_16081_out0;
wire v$C20_16082_out0;
wire v$C20_16083_out0;
wire v$C20_16084_out0;
wire v$C21_11258_out0;
wire v$C21_11259_out0;
wire v$C21_11260_out0;
wire v$C21_11261_out0;
wire v$C21_11262_out0;
wire v$C21_11263_out0;
wire v$C21_6608_out0;
wire v$C21_6609_out0;
wire v$C21_6610_out0;
wire v$C21_6611_out0;
wire v$C21_6612_out0;
wire v$C21_6613_out0;
wire v$C22_11488_out0;
wire v$C22_11489_out0;
wire v$C22_11490_out0;
wire v$C22_11491_out0;
wire v$C22_11492_out0;
wire v$C22_11493_out0;
wire v$C22_8714_out0;
wire v$C22_8715_out0;
wire v$C22_8716_out0;
wire v$C22_8717_out0;
wire v$C22_8718_out0;
wire v$C22_8719_out0;
wire v$C23_16758_out0;
wire v$C23_16759_out0;
wire v$C23_16760_out0;
wire v$C23_16761_out0;
wire v$C23_16762_out0;
wire v$C23_16763_out0;
wire v$C23_5056_out0;
wire v$C23_5057_out0;
wire v$C23_5058_out0;
wire v$C23_5059_out0;
wire v$C23_5060_out0;
wire v$C23_5061_out0;
wire v$C2_106_out0;
wire v$C2_11198_out0;
wire v$C2_11199_out0;
wire v$C2_111_out0;
wire v$C2_116_out0;
wire v$C2_119_out0;
wire v$C2_126_out0;
wire v$C2_129_out0;
wire v$C2_1317_out0;
wire v$C2_1318_out0;
wire v$C2_134_out0;
wire v$C2_137_out0;
wire v$C2_14082_out0;
wire v$C2_14083_out0;
wire v$C2_142_out0;
wire v$C2_147_out0;
wire v$C2_150_out0;
wire v$C2_15778_out0;
wire v$C2_15779_out0;
wire v$C2_15780_out0;
wire v$C2_15781_out0;
wire v$C2_157_out0;
wire v$C2_1607_out0;
wire v$C2_1608_out0;
wire v$C2_160_out0;
wire v$C2_165_out0;
wire v$C2_16851_out0;
wire v$C2_16852_out0;
wire v$C2_16894_out0;
wire v$C2_16895_out0;
wire v$C2_16896_out0;
wire v$C2_16897_out0;
wire v$C2_16946_out0;
wire v$C2_16947_out0;
wire v$C2_16948_out0;
wire v$C2_16949_out0;
wire v$C2_17614_out0;
wire v$C2_17615_out0;
wire v$C2_18777_out0;
wire v$C2_18778_out0;
wire v$C2_18779_out0;
wire v$C2_18780_out0;
wire v$C2_18781_out0;
wire v$C2_18782_out0;
wire v$C2_18926_out0;
wire v$C2_18927_out0;
wire v$C2_2863_out0;
wire v$C2_2864_out0;
wire v$C2_2884_out0;
wire v$C2_2885_out0;
wire v$C2_2886_out0;
wire v$C2_2887_out0;
wire v$C2_2888_out0;
wire v$C2_2889_out0;
wire v$C2_3185_out0;
wire v$C2_3186_out0;
wire v$C2_3818_out0;
wire v$C2_3819_out0;
wire v$C2_7951_out0;
wire v$C2_7952_out0;
wire v$C2_7953_out0;
wire v$C2_7954_out0;
wire v$C2_7955_out0;
wire v$C2_7956_out0;
wire v$C2_7957_out0;
wire v$C2_7958_out0;
wire v$C2_7959_out0;
wire v$C2_7960_out0;
wire v$C3_14090_out0;
wire v$C3_14091_out0;
wire v$C3_14092_out0;
wire v$C3_14093_out0;
wire v$C3_1525_out0;
wire v$C3_1526_out0;
wire v$C3_16323_out0;
wire v$C3_16324_out0;
wire v$C3_16325_out0;
wire v$C3_16326_out0;
wire v$C3_16327_out0;
wire v$C3_16328_out0;
wire v$C3_16420_out0;
wire v$C3_16421_out0;
wire v$C3_16422_out0;
wire v$C3_16423_out0;
wire v$C3_16424_out0;
wire v$C3_16425_out0;
wire v$C3_18739_out0;
wire v$C3_18740_out0;
wire v$C3_19163_out0;
wire v$C3_19164_out0;
wire v$C3_5628_out0;
wire v$C3_5629_out0;
wire v$C4_1413_out0;
wire v$C4_1414_out0;
wire v$C4_1415_out0;
wire v$C4_1416_out0;
wire v$C4_1417_out0;
wire v$C4_1418_out0;
wire v$C4_15440_out0;
wire v$C4_15441_out0;
wire v$C4_15442_out0;
wire v$C4_15443_out0;
wire v$C4_2038_out0;
wire v$C4_2039_out0;
wire v$C4_2040_out0;
wire v$C4_2041_out0;
wire v$C4_2042_out0;
wire v$C4_2043_out0;
wire v$C4_3127_out0;
wire v$C4_3128_out0;
wire v$C4_3935_out0;
wire v$C4_3936_out0;
wire v$C4_6606_out0;
wire v$C4_6607_out0;
wire v$C5_12253_out0;
wire v$C5_12254_out0;
wire v$C5_12255_out0;
wire v$C5_12256_out0;
wire v$C5_12257_out0;
wire v$C5_12258_out0;
wire v$C5_16519_out0;
wire v$C5_16520_out0;
wire v$C5_16521_out0;
wire v$C5_16522_out0;
wire v$C5_16523_out0;
wire v$C5_16524_out0;
wire v$C5_16705_out0;
wire v$C5_16706_out0;
wire v$C5_17519_out0;
wire v$C5_17521_out0;
wire v$C5_17523_out0;
wire v$C5_17525_out0;
wire v$C5_9112_out0;
wire v$C5_9113_out0;
wire v$C5_9114_out0;
wire v$C5_9115_out0;
wire v$C6_13145_out0;
wire v$C6_13146_out0;
wire v$C6_1725_out0;
wire v$C6_1726_out0;
wire v$C6_7341_out0;
wire v$C6_7342_out0;
wire v$C6_7343_out0;
wire v$C6_7344_out0;
wire v$C6_7345_out0;
wire v$C6_7346_out0;
wire v$C6_9182_out0;
wire v$C6_9183_out0;
wire v$C6_9966_out0;
wire v$C6_9967_out0;
wire v$C6_9968_out0;
wire v$C6_9969_out0;
wire v$C6_9970_out0;
wire v$C6_9971_out0;
wire v$C7_11475_out0;
wire v$C7_11476_out0;
wire v$C7_11477_out0;
wire v$C7_11478_out0;
wire v$C7_11479_out0;
wire v$C7_11480_out0;
wire v$C7_17051_out0;
wire v$C7_17052_out0;
wire v$C7_17053_out0;
wire v$C7_17054_out0;
wire v$C7_17055_out0;
wire v$C7_17056_out0;
wire v$C7_354_out0;
wire v$C7_355_out0;
wire v$C7_9871_out0;
wire v$C7_9872_out0;
wire v$C8_19107_out0;
wire v$C8_19108_out0;
wire v$C8_19109_out0;
wire v$C8_19110_out0;
wire v$C8_19111_out0;
wire v$C8_19112_out0;
wire v$C8_7748_out0;
wire v$C8_7749_out0;
wire v$C8_7750_out0;
wire v$C8_7751_out0;
wire v$C8_7752_out0;
wire v$C8_7753_out0;
wire v$C9_12716_out0;
wire v$C9_12717_out0;
wire v$C9_12718_out0;
wire v$C9_12719_out0;
wire v$C9_12720_out0;
wire v$C9_12721_out0;
wire v$C9_6216_out0;
wire v$C9_6217_out0;
wire v$C9_6218_out0;
wire v$C9_6219_out0;
wire v$C9_6220_out0;
wire v$C9_6221_out0;
wire v$CALCULATING_1647_out0;
wire v$CALCULATING_1648_out0;
wire v$CALCULATING_8122_out0;
wire v$CALCULATING_8123_out0;
wire v$CAPTURE_251_out0;
wire v$CAPTURE_252_out0;
wire v$CARRY_11411_out0;
wire v$CARRY_11412_out0;
wire v$CARRY_14027_out0;
wire v$CARRY_14028_out0;
wire v$CARRY_5219_out0;
wire v$CARRY_5220_out0;
wire v$CARRY_6582_out0;
wire v$CARRY_6583_out0;
wire v$CARRY_6584_out0;
wire v$CARRY_6585_out0;
wire v$CARRY_6586_out0;
wire v$CARRY_6587_out0;
wire v$CHECKPARITY_1489_out0;
wire v$CHECKPARITY_1490_out0;
wire v$CINA_8770_out0;
wire v$CINA_8771_out0;
wire v$CINA_8772_out0;
wire v$CINA_8773_out0;
wire v$CINA_8774_out0;
wire v$CINA_8775_out0;
wire v$CINA_8776_out0;
wire v$CINA_8777_out0;
wire v$CINA_8778_out0;
wire v$CINA_8779_out0;
wire v$CINA_8780_out0;
wire v$CINA_8781_out0;
wire v$CINA_8782_out0;
wire v$CINA_8783_out0;
wire v$CINA_8784_out0;
wire v$CINA_8785_out0;
wire v$CINA_8786_out0;
wire v$CINA_8787_out0;
wire v$CINA_8788_out0;
wire v$CINA_8789_out0;
wire v$CINA_8790_out0;
wire v$CINA_8791_out0;
wire v$CINA_8792_out0;
wire v$CINA_8793_out0;
wire v$CINA_8794_out0;
wire v$CINA_8795_out0;
wire v$CINA_8796_out0;
wire v$CINA_8797_out0;
wire v$CINA_8798_out0;
wire v$CINA_8799_out0;
wire v$CINA_8800_out0;
wire v$CINA_8801_out0;
wire v$CINA_8802_out0;
wire v$CINA_8803_out0;
wire v$CINA_8804_out0;
wire v$CINA_8805_out0;
wire v$CINA_8806_out0;
wire v$CINA_8807_out0;
wire v$CINA_8808_out0;
wire v$CINA_8809_out0;
wire v$CINA_8810_out0;
wire v$CINA_8811_out0;
wire v$CINA_8812_out0;
wire v$CINA_8813_out0;
wire v$CINA_8814_out0;
wire v$CINA_8815_out0;
wire v$CINA_8816_out0;
wire v$CINA_8817_out0;
wire v$CINA_8818_out0;
wire v$CINA_8819_out0;
wire v$CINA_8820_out0;
wire v$CINA_8821_out0;
wire v$CINA_8822_out0;
wire v$CINA_8823_out0;
wire v$CINA_8824_out0;
wire v$CINA_8825_out0;
wire v$CINA_8826_out0;
wire v$CINA_8827_out0;
wire v$CINA_8828_out0;
wire v$CINA_8829_out0;
wire v$CINA_8830_out0;
wire v$CINA_8831_out0;
wire v$CINA_8832_out0;
wire v$CINA_8833_out0;
wire v$CINA_8834_out0;
wire v$CINA_8835_out0;
wire v$CINA_8836_out0;
wire v$CINA_8837_out0;
wire v$CINA_8838_out0;
wire v$CINA_8839_out0;
wire v$CINA_8840_out0;
wire v$CINA_8841_out0;
wire v$CINA_8842_out0;
wire v$CINA_8843_out0;
wire v$CINA_8844_out0;
wire v$CINA_8845_out0;
wire v$CINA_8846_out0;
wire v$CINA_8847_out0;
wire v$CINA_8848_out0;
wire v$CINA_8849_out0;
wire v$CINA_8850_out0;
wire v$CINA_8851_out0;
wire v$CINA_8852_out0;
wire v$CINA_8853_out0;
wire v$CINA_8854_out0;
wire v$CINA_8855_out0;
wire v$CINA_8856_out0;
wire v$CINA_8857_out0;
wire v$CINA_8858_out0;
wire v$CINA_8859_out0;
wire v$CINA_8860_out0;
wire v$CINA_8861_out0;
wire v$CINA_8862_out0;
wire v$CINA_8863_out0;
wire v$CINA_8864_out0;
wire v$CINA_8865_out0;
wire v$CINA_8866_out0;
wire v$CINA_8867_out0;
wire v$CINA_8868_out0;
wire v$CINA_8869_out0;
wire v$CINA_8870_out0;
wire v$CINA_8871_out0;
wire v$CINA_8872_out0;
wire v$CINA_8873_out0;
wire v$CINA_8874_out0;
wire v$CINA_8875_out0;
wire v$CINA_8876_out0;
wire v$CINA_8877_out0;
wire v$CINA_8878_out0;
wire v$CINA_8879_out0;
wire v$CINA_8880_out0;
wire v$CINA_8881_out0;
wire v$CINA_8882_out0;
wire v$CINA_8883_out0;
wire v$CINA_8884_out0;
wire v$CINA_8885_out0;
wire v$CINA_8886_out0;
wire v$CINA_8887_out0;
wire v$CINA_8888_out0;
wire v$CINA_8889_out0;
wire v$CINA_8890_out0;
wire v$CINA_8891_out0;
wire v$CINA_8892_out0;
wire v$CINA_8893_out0;
wire v$CINA_8894_out0;
wire v$CINA_8895_out0;
wire v$CINA_8896_out0;
wire v$CINA_8897_out0;
wire v$CINA_8898_out0;
wire v$CINA_8899_out0;
wire v$CINA_8900_out0;
wire v$CINA_8901_out0;
wire v$CINA_8902_out0;
wire v$CINA_8903_out0;
wire v$CINA_8904_out0;
wire v$CINA_8905_out0;
wire v$CINA_8906_out0;
wire v$CINA_8907_out0;
wire v$CINA_8908_out0;
wire v$CINA_8909_out0;
wire v$CINA_8910_out0;
wire v$CINA_8911_out0;
wire v$CINA_8912_out0;
wire v$CINA_8913_out0;
wire v$CINA_8914_out0;
wire v$CINA_8915_out0;
wire v$CINA_8916_out0;
wire v$CINA_8917_out0;
wire v$CINA_8918_out0;
wire v$CINA_8919_out0;
wire v$CINA_8920_out0;
wire v$CINA_8921_out0;
wire v$CINA_8922_out0;
wire v$CINA_8923_out0;
wire v$CINA_8924_out0;
wire v$CINA_8925_out0;
wire v$CINA_8926_out0;
wire v$CINA_8927_out0;
wire v$CINA_8928_out0;
wire v$CINA_8929_out0;
wire v$CINA_8930_out0;
wire v$CINA_8931_out0;
wire v$CINA_8932_out0;
wire v$CINA_8933_out0;
wire v$CINA_8934_out0;
wire v$CINA_8935_out0;
wire v$CINA_8936_out0;
wire v$CINA_8937_out0;
wire v$CINA_8938_out0;
wire v$CINA_8939_out0;
wire v$CINA_8940_out0;
wire v$CINA_8941_out0;
wire v$CINA_8942_out0;
wire v$CINA_8943_out0;
wire v$CINA_8944_out0;
wire v$CINA_8945_out0;
wire v$CINA_8946_out0;
wire v$CINA_8947_out0;
wire v$CINA_8948_out0;
wire v$CINA_8949_out0;
wire v$CINA_8950_out0;
wire v$CINA_8951_out0;
wire v$CINA_8952_out0;
wire v$CINA_8953_out0;
wire v$CINA_8954_out0;
wire v$CINA_8955_out0;
wire v$CINA_8956_out0;
wire v$CINA_8957_out0;
wire v$CINA_8958_out0;
wire v$CINA_8959_out0;
wire v$CINA_8960_out0;
wire v$CINA_8961_out0;
wire v$CINA_8962_out0;
wire v$CINA_8963_out0;
wire v$CINA_8964_out0;
wire v$CINA_8965_out0;
wire v$CINA_8966_out0;
wire v$CINA_8967_out0;
wire v$CINA_8968_out0;
wire v$CINA_8969_out0;
wire v$CINA_8970_out0;
wire v$CINA_8971_out0;
wire v$CINA_8972_out0;
wire v$CINA_8973_out0;
wire v$CINA_8974_out0;
wire v$CINA_8975_out0;
wire v$CINA_8976_out0;
wire v$CINA_8977_out0;
wire v$CINA_8978_out0;
wire v$CINA_8979_out0;
wire v$CINA_8980_out0;
wire v$CINA_8981_out0;
wire v$CINA_8982_out0;
wire v$CINA_8983_out0;
wire v$CINA_8984_out0;
wire v$CINA_8985_out0;
wire v$CINA_8986_out0;
wire v$CINA_8987_out0;
wire v$CINA_8988_out0;
wire v$CINA_8989_out0;
wire v$CINA_8990_out0;
wire v$CINA_8991_out0;
wire v$CINA_8992_out0;
wire v$CINA_8993_out0;
wire v$CINA_8994_out0;
wire v$CINA_8995_out0;
wire v$CINA_8996_out0;
wire v$CINA_8997_out0;
wire v$CINA_8998_out0;
wire v$CINA_8999_out0;
wire v$CINA_9000_out0;
wire v$CINA_9001_out0;
wire v$CINA_9002_out0;
wire v$CINA_9003_out0;
wire v$CINA_9004_out0;
wire v$CINA_9005_out0;
wire v$CINA_9006_out0;
wire v$CINA_9007_out0;
wire v$CINA_9008_out0;
wire v$CINA_9009_out0;
wire v$CINA_9010_out0;
wire v$CINA_9011_out0;
wire v$CINA_9012_out0;
wire v$CINA_9013_out0;
wire v$CINA_9014_out0;
wire v$CINA_9015_out0;
wire v$CIN_15669_out0;
wire v$CIN_15670_out0;
wire v$CIN_15671_out0;
wire v$CIN_15672_out0;
wire v$CIN_15673_out0;
wire v$CIN_15674_out0;
wire v$CIN_16717_out0;
wire v$CIN_16718_out0;
wire v$CIN_16719_out0;
wire v$CIN_16720_out0;
wire v$CIN_16721_out0;
wire v$CIN_16722_out0;
wire v$CIN_17983_out0;
wire v$CIN_17984_out0;
wire v$CIN_17985_out0;
wire v$CIN_17986_out0;
wire v$CIN_17987_out0;
wire v$CIN_17988_out0;
wire v$CIN_18826_out0;
wire v$CIN_18827_out0;
wire v$CIN_18828_out0;
wire v$CIN_18829_out0;
wire v$CIN_18830_out0;
wire v$CIN_18831_out0;
wire v$CIN_18832_out0;
wire v$CIN_18833_out0;
wire v$CLEAR_19011_out0;
wire v$CLEAR_19012_out0;
wire v$CLK4_12779_out0;
wire v$CLK4_12780_out0;
wire v$CLK4_17354_out0;
wire v$CLK4_17355_out0;
wire v$CLK4_18601_out0;
wire v$CLK4_18602_out0;
wire v$CLK4_2728_out0;
wire v$CLK4_2729_out0;
wire v$CLK4_3873_out0;
wire v$CLK4_3874_out0;
wire v$CLK4_7347_out0;
wire v$CLK4_7348_out0;
wire v$CLK4_9180_out0;
wire v$CLK4_9181_out0;
wire v$CLRINTERRUPTS_356_out0;
wire v$CLRINTERRUPTS_357_out0;
wire v$CLR_4601_out0;
wire v$CLR_4602_out0;
wire v$COMP$H$OUT_6881_out0;
wire v$COMP$H$OUT_6882_out0;
wire v$COMP$L$OUT_12263_out0;
wire v$COMP$L$OUT_12264_out0;
wire v$CON1_4236_out0;
wire v$CON1_4237_out0;
wire v$CON1_4238_out0;
wire v$CON1_4239_out0;
wire v$CON1_4240_out0;
wire v$CON1_4241_out0;
wire v$CON2_14971_out0;
wire v$CON2_14972_out0;
wire v$CON2_14973_out0;
wire v$CON2_14974_out0;
wire v$CON2_14975_out0;
wire v$CON2_14976_out0;
wire v$CON3_8239_out0;
wire v$CON3_8240_out0;
wire v$CON3_8241_out0;
wire v$CON3_8242_out0;
wire v$CON3_8243_out0;
wire v$CON3_8244_out0;
wire v$CON4_17057_out0;
wire v$CON4_17058_out0;
wire v$CON4_17059_out0;
wire v$CON4_17060_out0;
wire v$CON4_17061_out0;
wire v$CON4_17062_out0;
wire v$CON5_11176_out0;
wire v$CON5_11177_out0;
wire v$CON5_11178_out0;
wire v$CON5_11179_out0;
wire v$CON5_11180_out0;
wire v$CON5_11181_out0;
wire v$CON6_13571_out0;
wire v$CON6_13572_out0;
wire v$CON6_13573_out0;
wire v$CON6_13574_out0;
wire v$CON6_13575_out0;
wire v$CON6_13576_out0;
wire v$CON7_2614_out0;
wire v$CON7_2615_out0;
wire v$CON7_2616_out0;
wire v$CON7_2617_out0;
wire v$CON7_2618_out0;
wire v$CON7_2619_out0;
wire v$COUNTEREN_14035_out0;
wire v$COUNTEREN_14036_out0;
wire v$COUNTEREN_1782_out0;
wire v$COUNTEREN_1783_out0;
wire v$COUNTERINTERRUPT_15460_out0;
wire v$COUNTERINTERRUPT_15461_out0;
wire v$COUTD_6930_out0;
wire v$COUTD_6931_out0;
wire v$COUTD_6932_out0;
wire v$COUTD_6933_out0;
wire v$COUTD_6934_out0;
wire v$COUTD_6935_out0;
wire v$COUTD_6936_out0;
wire v$COUTD_6937_out0;
wire v$COUTD_6938_out0;
wire v$COUTD_6939_out0;
wire v$COUTD_6940_out0;
wire v$COUTD_6941_out0;
wire v$COUTD_6942_out0;
wire v$COUTD_6943_out0;
wire v$COUTD_6944_out0;
wire v$COUTD_6945_out0;
wire v$COUTD_6946_out0;
wire v$COUTD_6947_out0;
wire v$COUTD_6948_out0;
wire v$COUTD_6949_out0;
wire v$COUTD_6950_out0;
wire v$COUTD_6951_out0;
wire v$COUTD_6952_out0;
wire v$COUTD_6953_out0;
wire v$COUTD_6954_out0;
wire v$COUTD_6955_out0;
wire v$COUTD_6956_out0;
wire v$COUTD_6957_out0;
wire v$COUTD_6958_out0;
wire v$COUTD_6959_out0;
wire v$COUTD_6960_out0;
wire v$COUTD_6961_out0;
wire v$COUTD_6962_out0;
wire v$COUTD_6963_out0;
wire v$COUTD_6964_out0;
wire v$COUTD_6965_out0;
wire v$COUTD_6966_out0;
wire v$COUTD_6967_out0;
wire v$COUTD_6968_out0;
wire v$COUTD_6969_out0;
wire v$COUTD_6970_out0;
wire v$COUTD_6971_out0;
wire v$COUTD_6972_out0;
wire v$COUTD_6973_out0;
wire v$COUTD_6974_out0;
wire v$COUTD_6975_out0;
wire v$COUTD_6976_out0;
wire v$COUTD_6977_out0;
wire v$COUTD_6978_out0;
wire v$COUTD_6979_out0;
wire v$COUTD_6980_out0;
wire v$COUTD_6981_out0;
wire v$COUTD_6982_out0;
wire v$COUTD_6983_out0;
wire v$COUTD_6984_out0;
wire v$COUTD_6985_out0;
wire v$COUTD_6986_out0;
wire v$COUTD_6987_out0;
wire v$COUTD_6988_out0;
wire v$COUTD_6989_out0;
wire v$COUTD_6990_out0;
wire v$COUTD_6991_out0;
wire v$COUTD_6992_out0;
wire v$COUTD_6993_out0;
wire v$COUTD_6994_out0;
wire v$COUTD_6995_out0;
wire v$COUTD_6996_out0;
wire v$COUTD_6997_out0;
wire v$COUTD_6998_out0;
wire v$COUTD_6999_out0;
wire v$COUTD_7000_out0;
wire v$COUTD_7001_out0;
wire v$COUTD_7002_out0;
wire v$COUTD_7003_out0;
wire v$COUTD_7004_out0;
wire v$COUTD_7005_out0;
wire v$COUTD_7006_out0;
wire v$COUTD_7007_out0;
wire v$COUTD_7008_out0;
wire v$COUTD_7009_out0;
wire v$COUTD_7010_out0;
wire v$COUTD_7011_out0;
wire v$COUTD_7012_out0;
wire v$COUTD_7013_out0;
wire v$COUTD_7014_out0;
wire v$COUTD_7015_out0;
wire v$COUTD_7016_out0;
wire v$COUTD_7017_out0;
wire v$COUTD_7018_out0;
wire v$COUTD_7019_out0;
wire v$COUTD_7020_out0;
wire v$COUTD_7021_out0;
wire v$COUTD_7022_out0;
wire v$COUTD_7023_out0;
wire v$COUTD_7024_out0;
wire v$COUTD_7025_out0;
wire v$COUTD_7026_out0;
wire v$COUTD_7027_out0;
wire v$COUTD_7028_out0;
wire v$COUTD_7029_out0;
wire v$COUTD_7030_out0;
wire v$COUTD_7031_out0;
wire v$COUTD_7032_out0;
wire v$COUTD_7033_out0;
wire v$COUTD_7034_out0;
wire v$COUTD_7035_out0;
wire v$COUTD_7036_out0;
wire v$COUTD_7037_out0;
wire v$COUTD_7038_out0;
wire v$COUTD_7039_out0;
wire v$COUTD_7040_out0;
wire v$COUTD_7041_out0;
wire v$COUTD_7042_out0;
wire v$COUTD_7043_out0;
wire v$COUTD_7044_out0;
wire v$COUTD_7045_out0;
wire v$COUTD_7046_out0;
wire v$COUTD_7047_out0;
wire v$COUTD_7048_out0;
wire v$COUTD_7049_out0;
wire v$COUTD_7050_out0;
wire v$COUTD_7051_out0;
wire v$COUTD_7052_out0;
wire v$COUTD_7053_out0;
wire v$COUTD_7054_out0;
wire v$COUTD_7055_out0;
wire v$COUTD_7056_out0;
wire v$COUTD_7057_out0;
wire v$COUTD_7058_out0;
wire v$COUTD_7059_out0;
wire v$COUTD_7060_out0;
wire v$COUTD_7061_out0;
wire v$COUTD_7062_out0;
wire v$COUTD_7063_out0;
wire v$COUTD_7064_out0;
wire v$COUTD_7065_out0;
wire v$COUTD_7066_out0;
wire v$COUTD_7067_out0;
wire v$COUTD_7068_out0;
wire v$COUTD_7069_out0;
wire v$COUTD_7070_out0;
wire v$COUTD_7071_out0;
wire v$COUTD_7072_out0;
wire v$COUTD_7073_out0;
wire v$COUTD_7074_out0;
wire v$COUTD_7075_out0;
wire v$COUTD_7076_out0;
wire v$COUTD_7077_out0;
wire v$COUTD_7078_out0;
wire v$COUTD_7079_out0;
wire v$COUTD_7080_out0;
wire v$COUTD_7081_out0;
wire v$COUTD_7082_out0;
wire v$COUTD_7083_out0;
wire v$COUTD_7084_out0;
wire v$COUTD_7085_out0;
wire v$COUTD_7086_out0;
wire v$COUTD_7087_out0;
wire v$COUTD_7088_out0;
wire v$COUTD_7089_out0;
wire v$COUTD_7090_out0;
wire v$COUTD_7091_out0;
wire v$COUTD_7092_out0;
wire v$COUTD_7093_out0;
wire v$COUTD_7094_out0;
wire v$COUTD_7095_out0;
wire v$COUTD_7096_out0;
wire v$COUTD_7097_out0;
wire v$COUTD_7098_out0;
wire v$COUTD_7099_out0;
wire v$COUTD_7100_out0;
wire v$COUTD_7101_out0;
wire v$COUTD_7102_out0;
wire v$COUTD_7103_out0;
wire v$COUTD_7104_out0;
wire v$COUTD_7105_out0;
wire v$COUTD_7106_out0;
wire v$COUTD_7107_out0;
wire v$COUTD_7108_out0;
wire v$COUTD_7109_out0;
wire v$COUTD_7110_out0;
wire v$COUTD_7111_out0;
wire v$COUTD_7112_out0;
wire v$COUTD_7113_out0;
wire v$COUTD_7114_out0;
wire v$COUTD_7115_out0;
wire v$COUTD_7116_out0;
wire v$COUTD_7117_out0;
wire v$COUTD_7118_out0;
wire v$COUTD_7119_out0;
wire v$COUTD_7120_out0;
wire v$COUTD_7121_out0;
wire v$COUTD_7122_out0;
wire v$COUTD_7123_out0;
wire v$COUTD_7124_out0;
wire v$COUTD_7125_out0;
wire v$COUTD_7126_out0;
wire v$COUTD_7127_out0;
wire v$COUTD_7128_out0;
wire v$COUTD_7129_out0;
wire v$COUTD_7130_out0;
wire v$COUTD_7131_out0;
wire v$COUTD_7132_out0;
wire v$COUTD_7133_out0;
wire v$COUTD_7134_out0;
wire v$COUTD_7135_out0;
wire v$COUTD_7136_out0;
wire v$COUTD_7137_out0;
wire v$COUTD_7138_out0;
wire v$COUTD_7139_out0;
wire v$COUTD_7140_out0;
wire v$COUTD_7141_out0;
wire v$COUTD_7142_out0;
wire v$COUTD_7143_out0;
wire v$COUTD_7144_out0;
wire v$COUTD_7145_out0;
wire v$COUTD_7146_out0;
wire v$COUTD_7147_out0;
wire v$COUTD_7148_out0;
wire v$COUTD_7149_out0;
wire v$COUTD_7150_out0;
wire v$COUTD_7151_out0;
wire v$COUTD_7152_out0;
wire v$COUTD_7153_out0;
wire v$COUTD_7154_out0;
wire v$COUTD_7155_out0;
wire v$COUTD_7156_out0;
wire v$COUTD_7157_out0;
wire v$COUTD_7158_out0;
wire v$COUTD_7159_out0;
wire v$COUTD_7160_out0;
wire v$COUTD_7161_out0;
wire v$COUTD_7162_out0;
wire v$COUTD_7163_out0;
wire v$COUTD_7164_out0;
wire v$COUTD_7165_out0;
wire v$COUTD_7166_out0;
wire v$COUTD_7167_out0;
wire v$COUTD_7168_out0;
wire v$COUTD_7169_out0;
wire v$COUTD_7170_out0;
wire v$COUTD_7171_out0;
wire v$COUTD_7172_out0;
wire v$COUTD_7173_out0;
wire v$COUTD_7174_out0;
wire v$COUTD_7175_out0;
wire v$COUT_14088_out0;
wire v$COUT_14089_out0;
wire v$COUT_8603_out0;
wire v$COUT_8604_out0;
wire v$C_16498_out0;
wire v$C_16499_out0;
wire v$C_3419_out0;
wire v$C_3420_out0;
wire v$C_3832_out0;
wire v$C_3833_out0;
wire v$C_6338_out0;
wire v$C_6339_out0;
wire v$C_9990_out0;
wire v$C_9991_out0;
wire v$CheckParity_19290_out0;
wire v$CheckParity_19291_out0;
wire v$Clear_13319_out0;
wire v$Clear_13320_out0;
wire v$Clear_15245_out0;
wire v$Clear_15246_out0;
wire v$D1_14709_out0;
wire v$D1_14709_out1;
wire v$D1_14709_out2;
wire v$D1_14709_out3;
wire v$D1_14710_out0;
wire v$D1_14710_out1;
wire v$D1_14710_out2;
wire v$D1_14710_out3;
wire v$DATA$DEPENDENCY_6422_out0;
wire v$DATA$DEPENDENCY_6423_out0;
wire v$DATA$PROCESS$WB_18439_out0;
wire v$DATA$PROCESS$WB_18440_out0;
wire v$DISABLEINTERRUPTS_15588_out0;
wire v$DISABLEINTERRUPTS_15589_out0;
wire v$DM1_16855_out0;
wire v$DM1_16855_out1;
wire v$EDGE0_4146_out0;
wire v$EDGE0_4147_out0;
wire v$EDGE0_6025_out0;
wire v$EDGE0_6026_out0;
wire v$EDGE1_15855_out0;
wire v$EDGE1_15856_out0;
wire v$EDGE1_18050_out0;
wire v$EDGE1_18051_out0;
wire v$EDGE2_18729_out0;
wire v$EDGE2_18730_out0;
wire v$EDGE2_7280_out0;
wire v$EDGE2_7281_out0;
wire v$EDGE3_11552_out0;
wire v$EDGE3_11553_out0;
wire v$EDGE3_2446_out0;
wire v$EDGE3_2447_out0;
wire v$ENABLEINTERRUPTS_13141_out0;
wire v$ENABLEINTERRUPTS_13142_out0;
wire v$ENABLEINTERRUPTS_17620_out0;
wire v$ENABLEINTERRUPTS_17621_out0;
wire v$ENCODED0_14632_out0;
wire v$ENCODED0_14633_out0;
wire v$ENCODED1_9898_out0;
wire v$ENCODED1_9899_out0;
wire v$END0_9721_out0;
wire v$END0_9722_out0;
wire v$END0_9723_out0;
wire v$END0_9724_out0;
wire v$END0_9725_out0;
wire v$END0_9726_out0;
wire v$END10_1295_out0;
wire v$END10_1296_out0;
wire v$END10_1297_out0;
wire v$END10_1298_out0;
wire v$END10_1299_out0;
wire v$END10_1300_out0;
wire v$END11_12655_out0;
wire v$END11_12656_out0;
wire v$END11_12657_out0;
wire v$END11_12658_out0;
wire v$END11_12659_out0;
wire v$END11_12660_out0;
wire v$END12_11274_out0;
wire v$END12_11275_out0;
wire v$END12_11276_out0;
wire v$END12_11277_out0;
wire v$END12_11278_out0;
wire v$END12_11279_out0;
wire v$END13_18673_out0;
wire v$END13_18674_out0;
wire v$END13_18675_out0;
wire v$END13_18676_out0;
wire v$END13_18677_out0;
wire v$END13_18678_out0;
wire v$END14_284_out0;
wire v$END14_285_out0;
wire v$END14_286_out0;
wire v$END14_287_out0;
wire v$END14_288_out0;
wire v$END14_289_out0;
wire v$END15_7696_out0;
wire v$END15_7697_out0;
wire v$END15_7698_out0;
wire v$END15_7699_out0;
wire v$END15_7700_out0;
wire v$END15_7701_out0;
wire v$END16_222_out0;
wire v$END16_223_out0;
wire v$END16_224_out0;
wire v$END16_225_out0;
wire v$END16_226_out0;
wire v$END16_227_out0;
wire v$END17_7965_out0;
wire v$END17_7966_out0;
wire v$END17_7967_out0;
wire v$END17_7968_out0;
wire v$END17_7969_out0;
wire v$END17_7970_out0;
wire v$END18_12519_out0;
wire v$END18_12520_out0;
wire v$END18_12521_out0;
wire v$END18_12522_out0;
wire v$END18_12523_out0;
wire v$END18_12524_out0;
wire v$END19_12218_out0;
wire v$END19_12219_out0;
wire v$END19_12220_out0;
wire v$END19_12221_out0;
wire v$END19_12222_out0;
wire v$END19_12223_out0;
wire v$END1_1450_out0;
wire v$END1_1451_out0;
wire v$END1_1452_out0;
wire v$END1_1453_out0;
wire v$END1_1454_out0;
wire v$END1_1455_out0;
wire v$END1_1697_out0;
wire v$END1_1698_out0;
wire v$END1_1699_out0;
wire v$END1_1700_out0;
wire v$END1_1701_out0;
wire v$END1_1702_out0;
wire v$END1_7241_out0;
wire v$END1_7242_out0;
wire v$END1_7268_out0;
wire v$END1_7269_out0;
wire v$END20_13847_out0;
wire v$END20_13848_out0;
wire v$END20_13849_out0;
wire v$END20_13850_out0;
wire v$END20_13851_out0;
wire v$END20_13852_out0;
wire v$END21_4504_out0;
wire v$END21_4505_out0;
wire v$END21_4506_out0;
wire v$END21_4507_out0;
wire v$END21_4508_out0;
wire v$END21_4509_out0;
wire v$END22_16073_out0;
wire v$END22_16074_out0;
wire v$END22_16075_out0;
wire v$END22_16076_out0;
wire v$END22_16077_out0;
wire v$END22_16078_out0;
wire v$END23_17336_out0;
wire v$END23_17337_out0;
wire v$END23_17338_out0;
wire v$END23_17339_out0;
wire v$END23_17340_out0;
wire v$END23_17341_out0;
wire v$END24_17022_out0;
wire v$END24_17023_out0;
wire v$END24_17024_out0;
wire v$END24_17025_out0;
wire v$END24_17026_out0;
wire v$END24_17027_out0;
wire v$END25_17666_out0;
wire v$END25_17667_out0;
wire v$END25_17668_out0;
wire v$END25_17669_out0;
wire v$END25_17670_out0;
wire v$END25_17671_out0;
wire v$END26_6678_out0;
wire v$END26_6679_out0;
wire v$END26_6680_out0;
wire v$END26_6681_out0;
wire v$END26_6682_out0;
wire v$END26_6683_out0;
wire v$END27_2414_out0;
wire v$END27_2415_out0;
wire v$END27_2416_out0;
wire v$END27_2417_out0;
wire v$END27_2418_out0;
wire v$END27_2419_out0;
wire v$END28_14248_out0;
wire v$END28_14249_out0;
wire v$END28_14250_out0;
wire v$END28_14251_out0;
wire v$END28_14252_out0;
wire v$END28_14253_out0;
wire v$END29_6161_out0;
wire v$END29_6162_out0;
wire v$END29_6163_out0;
wire v$END29_6164_out0;
wire v$END29_6165_out0;
wire v$END29_6166_out0;
wire v$END2_5449_out0;
wire v$END2_5450_out0;
wire v$END2_5451_out0;
wire v$END2_5452_out0;
wire v$END2_5453_out0;
wire v$END2_5454_out0;
wire v$END2_8068_out0;
wire v$END2_8069_out0;
wire v$END2_8070_out0;
wire v$END2_8071_out0;
wire v$END2_8072_out0;
wire v$END2_8073_out0;
wire v$END30_16309_out0;
wire v$END30_16310_out0;
wire v$END30_16311_out0;
wire v$END30_16312_out0;
wire v$END30_16313_out0;
wire v$END30_16314_out0;
wire v$END31_19131_out0;
wire v$END31_19132_out0;
wire v$END31_19133_out0;
wire v$END31_19134_out0;
wire v$END31_19135_out0;
wire v$END31_19136_out0;
wire v$END32_2664_out0;
wire v$END32_2665_out0;
wire v$END32_2666_out0;
wire v$END32_2667_out0;
wire v$END32_2668_out0;
wire v$END32_2669_out0;
wire v$END33_273_out0;
wire v$END33_274_out0;
wire v$END33_275_out0;
wire v$END33_276_out0;
wire v$END33_277_out0;
wire v$END33_278_out0;
wire v$END3_3655_out0;
wire v$END3_3656_out0;
wire v$END3_3657_out0;
wire v$END3_3658_out0;
wire v$END3_3659_out0;
wire v$END3_3660_out0;
wire v$END3_8257_out0;
wire v$END3_8258_out0;
wire v$END3_8259_out0;
wire v$END3_8260_out0;
wire v$END3_8261_out0;
wire v$END3_8262_out0;
wire v$END40_6062_out0;
wire v$END40_6063_out0;
wire v$END40_6064_out0;
wire v$END40_6065_out0;
wire v$END40_6066_out0;
wire v$END40_6067_out0;
wire v$END41_17286_out0;
wire v$END41_17287_out0;
wire v$END41_17288_out0;
wire v$END41_17289_out0;
wire v$END41_17290_out0;
wire v$END41_17291_out0;
wire v$END42_18916_out0;
wire v$END42_18917_out0;
wire v$END42_18918_out0;
wire v$END42_18919_out0;
wire v$END42_18920_out0;
wire v$END42_18921_out0;
wire v$END43_13771_out0;
wire v$END43_13772_out0;
wire v$END43_13773_out0;
wire v$END43_13774_out0;
wire v$END43_13775_out0;
wire v$END43_13776_out0;
wire v$END44_16258_out0;
wire v$END44_16259_out0;
wire v$END44_16260_out0;
wire v$END44_16261_out0;
wire v$END44_16262_out0;
wire v$END44_16263_out0;
wire v$END45_9383_out0;
wire v$END45_9384_out0;
wire v$END45_9385_out0;
wire v$END45_9386_out0;
wire v$END45_9387_out0;
wire v$END45_9388_out0;
wire v$END46_15663_out0;
wire v$END46_15664_out0;
wire v$END46_15665_out0;
wire v$END46_15666_out0;
wire v$END46_15667_out0;
wire v$END46_15668_out0;
wire v$END47_2876_out0;
wire v$END47_2877_out0;
wire v$END47_2878_out0;
wire v$END47_2879_out0;
wire v$END47_2880_out0;
wire v$END47_2881_out0;
wire v$END48_10827_out0;
wire v$END48_10828_out0;
wire v$END48_10829_out0;
wire v$END48_10830_out0;
wire v$END48_10831_out0;
wire v$END48_10832_out0;
wire v$END49_19059_out0;
wire v$END49_19060_out0;
wire v$END49_19061_out0;
wire v$END49_19062_out0;
wire v$END49_19063_out0;
wire v$END49_19064_out0;
wire v$END4_3491_out0;
wire v$END4_3492_out0;
wire v$END4_5463_out0;
wire v$END4_5464_out0;
wire v$END4_5465_out0;
wire v$END4_5466_out0;
wire v$END4_5467_out0;
wire v$END4_5468_out0;
wire v$END4_8432_out0;
wire v$END4_8433_out0;
wire v$END4_9737_out0;
wire v$END4_9738_out0;
wire v$END4_9739_out0;
wire v$END4_9740_out0;
wire v$END4_9741_out0;
wire v$END4_9742_out0;
wire v$END50_7729_out0;
wire v$END50_7730_out0;
wire v$END50_7731_out0;
wire v$END50_7732_out0;
wire v$END50_7733_out0;
wire v$END50_7734_out0;
wire v$END51_12242_out0;
wire v$END51_12243_out0;
wire v$END51_12244_out0;
wire v$END51_12245_out0;
wire v$END51_12246_out0;
wire v$END51_12247_out0;
wire v$END52_12549_out0;
wire v$END52_12550_out0;
wire v$END52_12551_out0;
wire v$END52_12552_out0;
wire v$END52_12553_out0;
wire v$END52_12554_out0;
wire v$END53_330_out0;
wire v$END53_331_out0;
wire v$END53_332_out0;
wire v$END53_333_out0;
wire v$END53_334_out0;
wire v$END53_335_out0;
wire v$END5_4301_out0;
wire v$END5_4302_out0;
wire v$END5_4303_out0;
wire v$END5_4304_out0;
wire v$END5_4305_out0;
wire v$END5_4306_out0;
wire v$END60_15741_out0;
wire v$END60_15742_out0;
wire v$END60_15743_out0;
wire v$END60_15744_out0;
wire v$END60_15745_out0;
wire v$END60_15746_out0;
wire v$END61_18570_out0;
wire v$END61_18571_out0;
wire v$END61_18572_out0;
wire v$END61_18573_out0;
wire v$END61_18574_out0;
wire v$END61_18575_out0;
wire v$END6_15831_out0;
wire v$END6_15832_out0;
wire v$END6_15833_out0;
wire v$END6_15834_out0;
wire v$END6_15835_out0;
wire v$END6_15836_out0;
wire v$END6_7866_out0;
wire v$END6_7867_out0;
wire v$END7_3582_out0;
wire v$END7_3583_out0;
wire v$END7_3584_out0;
wire v$END7_3585_out0;
wire v$END7_3586_out0;
wire v$END7_3587_out0;
wire v$END8_4070_out0;
wire v$END8_4071_out0;
wire v$END8_4072_out0;
wire v$END8_4073_out0;
wire v$END8_4074_out0;
wire v$END8_4075_out0;
wire v$END9_4392_out0;
wire v$END9_4393_out0;
wire v$END9_4394_out0;
wire v$END9_4395_out0;
wire v$END9_4396_out0;
wire v$END9_4397_out0;
wire v$END_16336_out0;
wire v$END_16337_out0;
wire v$END_17644_out0;
wire v$END_17645_out0;
wire v$END_18875_out0;
wire v$END_18876_out0;
wire v$END_18877_out0;
wire v$END_18878_out0;
wire v$END_18879_out0;
wire v$END_18880_out0;
wire v$END_3541_out0;
wire v$END_3542_out0;
wire v$END_3543_out0;
wire v$END_3544_out0;
wire v$END_3545_out0;
wire v$END_3546_out0;
wire v$END_8410_out0;
wire v$END_8411_out0;
wire v$ENDa_17183_out0;
wire v$ENDa_17184_out0;
wire v$ENDa_17185_out0;
wire v$ENDa_17186_out0;
wire v$ENDa_17187_out0;
wire v$ENDa_17188_out0;
wire v$ENDd_11330_out0;
wire v$ENDd_11331_out0;
wire v$ENDd_11332_out0;
wire v$ENDd_11333_out0;
wire v$ENDd_11334_out0;
wire v$ENDd_11335_out0;
wire v$ENDe_18504_out0;
wire v$ENDe_18505_out0;
wire v$ENDe_18506_out0;
wire v$ENDe_18507_out0;
wire v$ENDe_18508_out0;
wire v$ENDe_18509_out0;
wire v$ENDi_9030_out0;
wire v$ENDi_9031_out0;
wire v$ENDi_9032_out0;
wire v$ENDi_9033_out0;
wire v$ENDi_9034_out0;
wire v$ENDi_9035_out0;
wire v$ENDo_19304_out0;
wire v$ENDo_19305_out0;
wire v$ENDo_19306_out0;
wire v$ENDo_19307_out0;
wire v$ENDo_19308_out0;
wire v$ENDo_19309_out0;
wire v$ENDp_3409_out0;
wire v$ENDp_3410_out0;
wire v$ENDp_3411_out0;
wire v$ENDp_3412_out0;
wire v$ENDp_3413_out0;
wire v$ENDp_3414_out0;
wire v$ENDq_1609_out0;
wire v$ENDq_1610_out0;
wire v$ENDq_1611_out0;
wire v$ENDq_1612_out0;
wire v$ENDq_1613_out0;
wire v$ENDq_1614_out0;
wire v$ENDr_7842_out0;
wire v$ENDr_7843_out0;
wire v$ENDr_7844_out0;
wire v$ENDr_7845_out0;
wire v$ENDr_7846_out0;
wire v$ENDr_7847_out0;
wire v$ENDs_3435_out0;
wire v$ENDs_3436_out0;
wire v$ENDs_3437_out0;
wire v$ENDs_3438_out0;
wire v$ENDs_3439_out0;
wire v$ENDs_3440_out0;
wire v$ENDt_10711_out0;
wire v$ENDt_10712_out0;
wire v$ENDt_10713_out0;
wire v$ENDt_10714_out0;
wire v$ENDt_10715_out0;
wire v$ENDt_10716_out0;
wire v$ENDu_7313_out0;
wire v$ENDu_7314_out0;
wire v$ENDu_7315_out0;
wire v$ENDu_7316_out0;
wire v$ENDu_7317_out0;
wire v$ENDu_7318_out0;
wire v$ENDw_9930_out0;
wire v$ENDw_9931_out0;
wire v$ENDw_9932_out0;
wire v$ENDw_9933_out0;
wire v$ENDw_9934_out0;
wire v$ENDw_9935_out0;
wire v$ENDy_4271_out0;
wire v$ENDy_4272_out0;
wire v$ENDy_4273_out0;
wire v$ENDy_4274_out0;
wire v$ENDy_4275_out0;
wire v$ENDy_4276_out0;
wire v$ENMODE_15175_out0;
wire v$ENMODE_15176_out0;
wire v$ENMODE_8055_out0;
wire v$ENMODE_8056_out0;
wire v$EN_1493_out0;
wire v$EN_1494_out0;
wire v$EN_1495_out0;
wire v$EN_1496_out0;
wire v$EN_1497_out0;
wire v$EN_1498_out0;
wire v$EN_1499_out0;
wire v$EN_1500_out0;
wire v$EN_1501_out0;
wire v$EN_1502_out0;
wire v$EN_1503_out0;
wire v$EN_1504_out0;
wire v$EN_1505_out0;
wire v$EN_1506_out0;
wire v$EN_1507_out0;
wire v$EN_1508_out0;
wire v$EN_1509_out0;
wire v$EN_1510_out0;
wire v$EN_1511_out0;
wire v$EN_1512_out0;
wire v$EN_16500_out0;
wire v$EN_16501_out0;
wire v$EN_17004_out0;
wire v$EN_17005_out0;
wire v$EN_17006_out0;
wire v$EN_17007_out0;
wire v$EN_17008_out0;
wire v$EN_17009_out0;
wire v$EN_17010_out0;
wire v$EN_17011_out0;
wire v$EN_17561_out0;
wire v$EN_17562_out0;
wire v$EN_17563_out0;
wire v$EN_17564_out0;
wire v$EN_17565_out0;
wire v$EN_17566_out0;
wire v$EN_17567_out0;
wire v$EN_17568_out0;
wire v$EN_4054_out0;
wire v$EN_4055_out0;
wire v$EN_4056_out0;
wire v$EN_4057_out0;
wire v$EN_4058_out0;
wire v$EN_4059_out0;
wire v$EN_4963_out0;
wire v$EN_4964_out0;
wire v$EN_4965_out0;
wire v$EN_4966_out0;
wire v$EN_4967_out0;
wire v$EN_4968_out0;
wire v$EN_4969_out0;
wire v$EN_4970_out0;
wire v$EN_4971_out0;
wire v$EN_4972_out0;
wire v$EN_4973_out0;
wire v$EN_4974_out0;
wire v$EN_5427_out0;
wire v$EN_5428_out0;
wire v$EN_5429_out0;
wire v$EN_5430_out0;
wire v$EN_5431_out0;
wire v$EN_5432_out0;
wire v$EN_5433_out0;
wire v$EN_5434_out0;
wire v$EN_5435_out0;
wire v$EN_5436_out0;
wire v$EN_5437_out0;
wire v$EN_5438_out0;
wire v$EN_8199_out0;
wire v$EN_8200_out0;
wire v$EN_8201_out0;
wire v$EN_8202_out0;
wire v$EN_8203_out0;
wire v$EN_8204_out0;
wire v$EN_8205_out0;
wire v$EN_8206_out0;
wire v$EN_8207_out0;
wire v$EN_8208_out0;
wire v$EN_8209_out0;
wire v$EN_8210_out0;
wire v$EN_9408_out0;
wire v$EN_9409_out0;
wire v$EPARITY_18914_out0;
wire v$EPARITY_18915_out0;
wire v$EQ$LDST_18074_out0;
wire v$EQ$LDST_18075_out0;
wire v$EQ10_10285_out0;
wire v$EQ10_10286_out0;
wire v$EQ10_13993_out0;
wire v$EQ10_13994_out0;
wire v$EQ10_6169_out0;
wire v$EQ10_6170_out0;
wire v$EQ10_6171_out0;
wire v$EQ10_6172_out0;
wire v$EQ11_12455_out0;
wire v$EQ11_12456_out0;
wire v$EQ11_14182_out0;
wire v$EQ11_14183_out0;
wire v$EQ11_6408_out0;
wire v$EQ11_6409_out0;
wire v$EQ11_6410_out0;
wire v$EQ11_6411_out0;
wire v$EQ12_13843_out0;
wire v$EQ12_13844_out0;
wire v$EQ12_14427_out0;
wire v$EQ12_14428_out0;
wire v$EQ12_14429_out0;
wire v$EQ12_14430_out0;
wire v$EQ12_15715_out0;
wire v$EQ12_15716_out0;
wire v$EQ12_1693_out0;
wire v$EQ12_1694_out0;
wire v$EQ13_19159_out0;
wire v$EQ13_19160_out0;
wire v$EQ13_5469_out0;
wire v$EQ13_5470_out0;
wire v$EQ13_9710_out0;
wire v$EQ13_9711_out0;
wire v$EQ13_9893_out0;
wire v$EQ13_9894_out0;
wire v$EQ13_9895_out0;
wire v$EQ13_9896_out0;
wire v$EQ14_12688_out0;
wire v$EQ14_12689_out0;
wire v$EQ14_5642_out0;
wire v$EQ14_5643_out0;
wire v$EQ14_5644_out0;
wire v$EQ14_5645_out0;
wire v$EQ14_5729_out0;
wire v$EQ14_5730_out0;
wire v$EQ15_16391_out0;
wire v$EQ15_16392_out0;
wire v$EQ15_16574_out0;
wire v$EQ15_16575_out0;
wire v$EQ15_16576_out0;
wire v$EQ15_16577_out0;
wire v$EQ15_17642_out0;
wire v$EQ15_17643_out0;
wire v$EQ16_11237_out0;
wire v$EQ16_11238_out0;
wire v$EQ16_1739_out0;
wire v$EQ16_1740_out0;
wire v$EQ16_8597_out0;
wire v$EQ16_8598_out0;
wire v$EQ16_8599_out0;
wire v$EQ16_8600_out0;
wire v$EQ17_6155_out0;
wire v$EQ17_6156_out0;
wire v$EQ17_6157_out0;
wire v$EQ17_6158_out0;
wire v$EQ18_13375_out0;
wire v$EQ18_13376_out0;
wire v$EQ18_13377_out0;
wire v$EQ18_13378_out0;
wire v$EQ19_5682_out0;
wire v$EQ19_5683_out0;
wire v$EQ19_5684_out0;
wire v$EQ19_5685_out0;
wire v$EQ1_10860_out0;
wire v$EQ1_10861_out0;
wire v$EQ1_12187_out0;
wire v$EQ1_12188_out0;
wire v$EQ1_13516_out0;
wire v$EQ1_13517_out0;
wire v$EQ1_13938_out0;
wire v$EQ1_13939_out0;
wire v$EQ1_13999_out0;
wire v$EQ1_14000_out0;
wire v$EQ1_14001_out0;
wire v$EQ1_14002_out0;
wire v$EQ1_14926_out0;
wire v$EQ1_14927_out0;
wire v$EQ1_15873_out0;
wire v$EQ1_15874_out0;
wire v$EQ1_15907_out0;
wire v$EQ1_15908_out0;
wire v$EQ1_16735_out0;
wire v$EQ1_16736_out0;
wire v$EQ1_16829_out0;
wire v$EQ1_16830_out0;
wire v$EQ1_16882_out0;
wire v$EQ1_16883_out0;
wire v$EQ1_18042_out0;
wire v$EQ1_18043_out0;
wire v$EQ1_19203_out0;
wire v$EQ1_19204_out0;
wire v$EQ1_2712_out0;
wire v$EQ1_2713_out0;
wire v$EQ1_3042_out0;
wire v$EQ1_3043_out0;
wire v$EQ1_3162_out0;
wire v$EQ1_3163_out0;
wire v$EQ1_3433_out0;
wire v$EQ1_3434_out0;
wire v$EQ1_4267_out0;
wire v$EQ1_4268_out0;
wire v$EQ1_5291_out0;
wire v$EQ1_5292_out0;
wire v$EQ1_5299_out0;
wire v$EQ1_5300_out0;
wire v$EQ1_7213_out0;
wire v$EQ1_7214_out0;
wire v$EQ1_7756_out0;
wire v$EQ1_7757_out0;
wire v$EQ1_8110_out0;
wire v$EQ1_8111_out0;
wire v$EQ20_10370_out0;
wire v$EQ20_10371_out0;
wire v$EQ20_10372_out0;
wire v$EQ20_10373_out0;
wire v$EQ21_3547_out0;
wire v$EQ21_3548_out0;
wire v$EQ21_3549_out0;
wire v$EQ21_3550_out0;
wire v$EQ22_3060_out0;
wire v$EQ22_3061_out0;
wire v$EQ22_3062_out0;
wire v$EQ22_3063_out0;
wire v$EQ23_3415_out0;
wire v$EQ23_3416_out0;
wire v$EQ23_3417_out0;
wire v$EQ23_3418_out0;
wire v$EQ24_2732_out0;
wire v$EQ24_2733_out0;
wire v$EQ24_2734_out0;
wire v$EQ24_2735_out0;
wire v$EQ2_11292_out0;
wire v$EQ2_11293_out0;
wire v$EQ2_12176_out0;
wire v$EQ2_12177_out0;
wire v$EQ2_13445_out0;
wire v$EQ2_13446_out0;
wire v$EQ2_14201_out0;
wire v$EQ2_14202_out0;
wire v$EQ2_14810_out0;
wire v$EQ2_14811_out0;
wire v$EQ2_14812_out0;
wire v$EQ2_14813_out0;
wire v$EQ2_14904_out0;
wire v$EQ2_14905_out0;
wire v$EQ2_16405_out0;
wire v$EQ2_16406_out0;
wire v$EQ2_16766_out0;
wire v$EQ2_16767_out0;
wire v$EQ2_17012_out0;
wire v$EQ2_17013_out0;
wire v$EQ2_17513_out0;
wire v$EQ2_17514_out0;
wire v$EQ2_19266_out0;
wire v$EQ2_19267_out0;
wire v$EQ2_3431_out0;
wire v$EQ2_3432_out0;
wire v$EQ2_4388_out0;
wire v$EQ2_4389_out0;
wire v$EQ2_8279_out0;
wire v$EQ2_8280_out0;
wire v$EQ3_12280_out0;
wire v$EQ3_12281_out0;
wire v$EQ3_12702_out0;
wire v$EQ3_12703_out0;
wire v$EQ3_14381_out0;
wire v$EQ3_14382_out0;
wire v$EQ3_14906_out0;
wire v$EQ3_14907_out0;
wire v$EQ3_15864_out0;
wire v$EQ3_15865_out0;
wire v$EQ3_16095_out0;
wire v$EQ3_16096_out0;
wire v$EQ3_17164_out0;
wire v$EQ3_17165_out0;
wire v$EQ3_18535_out0;
wire v$EQ3_18536_out0;
wire v$EQ3_1977_out0;
wire v$EQ3_1978_out0;
wire v$EQ3_1979_out0;
wire v$EQ3_1980_out0;
wire v$EQ3_2808_out0;
wire v$EQ3_2809_out0;
wire v$EQ3_4362_out0;
wire v$EQ3_4363_out0;
wire v$EQ3_5676_out0;
wire v$EQ3_5677_out0;
wire v$EQ3_6015_out0;
wire v$EQ3_6016_out0;
wire v$EQ3_7548_out0;
wire v$EQ3_7549_out0;
wire v$EQ3_8225_out0;
wire v$EQ3_8226_out0;
wire v$EQ4_10007_out0;
wire v$EQ4_10008_out0;
wire v$EQ4_13295_out0;
wire v$EQ4_13296_out0;
wire v$EQ4_17130_out0;
wire v$EQ4_17131_out0;
wire v$EQ4_17198_out0;
wire v$EQ4_17199_out0;
wire v$EQ4_17319_out0;
wire v$EQ4_17320_out0;
wire v$EQ4_19209_out0;
wire v$EQ4_19210_out0;
wire v$EQ4_19211_out0;
wire v$EQ4_19212_out0;
wire v$EQ4_2813_out0;
wire v$EQ4_2814_out0;
wire v$EQ4_3217_out0;
wire v$EQ4_3218_out0;
wire v$EQ4_5656_out0;
wire v$EQ4_5657_out0;
wire v$EQ4_9727_out0;
wire v$EQ4_9728_out0;
wire v$EQ5_10454_out0;
wire v$EQ5_10455_out0;
wire v$EQ5_14979_out0;
wire v$EQ5_14980_out0;
wire v$EQ5_1657_out0;
wire v$EQ5_1658_out0;
wire v$EQ5_2074_out0;
wire v$EQ5_2075_out0;
wire v$EQ5_3178_out0;
wire v$EQ5_3179_out0;
wire v$EQ5_3537_out0;
wire v$EQ5_3538_out0;
wire v$EQ5_3539_out0;
wire v$EQ5_3540_out0;
wire v$EQ5_3752_out0;
wire v$EQ5_3753_out0;
wire v$EQ5_5070_out0;
wire v$EQ5_5071_out0;
wire v$EQ5_9433_out0;
wire v$EQ5_9434_out0;
wire v$EQ6_16480_out0;
wire v$EQ6_16481_out0;
wire v$EQ6_16860_out0;
wire v$EQ6_16861_out0;
wire v$EQ6_1723_out0;
wire v$EQ6_1724_out0;
wire v$EQ6_4128_out0;
wire v$EQ6_4129_out0;
wire v$EQ6_5666_out0;
wire v$EQ6_5667_out0;
wire v$EQ6_5668_out0;
wire v$EQ6_5669_out0;
wire v$EQ6_6654_out0;
wire v$EQ6_6655_out0;
wire v$EQ7_14178_out0;
wire v$EQ7_14179_out0;
wire v$EQ7_17509_out0;
wire v$EQ7_17510_out0;
wire v$EQ7_19241_out0;
wire v$EQ7_19242_out0;
wire v$EQ7_239_out0;
wire v$EQ7_240_out0;
wire v$EQ7_3706_out0;
wire v$EQ7_3707_out0;
wire v$EQ7_4242_out0;
wire v$EQ7_4243_out0;
wire v$EQ7_4244_out0;
wire v$EQ7_4245_out0;
wire v$EQ8_14932_out0;
wire v$EQ8_14933_out0;
wire v$EQ8_15018_out0;
wire v$EQ8_15019_out0;
wire v$EQ8_15020_out0;
wire v$EQ8_15021_out0;
wire v$EQ8_16631_out0;
wire v$EQ8_16632_out0;
wire v$EQ8_261_out0;
wire v$EQ8_262_out0;
wire v$EQ9_14361_out0;
wire v$EQ9_14362_out0;
wire v$EQ9_14363_out0;
wire v$EQ9_14364_out0;
wire v$EQ9_18380_out0;
wire v$EQ9_18381_out0;
wire v$EQ9_18887_out0;
wire v$EQ9_18888_out0;
wire v$EQ9_8295_out0;
wire v$EQ9_8296_out0;
wire v$EQUAL_12184_out0;
wire v$EQUAL_12185_out0;
wire v$EQUAL_16432_out0;
wire v$EQUAL_16433_out0;
wire v$EQ_14007_out0;
wire v$EQ_14008_out0;
wire v$EQ_15177_out0;
wire v$EQ_15178_out0;
wire v$EQ_3677_out0;
wire v$EQ_3678_out0;
wire v$EQ_3889_out0;
wire v$EQ_3890_out0;
wire v$EQ_4490_out0;
wire v$EQ_4491_out0;
wire v$EQ_450_out0;
wire v$EQ_451_out0;
wire v$EQ_6416_out0;
wire v$EQ_6417_out0;
wire v$ERR_13343_out0;
wire v$ERR_13344_out0;
wire v$EVENPARITY_14162_out0;
wire v$EVENPARITY_14163_out0;
wire v$EXEC1$FPU_14256_out0;
wire v$EXEC1$FPU_14257_out0;
wire v$EXEC1_10709_out0;
wire v$EXEC1_10710_out0;
wire v$EXEC2_10281_out0;
wire v$EXEC2_10282_out0;
wire v$EXEC2_1313_out0;
wire v$EXEC2_1314_out0;
wire v$EXEC2_1621_out0;
wire v$EXEC2_1622_out0;
wire v$EXEC2_16486_out0;
wire v$EXEC2_16487_out0;
wire v$EXEC2_16981_out0;
wire v$EXEC2_16982_out0;
wire v$EXEC2_18249_out0;
wire v$EXEC2_18250_out0;
wire v$EXEC2_2109_out0;
wire v$EXEC2_2110_out0;
wire v$EXEC2_4154_out0;
wire v$EXEC2_4155_out0;
wire v$EXEC2_448_out0;
wire v$EXEC2_449_out0;
wire v$EXEC2_4552_out0;
wire v$EXEC2_4553_out0;
wire v$EXEC2_8333_out0;
wire v$EXEC2_8334_out0;
wire v$EXEC2_8362_out0;
wire v$EXEC2_8363_out0;
wire v$EXEC2_9813_out0;
wire v$EXEC2_9814_out0;
wire v$EXP$SAME_1006_out0;
wire v$EXP$SAME_1007_out0;
wire v$EXP$SAME_17166_out0;
wire v$EXP$SAME_17167_out0;
wire v$EXP$SAME_3349_out0;
wire v$EXP$SAME_3350_out0;
wire v$EXTHALT_18494_out0;
wire v$EXTHALT_18495_out0;
wire v$EXTHALT_6705_out0;
wire v$EXTHALT_6706_out0;
wire v$E_17993_out0;
wire v$E_17994_out0;
wire v$Error_3949_out0;
wire v$Error_3950_out0;
wire v$F0_16438_out0;
wire v$F0_16439_out0;
wire v$F1_3687_out0;
wire v$F1_3688_out0;
wire v$F2_12662_out0;
wire v$F2_12663_out0;
wire v$F3_8557_out0;
wire v$F3_8558_out0;
wire v$FINISHED_11360_out0;
wire v$FINISHED_11361_out0;
wire v$FINISHED_12202_out0;
wire v$FINISHED_12203_out0;
wire v$FINISHED_14451_out0;
wire v$FINISHED_14452_out0;
wire v$FINISHED_19280_out0;
wire v$FINISHED_19281_out0;
wire v$FINISHED_2461_out0;
wire v$FINISHED_2462_out0;
wire v$FINISHED_7284_out0;
wire v$FINISHED_7285_out0;
wire v$FINISHED_8327_out0;
wire v$FINISHED_8328_out0;
wire v$FMUL$FINISHED$VIEWER_3381_out0;
wire v$FMUL$FINISHED$VIEWER_3382_out0;
wire v$FMUL$FINISHED_15076_out0;
wire v$FMUL$FINISHED_15077_out0;
wire v$FMUL$FINISHED_202_out0;
wire v$FMUL$FINISHED_203_out0;
wire v$FPU$32$BIT$DATAPATH_18334_out0;
wire v$FPU$32$BIT$DATAPATH_18335_out0;
wire v$FPU$32$BIT$MUL$PIPELINED_3712_out0;
wire v$FPU$32$BIT$MUL$PIPELINED_3713_out0;
wire v$FPU$A$EN_12236_out0;
wire v$FPU$A$EN_12237_out0;
wire v$FPU$LOAD$B_12310_out0;
wire v$FPU$LOAD$B_12311_out0;
wire v$FPU$LOAD$STORE_11486_out0;
wire v$FPU$LOAD$STORE_11487_out0;
wire v$F_2133_out0;
wire v$F_2134_out0;
wire v$G$AB_9464_out0;
wire v$G$AB_9465_out0;
wire v$G$AB_9466_out0;
wire v$G$AB_9467_out0;
wire v$G$AB_9468_out0;
wire v$G$AB_9469_out0;
wire v$G$AB_9470_out0;
wire v$G$AB_9471_out0;
wire v$G$AB_9472_out0;
wire v$G$AB_9473_out0;
wire v$G$AB_9474_out0;
wire v$G$AB_9475_out0;
wire v$G$AB_9476_out0;
wire v$G$AB_9477_out0;
wire v$G$AB_9478_out0;
wire v$G$AB_9479_out0;
wire v$G$AB_9480_out0;
wire v$G$AB_9481_out0;
wire v$G$AB_9482_out0;
wire v$G$AB_9483_out0;
wire v$G$AB_9484_out0;
wire v$G$AB_9485_out0;
wire v$G$AB_9486_out0;
wire v$G$AB_9487_out0;
wire v$G$AB_9488_out0;
wire v$G$AB_9489_out0;
wire v$G$AB_9490_out0;
wire v$G$AB_9491_out0;
wire v$G$AB_9492_out0;
wire v$G$AB_9493_out0;
wire v$G$AB_9494_out0;
wire v$G$AB_9495_out0;
wire v$G$AB_9496_out0;
wire v$G$AB_9497_out0;
wire v$G$AB_9498_out0;
wire v$G$AB_9499_out0;
wire v$G$AB_9500_out0;
wire v$G$AB_9501_out0;
wire v$G$AB_9502_out0;
wire v$G$AB_9503_out0;
wire v$G$AB_9504_out0;
wire v$G$AB_9505_out0;
wire v$G$AB_9506_out0;
wire v$G$AB_9507_out0;
wire v$G$AB_9508_out0;
wire v$G$AB_9509_out0;
wire v$G$AB_9510_out0;
wire v$G$AB_9511_out0;
wire v$G$AB_9512_out0;
wire v$G$AB_9513_out0;
wire v$G$AB_9514_out0;
wire v$G$AB_9515_out0;
wire v$G$AB_9516_out0;
wire v$G$AB_9517_out0;
wire v$G$AB_9518_out0;
wire v$G$AB_9519_out0;
wire v$G$AB_9520_out0;
wire v$G$AB_9521_out0;
wire v$G$AB_9522_out0;
wire v$G$AB_9523_out0;
wire v$G$AB_9524_out0;
wire v$G$AB_9525_out0;
wire v$G$AB_9526_out0;
wire v$G$AB_9527_out0;
wire v$G$AB_9528_out0;
wire v$G$AB_9529_out0;
wire v$G$AB_9530_out0;
wire v$G$AB_9531_out0;
wire v$G$AB_9532_out0;
wire v$G$AB_9533_out0;
wire v$G$AB_9534_out0;
wire v$G$AB_9535_out0;
wire v$G$AB_9536_out0;
wire v$G$AB_9537_out0;
wire v$G$AB_9538_out0;
wire v$G$AB_9539_out0;
wire v$G$AB_9540_out0;
wire v$G$AB_9541_out0;
wire v$G$AB_9542_out0;
wire v$G$AB_9543_out0;
wire v$G$AB_9544_out0;
wire v$G$AB_9545_out0;
wire v$G$AB_9546_out0;
wire v$G$AB_9547_out0;
wire v$G$AB_9548_out0;
wire v$G$AB_9549_out0;
wire v$G$AB_9550_out0;
wire v$G$AB_9551_out0;
wire v$G$AB_9552_out0;
wire v$G$AB_9553_out0;
wire v$G$AB_9554_out0;
wire v$G$AB_9555_out0;
wire v$G$AB_9556_out0;
wire v$G$AB_9557_out0;
wire v$G$AB_9558_out0;
wire v$G$AB_9559_out0;
wire v$G$AB_9560_out0;
wire v$G$AB_9561_out0;
wire v$G$AB_9562_out0;
wire v$G$AB_9563_out0;
wire v$G$AB_9564_out0;
wire v$G$AB_9565_out0;
wire v$G$AB_9566_out0;
wire v$G$AB_9567_out0;
wire v$G$AB_9568_out0;
wire v$G$AB_9569_out0;
wire v$G$AB_9570_out0;
wire v$G$AB_9571_out0;
wire v$G$AB_9572_out0;
wire v$G$AB_9573_out0;
wire v$G$AB_9574_out0;
wire v$G$AB_9575_out0;
wire v$G$AB_9576_out0;
wire v$G$AB_9577_out0;
wire v$G$AB_9578_out0;
wire v$G$AB_9579_out0;
wire v$G$AB_9580_out0;
wire v$G$AB_9581_out0;
wire v$G$AB_9582_out0;
wire v$G$AB_9583_out0;
wire v$G$AB_9584_out0;
wire v$G$AB_9585_out0;
wire v$G$AB_9586_out0;
wire v$G$AB_9587_out0;
wire v$G$AB_9588_out0;
wire v$G$AB_9589_out0;
wire v$G$AB_9590_out0;
wire v$G$AB_9591_out0;
wire v$G$AB_9592_out0;
wire v$G$AB_9593_out0;
wire v$G$AB_9594_out0;
wire v$G$AB_9595_out0;
wire v$G$AB_9596_out0;
wire v$G$AB_9597_out0;
wire v$G$AB_9598_out0;
wire v$G$AB_9599_out0;
wire v$G$AB_9600_out0;
wire v$G$AB_9601_out0;
wire v$G$AB_9602_out0;
wire v$G$AB_9603_out0;
wire v$G$AB_9604_out0;
wire v$G$AB_9605_out0;
wire v$G$AB_9606_out0;
wire v$G$AB_9607_out0;
wire v$G$AB_9608_out0;
wire v$G$AB_9609_out0;
wire v$G$AB_9610_out0;
wire v$G$AB_9611_out0;
wire v$G$AB_9612_out0;
wire v$G$AB_9613_out0;
wire v$G$AB_9614_out0;
wire v$G$AB_9615_out0;
wire v$G$AB_9616_out0;
wire v$G$AB_9617_out0;
wire v$G$AB_9618_out0;
wire v$G$AB_9619_out0;
wire v$G$AB_9620_out0;
wire v$G$AB_9621_out0;
wire v$G$AB_9622_out0;
wire v$G$AB_9623_out0;
wire v$G$AB_9624_out0;
wire v$G$AB_9625_out0;
wire v$G$AB_9626_out0;
wire v$G$AB_9627_out0;
wire v$G$AB_9628_out0;
wire v$G$AB_9629_out0;
wire v$G$AB_9630_out0;
wire v$G$AB_9631_out0;
wire v$G$AB_9632_out0;
wire v$G$AB_9633_out0;
wire v$G$AB_9634_out0;
wire v$G$AB_9635_out0;
wire v$G$AB_9636_out0;
wire v$G$AB_9637_out0;
wire v$G$AB_9638_out0;
wire v$G$AB_9639_out0;
wire v$G$AB_9640_out0;
wire v$G$AB_9641_out0;
wire v$G$AB_9642_out0;
wire v$G$AB_9643_out0;
wire v$G$AB_9644_out0;
wire v$G$AB_9645_out0;
wire v$G$AB_9646_out0;
wire v$G$AB_9647_out0;
wire v$G$AB_9648_out0;
wire v$G$AB_9649_out0;
wire v$G$AB_9650_out0;
wire v$G$AB_9651_out0;
wire v$G$AB_9652_out0;
wire v$G$AB_9653_out0;
wire v$G$AB_9654_out0;
wire v$G$AB_9655_out0;
wire v$G$AB_9656_out0;
wire v$G$AB_9657_out0;
wire v$G$AB_9658_out0;
wire v$G$AB_9659_out0;
wire v$G$AB_9660_out0;
wire v$G$AB_9661_out0;
wire v$G$AB_9662_out0;
wire v$G$AB_9663_out0;
wire v$G$AB_9664_out0;
wire v$G$AB_9665_out0;
wire v$G$AB_9666_out0;
wire v$G$AB_9667_out0;
wire v$G$AB_9668_out0;
wire v$G$AB_9669_out0;
wire v$G$AB_9670_out0;
wire v$G$AB_9671_out0;
wire v$G$AB_9672_out0;
wire v$G$AB_9673_out0;
wire v$G$AB_9674_out0;
wire v$G$AB_9675_out0;
wire v$G$AB_9676_out0;
wire v$G$AB_9677_out0;
wire v$G$AB_9678_out0;
wire v$G$AB_9679_out0;
wire v$G$AB_9680_out0;
wire v$G$AB_9681_out0;
wire v$G$AB_9682_out0;
wire v$G$AB_9683_out0;
wire v$G$AB_9684_out0;
wire v$G$AB_9685_out0;
wire v$G$AB_9686_out0;
wire v$G$AB_9687_out0;
wire v$G$AB_9688_out0;
wire v$G$AB_9689_out0;
wire v$G$AB_9690_out0;
wire v$G$AB_9691_out0;
wire v$G$AB_9692_out0;
wire v$G$AB_9693_out0;
wire v$G$AB_9694_out0;
wire v$G$AB_9695_out0;
wire v$G$AB_9696_out0;
wire v$G$AB_9697_out0;
wire v$G$AB_9698_out0;
wire v$G$AB_9699_out0;
wire v$G$AB_9700_out0;
wire v$G$AB_9701_out0;
wire v$G$AB_9702_out0;
wire v$G$AB_9703_out0;
wire v$G$AB_9704_out0;
wire v$G$AB_9705_out0;
wire v$G$AB_9706_out0;
wire v$G$AB_9707_out0;
wire v$G$AB_9708_out0;
wire v$G$AB_9709_out0;
wire v$G$AD_17684_out0;
wire v$G$AD_17685_out0;
wire v$G$AD_17686_out0;
wire v$G$AD_17687_out0;
wire v$G$AD_17688_out0;
wire v$G$AD_17689_out0;
wire v$G$AD_17690_out0;
wire v$G$AD_17691_out0;
wire v$G$AD_17692_out0;
wire v$G$AD_17693_out0;
wire v$G$AD_17694_out0;
wire v$G$AD_17695_out0;
wire v$G$AD_17696_out0;
wire v$G$AD_17697_out0;
wire v$G$AD_17698_out0;
wire v$G$AD_17699_out0;
wire v$G$AD_17700_out0;
wire v$G$AD_17701_out0;
wire v$G$AD_17702_out0;
wire v$G$AD_17703_out0;
wire v$G$AD_17704_out0;
wire v$G$AD_17705_out0;
wire v$G$AD_17706_out0;
wire v$G$AD_17707_out0;
wire v$G$AD_17708_out0;
wire v$G$AD_17709_out0;
wire v$G$AD_17710_out0;
wire v$G$AD_17711_out0;
wire v$G$AD_17712_out0;
wire v$G$AD_17713_out0;
wire v$G$AD_17714_out0;
wire v$G$AD_17715_out0;
wire v$G$AD_17716_out0;
wire v$G$AD_17717_out0;
wire v$G$AD_17718_out0;
wire v$G$AD_17719_out0;
wire v$G$AD_17720_out0;
wire v$G$AD_17721_out0;
wire v$G$AD_17722_out0;
wire v$G$AD_17723_out0;
wire v$G$AD_17724_out0;
wire v$G$AD_17725_out0;
wire v$G$AD_17726_out0;
wire v$G$AD_17727_out0;
wire v$G$AD_17728_out0;
wire v$G$AD_17729_out0;
wire v$G$AD_17730_out0;
wire v$G$AD_17731_out0;
wire v$G$AD_17732_out0;
wire v$G$AD_17733_out0;
wire v$G$AD_17734_out0;
wire v$G$AD_17735_out0;
wire v$G$AD_17736_out0;
wire v$G$AD_17737_out0;
wire v$G$AD_17738_out0;
wire v$G$AD_17739_out0;
wire v$G$AD_17740_out0;
wire v$G$AD_17741_out0;
wire v$G$AD_17742_out0;
wire v$G$AD_17743_out0;
wire v$G$AD_17744_out0;
wire v$G$AD_17745_out0;
wire v$G$AD_17746_out0;
wire v$G$AD_17747_out0;
wire v$G$AD_17748_out0;
wire v$G$AD_17749_out0;
wire v$G$AD_17750_out0;
wire v$G$AD_17751_out0;
wire v$G$AD_17752_out0;
wire v$G$AD_17753_out0;
wire v$G$AD_17754_out0;
wire v$G$AD_17755_out0;
wire v$G$AD_17756_out0;
wire v$G$AD_17757_out0;
wire v$G$AD_17758_out0;
wire v$G$AD_17759_out0;
wire v$G$AD_17760_out0;
wire v$G$AD_17761_out0;
wire v$G$AD_17762_out0;
wire v$G$AD_17763_out0;
wire v$G$AD_17764_out0;
wire v$G$AD_17765_out0;
wire v$G$AD_17766_out0;
wire v$G$AD_17767_out0;
wire v$G$AD_17768_out0;
wire v$G$AD_17769_out0;
wire v$G$AD_17770_out0;
wire v$G$AD_17771_out0;
wire v$G$AD_17772_out0;
wire v$G$AD_17773_out0;
wire v$G$AD_17774_out0;
wire v$G$AD_17775_out0;
wire v$G$AD_17776_out0;
wire v$G$AD_17777_out0;
wire v$G$AD_17778_out0;
wire v$G$AD_17779_out0;
wire v$G$AD_17780_out0;
wire v$G$AD_17781_out0;
wire v$G$AD_17782_out0;
wire v$G$AD_17783_out0;
wire v$G$AD_17784_out0;
wire v$G$AD_17785_out0;
wire v$G$AD_17786_out0;
wire v$G$AD_17787_out0;
wire v$G$AD_17788_out0;
wire v$G$AD_17789_out0;
wire v$G$AD_17790_out0;
wire v$G$AD_17791_out0;
wire v$G$AD_17792_out0;
wire v$G$AD_17793_out0;
wire v$G$AD_17794_out0;
wire v$G$AD_17795_out0;
wire v$G$AD_17796_out0;
wire v$G$AD_17797_out0;
wire v$G$AD_17798_out0;
wire v$G$AD_17799_out0;
wire v$G$AD_17800_out0;
wire v$G$AD_17801_out0;
wire v$G$AD_17802_out0;
wire v$G$AD_17803_out0;
wire v$G$AD_17804_out0;
wire v$G$AD_17805_out0;
wire v$G$AD_17806_out0;
wire v$G$AD_17807_out0;
wire v$G$AD_17808_out0;
wire v$G$AD_17809_out0;
wire v$G$AD_17810_out0;
wire v$G$AD_17811_out0;
wire v$G$AD_17812_out0;
wire v$G$AD_17813_out0;
wire v$G$AD_17814_out0;
wire v$G$AD_17815_out0;
wire v$G$AD_17816_out0;
wire v$G$AD_17817_out0;
wire v$G$AD_17818_out0;
wire v$G$AD_17819_out0;
wire v$G$AD_17820_out0;
wire v$G$AD_17821_out0;
wire v$G$AD_17822_out0;
wire v$G$AD_17823_out0;
wire v$G$AD_17824_out0;
wire v$G$AD_17825_out0;
wire v$G$AD_17826_out0;
wire v$G$AD_17827_out0;
wire v$G$AD_17828_out0;
wire v$G$AD_17829_out0;
wire v$G$AD_17830_out0;
wire v$G$AD_17831_out0;
wire v$G$AD_17832_out0;
wire v$G$AD_17833_out0;
wire v$G$AD_17834_out0;
wire v$G$AD_17835_out0;
wire v$G$AD_17836_out0;
wire v$G$AD_17837_out0;
wire v$G$AD_17838_out0;
wire v$G$AD_17839_out0;
wire v$G$AD_17840_out0;
wire v$G$AD_17841_out0;
wire v$G$AD_17842_out0;
wire v$G$AD_17843_out0;
wire v$G$AD_17844_out0;
wire v$G$AD_17845_out0;
wire v$G$AD_17846_out0;
wire v$G$AD_17847_out0;
wire v$G$AD_17848_out0;
wire v$G$AD_17849_out0;
wire v$G$AD_17850_out0;
wire v$G$AD_17851_out0;
wire v$G$AD_17852_out0;
wire v$G$AD_17853_out0;
wire v$G$AD_17854_out0;
wire v$G$AD_17855_out0;
wire v$G$AD_17856_out0;
wire v$G$AD_17857_out0;
wire v$G$AD_17858_out0;
wire v$G$AD_17859_out0;
wire v$G$AD_17860_out0;
wire v$G$AD_17861_out0;
wire v$G$AD_17862_out0;
wire v$G$AD_17863_out0;
wire v$G$AD_17864_out0;
wire v$G$AD_17865_out0;
wire v$G$AD_17866_out0;
wire v$G$AD_17867_out0;
wire v$G$AD_17868_out0;
wire v$G$AD_17869_out0;
wire v$G$AD_17870_out0;
wire v$G$AD_17871_out0;
wire v$G$AD_17872_out0;
wire v$G$AD_17873_out0;
wire v$G$AD_17874_out0;
wire v$G$AD_17875_out0;
wire v$G$AD_17876_out0;
wire v$G$AD_17877_out0;
wire v$G$AD_17878_out0;
wire v$G$AD_17879_out0;
wire v$G$AD_17880_out0;
wire v$G$AD_17881_out0;
wire v$G$AD_17882_out0;
wire v$G$AD_17883_out0;
wire v$G$AD_17884_out0;
wire v$G$AD_17885_out0;
wire v$G$AD_17886_out0;
wire v$G$AD_17887_out0;
wire v$G$AD_17888_out0;
wire v$G$AD_17889_out0;
wire v$G$AD_17890_out0;
wire v$G$AD_17891_out0;
wire v$G$AD_17892_out0;
wire v$G$AD_17893_out0;
wire v$G$AD_17894_out0;
wire v$G$AD_17895_out0;
wire v$G$AD_17896_out0;
wire v$G$AD_17897_out0;
wire v$G$AD_17898_out0;
wire v$G$AD_17899_out0;
wire v$G$AD_17900_out0;
wire v$G$AD_17901_out0;
wire v$G$AD_17902_out0;
wire v$G$AD_17903_out0;
wire v$G$AD_17904_out0;
wire v$G$AD_17905_out0;
wire v$G$AD_17906_out0;
wire v$G$AD_17907_out0;
wire v$G$AD_17908_out0;
wire v$G$AD_17909_out0;
wire v$G$AD_17910_out0;
wire v$G$AD_17911_out0;
wire v$G$AD_17912_out0;
wire v$G$AD_17913_out0;
wire v$G$AD_17914_out0;
wire v$G$AD_17915_out0;
wire v$G$AD_17916_out0;
wire v$G$AD_17917_out0;
wire v$G$AD_17918_out0;
wire v$G$AD_17919_out0;
wire v$G$AD_17920_out0;
wire v$G$AD_17921_out0;
wire v$G$AD_17922_out0;
wire v$G$AD_17923_out0;
wire v$G$AD_17924_out0;
wire v$G$AD_17925_out0;
wire v$G$AD_17926_out0;
wire v$G$AD_17927_out0;
wire v$G$AD_17928_out0;
wire v$G$AD_17929_out0;
wire v$G$CD_1017_out0;
wire v$G$CD_1018_out0;
wire v$G$CD_1019_out0;
wire v$G$CD_1020_out0;
wire v$G$CD_1021_out0;
wire v$G$CD_1022_out0;
wire v$G$CD_1023_out0;
wire v$G$CD_1024_out0;
wire v$G$CD_1025_out0;
wire v$G$CD_1026_out0;
wire v$G$CD_1027_out0;
wire v$G$CD_1028_out0;
wire v$G$CD_1029_out0;
wire v$G$CD_1030_out0;
wire v$G$CD_1031_out0;
wire v$G$CD_1032_out0;
wire v$G$CD_1033_out0;
wire v$G$CD_1034_out0;
wire v$G$CD_1035_out0;
wire v$G$CD_1036_out0;
wire v$G$CD_1037_out0;
wire v$G$CD_1038_out0;
wire v$G$CD_1039_out0;
wire v$G$CD_1040_out0;
wire v$G$CD_1041_out0;
wire v$G$CD_1042_out0;
wire v$G$CD_1043_out0;
wire v$G$CD_1044_out0;
wire v$G$CD_1045_out0;
wire v$G$CD_1046_out0;
wire v$G$CD_1047_out0;
wire v$G$CD_1048_out0;
wire v$G$CD_1049_out0;
wire v$G$CD_1050_out0;
wire v$G$CD_1051_out0;
wire v$G$CD_1052_out0;
wire v$G$CD_1053_out0;
wire v$G$CD_1054_out0;
wire v$G$CD_1055_out0;
wire v$G$CD_1056_out0;
wire v$G$CD_1057_out0;
wire v$G$CD_1058_out0;
wire v$G$CD_1059_out0;
wire v$G$CD_1060_out0;
wire v$G$CD_1061_out0;
wire v$G$CD_1062_out0;
wire v$G$CD_1063_out0;
wire v$G$CD_1064_out0;
wire v$G$CD_1065_out0;
wire v$G$CD_1066_out0;
wire v$G$CD_1067_out0;
wire v$G$CD_1068_out0;
wire v$G$CD_1069_out0;
wire v$G$CD_1070_out0;
wire v$G$CD_1071_out0;
wire v$G$CD_1072_out0;
wire v$G$CD_1073_out0;
wire v$G$CD_1074_out0;
wire v$G$CD_1075_out0;
wire v$G$CD_1076_out0;
wire v$G$CD_1077_out0;
wire v$G$CD_1078_out0;
wire v$G$CD_1079_out0;
wire v$G$CD_1080_out0;
wire v$G$CD_1081_out0;
wire v$G$CD_1082_out0;
wire v$G$CD_1083_out0;
wire v$G$CD_1084_out0;
wire v$G$CD_1085_out0;
wire v$G$CD_1086_out0;
wire v$G$CD_1087_out0;
wire v$G$CD_1088_out0;
wire v$G$CD_1089_out0;
wire v$G$CD_1090_out0;
wire v$G$CD_1091_out0;
wire v$G$CD_1092_out0;
wire v$G$CD_1093_out0;
wire v$G$CD_1094_out0;
wire v$G$CD_1095_out0;
wire v$G$CD_1096_out0;
wire v$G$CD_1097_out0;
wire v$G$CD_1098_out0;
wire v$G$CD_1099_out0;
wire v$G$CD_1100_out0;
wire v$G$CD_1101_out0;
wire v$G$CD_1102_out0;
wire v$G$CD_1103_out0;
wire v$G$CD_1104_out0;
wire v$G$CD_1105_out0;
wire v$G$CD_1106_out0;
wire v$G$CD_1107_out0;
wire v$G$CD_1108_out0;
wire v$G$CD_1109_out0;
wire v$G$CD_1110_out0;
wire v$G$CD_1111_out0;
wire v$G$CD_1112_out0;
wire v$G$CD_1113_out0;
wire v$G$CD_1114_out0;
wire v$G$CD_1115_out0;
wire v$G$CD_1116_out0;
wire v$G$CD_1117_out0;
wire v$G$CD_1118_out0;
wire v$G$CD_1119_out0;
wire v$G$CD_1120_out0;
wire v$G$CD_1121_out0;
wire v$G$CD_1122_out0;
wire v$G$CD_1123_out0;
wire v$G$CD_1124_out0;
wire v$G$CD_1125_out0;
wire v$G$CD_1126_out0;
wire v$G$CD_1127_out0;
wire v$G$CD_1128_out0;
wire v$G$CD_1129_out0;
wire v$G$CD_1130_out0;
wire v$G$CD_1131_out0;
wire v$G$CD_1132_out0;
wire v$G$CD_1133_out0;
wire v$G$CD_1134_out0;
wire v$G$CD_1135_out0;
wire v$G$CD_1136_out0;
wire v$G$CD_1137_out0;
wire v$G$CD_1138_out0;
wire v$G$CD_1139_out0;
wire v$G$CD_1140_out0;
wire v$G$CD_1141_out0;
wire v$G$CD_1142_out0;
wire v$G$CD_1143_out0;
wire v$G$CD_1144_out0;
wire v$G$CD_1145_out0;
wire v$G$CD_1146_out0;
wire v$G$CD_1147_out0;
wire v$G$CD_1148_out0;
wire v$G$CD_1149_out0;
wire v$G$CD_1150_out0;
wire v$G$CD_1151_out0;
wire v$G$CD_1152_out0;
wire v$G$CD_1153_out0;
wire v$G$CD_1154_out0;
wire v$G$CD_1155_out0;
wire v$G$CD_1156_out0;
wire v$G$CD_1157_out0;
wire v$G$CD_1158_out0;
wire v$G$CD_1159_out0;
wire v$G$CD_1160_out0;
wire v$G$CD_1161_out0;
wire v$G$CD_1162_out0;
wire v$G$CD_1163_out0;
wire v$G$CD_1164_out0;
wire v$G$CD_1165_out0;
wire v$G$CD_1166_out0;
wire v$G$CD_1167_out0;
wire v$G$CD_1168_out0;
wire v$G$CD_1169_out0;
wire v$G$CD_1170_out0;
wire v$G$CD_1171_out0;
wire v$G$CD_1172_out0;
wire v$G$CD_1173_out0;
wire v$G$CD_1174_out0;
wire v$G$CD_1175_out0;
wire v$G$CD_1176_out0;
wire v$G$CD_1177_out0;
wire v$G$CD_1178_out0;
wire v$G$CD_1179_out0;
wire v$G$CD_1180_out0;
wire v$G$CD_1181_out0;
wire v$G$CD_1182_out0;
wire v$G$CD_1183_out0;
wire v$G$CD_1184_out0;
wire v$G$CD_1185_out0;
wire v$G$CD_1186_out0;
wire v$G$CD_1187_out0;
wire v$G$CD_1188_out0;
wire v$G$CD_1189_out0;
wire v$G$CD_1190_out0;
wire v$G$CD_1191_out0;
wire v$G$CD_1192_out0;
wire v$G$CD_1193_out0;
wire v$G$CD_1194_out0;
wire v$G$CD_1195_out0;
wire v$G$CD_1196_out0;
wire v$G$CD_1197_out0;
wire v$G$CD_1198_out0;
wire v$G$CD_1199_out0;
wire v$G$CD_1200_out0;
wire v$G$CD_1201_out0;
wire v$G$CD_1202_out0;
wire v$G$CD_1203_out0;
wire v$G$CD_1204_out0;
wire v$G$CD_1205_out0;
wire v$G$CD_1206_out0;
wire v$G$CD_1207_out0;
wire v$G$CD_1208_out0;
wire v$G$CD_1209_out0;
wire v$G$CD_1210_out0;
wire v$G$CD_1211_out0;
wire v$G$CD_1212_out0;
wire v$G$CD_1213_out0;
wire v$G$CD_1214_out0;
wire v$G$CD_1215_out0;
wire v$G$CD_1216_out0;
wire v$G$CD_1217_out0;
wire v$G$CD_1218_out0;
wire v$G$CD_1219_out0;
wire v$G$CD_1220_out0;
wire v$G$CD_1221_out0;
wire v$G$CD_1222_out0;
wire v$G$CD_1223_out0;
wire v$G$CD_1224_out0;
wire v$G$CD_1225_out0;
wire v$G$CD_1226_out0;
wire v$G$CD_1227_out0;
wire v$G$CD_1228_out0;
wire v$G$CD_1229_out0;
wire v$G$CD_1230_out0;
wire v$G$CD_1231_out0;
wire v$G$CD_1232_out0;
wire v$G$CD_1233_out0;
wire v$G$CD_1234_out0;
wire v$G$CD_1235_out0;
wire v$G$CD_1236_out0;
wire v$G$CD_1237_out0;
wire v$G$CD_1238_out0;
wire v$G$CD_1239_out0;
wire v$G$CD_1240_out0;
wire v$G$CD_1241_out0;
wire v$G$CD_1242_out0;
wire v$G$CD_1243_out0;
wire v$G$CD_1244_out0;
wire v$G$CD_1245_out0;
wire v$G$CD_1246_out0;
wire v$G$CD_1247_out0;
wire v$G$CD_1248_out0;
wire v$G$CD_1249_out0;
wire v$G$CD_1250_out0;
wire v$G$CD_1251_out0;
wire v$G$CD_1252_out0;
wire v$G$CD_1253_out0;
wire v$G$CD_1254_out0;
wire v$G$CD_1255_out0;
wire v$G$CD_1256_out0;
wire v$G$CD_1257_out0;
wire v$G$CD_1258_out0;
wire v$G$CD_1259_out0;
wire v$G$CD_1260_out0;
wire v$G$CD_1261_out0;
wire v$G$CD_1262_out0;
wire v$G0_16548_out0;
wire v$G0_16549_out0;
wire v$G0_16550_out0;
wire v$G0_16551_out0;
wire v$G0_16552_out0;
wire v$G0_16553_out0;
wire v$G10_10725_out0;
wire v$G10_10726_out0;
wire v$G10_1329_out0;
wire v$G10_1330_out0;
wire v$G10_13900_out0;
wire v$G10_13901_out0;
wire v$G10_15166_out0;
wire v$G10_15167_out0;
wire v$G10_15189_out0;
wire v$G10_15190_out0;
wire v$G10_1543_out0;
wire v$G10_1544_out0;
wire v$G10_1545_out0;
wire v$G10_1546_out0;
wire v$G10_1547_out0;
wire v$G10_1548_out0;
wire v$G10_1549_out0;
wire v$G10_15507_out0;
wire v$G10_15508_out0;
wire v$G10_1550_out0;
wire v$G10_1551_out0;
wire v$G10_1552_out0;
wire v$G10_1553_out0;
wire v$G10_1554_out0;
wire v$G10_1555_out0;
wire v$G10_1556_out0;
wire v$G10_1557_out0;
wire v$G10_1558_out0;
wire v$G10_1559_out0;
wire v$G10_1560_out0;
wire v$G10_1561_out0;
wire v$G10_1562_out0;
wire v$G10_1563_out0;
wire v$G10_1564_out0;
wire v$G10_1565_out0;
wire v$G10_1566_out0;
wire v$G10_1567_out0;
wire v$G10_1568_out0;
wire v$G10_1569_out0;
wire v$G10_1570_out0;
wire v$G10_1571_out0;
wire v$G10_1572_out0;
wire v$G10_1573_out0;
wire v$G10_1574_out0;
wire v$G10_1575_out0;
wire v$G10_1576_out0;
wire v$G10_1577_out0;
wire v$G10_1578_out0;
wire v$G10_17126_out0;
wire v$G10_17127_out0;
wire v$G10_18785_out0;
wire v$G10_18786_out0;
wire v$G10_19095_out0;
wire v$G10_19096_out0;
wire v$G10_1993_out0;
wire v$G10_1994_out0;
wire v$G10_1995_out0;
wire v$G10_1996_out0;
wire v$G10_1997_out0;
wire v$G10_1998_out0;
wire v$G10_2161_out0;
wire v$G10_2162_out0;
wire v$G10_3112_out0;
wire v$G10_3113_out0;
wire v$G10_3985_out0;
wire v$G10_3986_out0;
wire v$G10_6926_out0;
wire v$G10_6927_out0;
wire v$G11_11575_out0;
wire v$G11_11576_out0;
wire v$G11_11577_out0;
wire v$G11_11578_out0;
wire v$G11_11579_out0;
wire v$G11_11580_out0;
wire v$G11_12417_out0;
wire v$G11_12418_out0;
wire v$G11_13991_out0;
wire v$G11_13992_out0;
wire v$G11_15185_out0;
wire v$G11_15186_out0;
wire v$G11_16230_out0;
wire v$G11_16231_out0;
wire v$G11_16232_out0;
wire v$G11_16233_out0;
wire v$G11_16234_out0;
wire v$G11_16235_out0;
wire v$G11_16236_out0;
wire v$G11_16237_out0;
wire v$G11_16238_out0;
wire v$G11_16239_out0;
wire v$G11_16240_out0;
wire v$G11_16241_out0;
wire v$G11_16242_out0;
wire v$G11_16243_out0;
wire v$G11_16244_out0;
wire v$G11_16245_out0;
wire v$G11_16246_out0;
wire v$G11_16247_out0;
wire v$G11_16248_out0;
wire v$G11_16249_out0;
wire v$G11_16250_out0;
wire v$G11_16251_out0;
wire v$G11_16252_out0;
wire v$G11_16253_out0;
wire v$G11_1775_out0;
wire v$G11_1776_out0;
wire v$G11_18621_out0;
wire v$G11_18622_out0;
wire v$G11_2491_out0;
wire v$G11_2492_out0;
wire v$G11_3188_out0;
wire v$G11_3189_out0;
wire v$G11_3223_out0;
wire v$G11_3224_out0;
wire v$G11_3475_out0;
wire v$G11_3476_out0;
wire v$G11_5080_out0;
wire v$G11_5081_out0;
wire v$G11_8511_out0;
wire v$G11_8512_out0;
wire v$G11_8539_out0;
wire v$G11_8540_out0;
wire v$G11_8572_out0;
wire v$G11_8573_out0;
wire v$G11_9189_out0;
wire v$G11_9190_out0;
wire v$G11_9191_out0;
wire v$G11_9192_out0;
wire v$G11_9193_out0;
wire v$G11_9194_out0;
wire v$G11_9195_out0;
wire v$G11_9196_out0;
wire v$G11_9197_out0;
wire v$G11_9198_out0;
wire v$G11_9199_out0;
wire v$G11_9200_out0;
wire v$G11_9201_out0;
wire v$G11_9202_out0;
wire v$G11_9203_out0;
wire v$G11_9204_out0;
wire v$G11_9205_out0;
wire v$G11_9206_out0;
wire v$G11_9207_out0;
wire v$G11_9208_out0;
wire v$G11_9209_out0;
wire v$G11_9210_out0;
wire v$G11_9211_out0;
wire v$G11_9212_out0;
wire v$G11_9213_out0;
wire v$G11_9214_out0;
wire v$G11_9215_out0;
wire v$G11_9216_out0;
wire v$G11_9217_out0;
wire v$G11_9218_out0;
wire v$G11_9219_out0;
wire v$G11_9220_out0;
wire v$G11_9221_out0;
wire v$G11_9222_out0;
wire v$G11_9223_out0;
wire v$G11_9224_out0;
wire v$G11_9984_out0;
wire v$G11_9985_out0;
wire v$G12_10366_out0;
wire v$G12_10367_out0;
wire v$G12_12470_out0;
wire v$G12_12471_out0;
wire v$G12_12555_out0;
wire v$G12_12556_out0;
wire v$G12_14383_out0;
wire v$G12_14384_out0;
wire v$G12_15311_out0;
wire v$G12_15312_out0;
wire v$G12_16862_out0;
wire v$G12_16863_out0;
wire v$G12_17094_out0;
wire v$G12_17095_out0;
wire v$G12_17096_out0;
wire v$G12_17097_out0;
wire v$G12_17098_out0;
wire v$G12_17099_out0;
wire v$G12_17100_out0;
wire v$G12_17101_out0;
wire v$G12_17102_out0;
wire v$G12_17103_out0;
wire v$G12_17104_out0;
wire v$G12_17105_out0;
wire v$G12_17106_out0;
wire v$G12_17107_out0;
wire v$G12_17108_out0;
wire v$G12_17109_out0;
wire v$G12_17110_out0;
wire v$G12_17111_out0;
wire v$G12_17112_out0;
wire v$G12_17113_out0;
wire v$G12_17114_out0;
wire v$G12_17115_out0;
wire v$G12_17116_out0;
wire v$G12_17117_out0;
wire v$G12_1981_out0;
wire v$G12_1982_out0;
wire v$G12_2420_out0;
wire v$G12_2421_out0;
wire v$G12_3804_out0;
wire v$G12_3805_out0;
wire v$G12_5046_out0;
wire v$G12_5047_out0;
wire v$G12_6432_out0;
wire v$G12_6433_out0;
wire v$G12_7327_out0;
wire v$G12_7328_out0;
wire v$G12_7329_out0;
wire v$G12_7330_out0;
wire v$G12_7331_out0;
wire v$G12_7332_out0;
wire v$G13_10681_out0;
wire v$G13_10682_out0;
wire v$G13_12722_out0;
wire v$G13_12723_out0;
wire v$G13_14029_out0;
wire v$G13_14030_out0;
wire v$G13_15463_out0;
wire v$G13_15464_out0;
wire v$G13_15713_out0;
wire v$G13_15714_out0;
wire v$G13_17152_out0;
wire v$G13_17153_out0;
wire v$G13_1847_out0;
wire v$G13_1848_out0;
wire v$G13_200_out0;
wire v$G13_201_out0;
wire v$G13_3052_out0;
wire v$G13_3053_out0;
wire v$G13_3054_out0;
wire v$G13_3055_out0;
wire v$G13_3056_out0;
wire v$G13_3057_out0;
wire v$G13_4516_out0;
wire v$G13_4517_out0;
wire v$G13_4564_out0;
wire v$G13_4565_out0;
wire v$G13_4566_out0;
wire v$G13_4567_out0;
wire v$G13_4568_out0;
wire v$G13_4569_out0;
wire v$G13_4570_out0;
wire v$G13_4571_out0;
wire v$G13_4572_out0;
wire v$G13_4573_out0;
wire v$G13_4574_out0;
wire v$G13_4575_out0;
wire v$G13_4576_out0;
wire v$G13_4577_out0;
wire v$G13_4578_out0;
wire v$G13_4579_out0;
wire v$G13_4580_out0;
wire v$G13_4581_out0;
wire v$G13_4582_out0;
wire v$G13_4583_out0;
wire v$G13_4584_out0;
wire v$G13_4585_out0;
wire v$G13_4586_out0;
wire v$G13_4587_out0;
wire v$G13_8221_out0;
wire v$G13_8222_out0;
wire v$G14_12611_out0;
wire v$G14_12612_out0;
wire v$G14_13227_out0;
wire v$G14_13228_out0;
wire v$G14_13229_out0;
wire v$G14_13230_out0;
wire v$G14_15285_out0;
wire v$G14_15286_out0;
wire v$G14_15875_out0;
wire v$G14_15876_out0;
wire v$G14_16418_out0;
wire v$G14_16419_out0;
wire v$G14_17632_out0;
wire v$G14_17633_out0;
wire v$G14_1831_out0;
wire v$G14_1832_out0;
wire v$G14_18593_out0;
wire v$G14_18594_out0;
wire v$G14_18595_out0;
wire v$G14_18596_out0;
wire v$G14_18597_out0;
wire v$G14_18598_out0;
wire v$G14_19043_out0;
wire v$G14_19044_out0;
wire v$G14_5346_out0;
wire v$G14_5347_out0;
wire v$G14_5626_out0;
wire v$G14_5627_out0;
wire v$G14_6392_out0;
wire v$G14_6393_out0;
wire v$G14_6671_out0;
wire v$G14_6672_out0;
wire v$G15_11541_out0;
wire v$G15_11542_out0;
wire v$G15_11543_out0;
wire v$G15_11544_out0;
wire v$G15_11545_out0;
wire v$G15_11546_out0;
wire v$G15_13976_out0;
wire v$G15_13977_out0;
wire v$G15_14005_out0;
wire v$G15_14006_out0;
wire v$G15_14180_out0;
wire v$G15_14181_out0;
wire v$G15_14222_out0;
wire v$G15_14223_out0;
wire v$G15_14224_out0;
wire v$G15_14225_out0;
wire v$G15_14226_out0;
wire v$G15_14227_out0;
wire v$G15_14228_out0;
wire v$G15_14229_out0;
wire v$G15_14230_out0;
wire v$G15_14231_out0;
wire v$G15_14232_out0;
wire v$G15_14233_out0;
wire v$G15_14234_out0;
wire v$G15_14235_out0;
wire v$G15_14236_out0;
wire v$G15_14237_out0;
wire v$G15_14238_out0;
wire v$G15_14239_out0;
wire v$G15_14240_out0;
wire v$G15_14241_out0;
wire v$G15_14242_out0;
wire v$G15_14243_out0;
wire v$G15_14244_out0;
wire v$G15_14245_out0;
wire v$G15_15183_out0;
wire v$G15_15184_out0;
wire v$G15_18435_out0;
wire v$G15_18436_out0;
wire v$G15_19147_out0;
wire v$G15_19148_out0;
wire v$G15_2030_out0;
wire v$G15_2031_out0;
wire v$G15_2874_out0;
wire v$G15_2875_out0;
wire v$G15_4364_out0;
wire v$G15_4365_out0;
wire v$G15_5719_out0;
wire v$G15_5720_out0;
wire v$G16_12541_out0;
wire v$G16_12542_out0;
wire v$G16_1476_out0;
wire v$G16_1477_out0;
wire v$G16_17071_out0;
wire v$G16_17072_out0;
wire v$G16_17073_out0;
wire v$G16_17074_out0;
wire v$G16_17075_out0;
wire v$G16_17076_out0;
wire v$G16_17473_out0;
wire v$G16_17474_out0;
wire v$G16_17475_out0;
wire v$G16_17476_out0;
wire v$G16_17477_out0;
wire v$G16_17478_out0;
wire v$G16_17479_out0;
wire v$G16_17480_out0;
wire v$G16_17481_out0;
wire v$G16_17482_out0;
wire v$G16_17483_out0;
wire v$G16_17484_out0;
wire v$G16_17485_out0;
wire v$G16_17486_out0;
wire v$G16_17487_out0;
wire v$G16_17488_out0;
wire v$G16_17489_out0;
wire v$G16_17490_out0;
wire v$G16_17491_out0;
wire v$G16_17492_out0;
wire v$G16_17493_out0;
wire v$G16_17494_out0;
wire v$G16_17495_out0;
wire v$G16_17496_out0;
wire v$G16_17575_out0;
wire v$G16_17576_out0;
wire v$G16_17588_out0;
wire v$G16_17589_out0;
wire v$G16_19392_out0;
wire v$G16_19393_out0;
wire v$G16_3233_out0;
wire v$G16_3234_out0;
wire v$G16_3720_out0;
wire v$G16_3721_out0;
wire v$G16_4639_out0;
wire v$G16_4640_out0;
wire v$G16_6632_out0;
wire v$G16_6633_out0;
wire v$G16_6650_out0;
wire v$G16_6651_out0;
wire v$G17_12250_out0;
wire v$G17_12251_out0;
wire v$G17_12704_out0;
wire v$G17_12705_out0;
wire v$G17_14419_out0;
wire v$G17_14420_out0;
wire v$G17_15402_out0;
wire v$G17_15403_out0;
wire v$G17_381_out0;
wire v$G17_382_out0;
wire v$G17_5699_out0;
wire v$G17_5700_out0;
wire v$G17_5717_out0;
wire v$G17_5718_out0;
wire v$G17_8487_out0;
wire v$G17_8488_out0;
wire v$G17_8489_out0;
wire v$G17_8490_out0;
wire v$G17_8491_out0;
wire v$G17_8492_out0;
wire v$G17_8493_out0;
wire v$G17_8494_out0;
wire v$G17_8495_out0;
wire v$G17_8496_out0;
wire v$G17_8497_out0;
wire v$G17_8498_out0;
wire v$G17_8499_out0;
wire v$G17_8500_out0;
wire v$G17_8501_out0;
wire v$G17_8502_out0;
wire v$G17_8503_out0;
wire v$G17_8504_out0;
wire v$G17_8505_out0;
wire v$G17_8506_out0;
wire v$G17_8507_out0;
wire v$G17_8508_out0;
wire v$G17_8509_out0;
wire v$G17_8510_out0;
wire v$G17_9176_out0;
wire v$G17_9177_out0;
wire v$G17_9229_out0;
wire v$G17_9230_out0;
wire v$G17_9714_out0;
wire v$G17_9715_out0;
wire v$G17_9716_out0;
wire v$G17_9717_out0;
wire v$G17_9718_out0;
wire v$G17_9719_out0;
wire v$G18_10707_out0;
wire v$G18_10708_out0;
wire v$G18_11539_out0;
wire v$G18_11540_out0;
wire v$G18_13508_out0;
wire v$G18_13509_out0;
wire v$G18_13510_out0;
wire v$G18_13511_out0;
wire v$G18_13512_out0;
wire v$G18_13513_out0;
wire v$G18_14086_out0;
wire v$G18_14087_out0;
wire v$G18_14176_out0;
wire v$G18_14177_out0;
wire v$G18_18705_out0;
wire v$G18_18706_out0;
wire v$G18_3199_out0;
wire v$G18_3200_out0;
wire v$G18_3607_out0;
wire v$G18_3608_out0;
wire v$G18_5188_out0;
wire v$G18_5189_out0;
wire v$G18_5190_out0;
wire v$G18_5191_out0;
wire v$G18_5192_out0;
wire v$G18_5193_out0;
wire v$G18_5194_out0;
wire v$G18_5195_out0;
wire v$G18_5196_out0;
wire v$G18_5197_out0;
wire v$G18_5198_out0;
wire v$G18_5199_out0;
wire v$G18_5200_out0;
wire v$G18_5201_out0;
wire v$G18_5202_out0;
wire v$G18_5203_out0;
wire v$G18_5204_out0;
wire v$G18_5205_out0;
wire v$G18_5206_out0;
wire v$G18_5207_out0;
wire v$G18_5208_out0;
wire v$G18_5209_out0;
wire v$G18_5210_out0;
wire v$G18_5211_out0;
wire v$G18_8726_out0;
wire v$G18_8727_out0;
wire v$G19_10699_out0;
wire v$G19_10700_out0;
wire v$G19_10701_out0;
wire v$G19_10702_out0;
wire v$G19_14605_out0;
wire v$G19_14606_out0;
wire v$G19_16478_out0;
wire v$G19_16479_out0;
wire v$G19_16556_out0;
wire v$G19_16557_out0;
wire v$G19_16657_out0;
wire v$G19_16658_out0;
wire v$G19_17314_out0;
wire v$G19_17315_out0;
wire v$G19_2044_out0;
wire v$G19_2045_out0;
wire v$G19_2046_out0;
wire v$G19_2047_out0;
wire v$G19_2048_out0;
wire v$G19_2049_out0;
wire v$G19_2605_out0;
wire v$G19_2606_out0;
wire v$G19_3050_out0;
wire v$G19_3051_out0;
wire v$G19_352_out0;
wire v$G19_353_out0;
wire v$G19_8570_out0;
wire v$G19_8571_out0;
wire v$G1_10773_out0;
wire v$G1_10774_out0;
wire v$G1_12690_out0;
wire v$G1_12691_out0;
wire v$G1_12789_out0;
wire v$G1_12790_out0;
wire v$G1_12902_out0;
wire v$G1_12903_out0;
wire v$G1_12904_out0;
wire v$G1_12905_out0;
wire v$G1_12906_out0;
wire v$G1_12907_out0;
wire v$G1_12908_out0;
wire v$G1_12909_out0;
wire v$G1_12910_out0;
wire v$G1_12911_out0;
wire v$G1_12912_out0;
wire v$G1_12913_out0;
wire v$G1_12914_out0;
wire v$G1_12915_out0;
wire v$G1_12916_out0;
wire v$G1_12917_out0;
wire v$G1_12918_out0;
wire v$G1_12919_out0;
wire v$G1_12920_out0;
wire v$G1_12921_out0;
wire v$G1_12922_out0;
wire v$G1_12923_out0;
wire v$G1_12924_out0;
wire v$G1_12925_out0;
wire v$G1_12926_out0;
wire v$G1_12927_out0;
wire v$G1_12928_out0;
wire v$G1_12929_out0;
wire v$G1_12930_out0;
wire v$G1_12931_out0;
wire v$G1_12932_out0;
wire v$G1_12933_out0;
wire v$G1_12934_out0;
wire v$G1_12935_out0;
wire v$G1_12936_out0;
wire v$G1_12937_out0;
wire v$G1_12938_out0;
wire v$G1_12939_out0;
wire v$G1_12940_out0;
wire v$G1_12941_out0;
wire v$G1_12942_out0;
wire v$G1_12943_out0;
wire v$G1_12944_out0;
wire v$G1_12945_out0;
wire v$G1_12946_out0;
wire v$G1_12947_out0;
wire v$G1_12948_out0;
wire v$G1_12949_out0;
wire v$G1_12950_out0;
wire v$G1_12951_out0;
wire v$G1_12952_out0;
wire v$G1_12953_out0;
wire v$G1_12954_out0;
wire v$G1_12955_out0;
wire v$G1_12956_out0;
wire v$G1_12957_out0;
wire v$G1_12958_out0;
wire v$G1_12959_out0;
wire v$G1_12960_out0;
wire v$G1_12961_out0;
wire v$G1_12962_out0;
wire v$G1_12963_out0;
wire v$G1_12964_out0;
wire v$G1_12965_out0;
wire v$G1_12966_out0;
wire v$G1_12967_out0;
wire v$G1_12968_out0;
wire v$G1_12969_out0;
wire v$G1_12970_out0;
wire v$G1_12971_out0;
wire v$G1_12972_out0;
wire v$G1_12973_out0;
wire v$G1_12974_out0;
wire v$G1_12975_out0;
wire v$G1_12976_out0;
wire v$G1_12977_out0;
wire v$G1_12978_out0;
wire v$G1_12979_out0;
wire v$G1_12980_out0;
wire v$G1_12981_out0;
wire v$G1_12982_out0;
wire v$G1_12983_out0;
wire v$G1_12984_out0;
wire v$G1_12985_out0;
wire v$G1_12986_out0;
wire v$G1_12987_out0;
wire v$G1_12988_out0;
wire v$G1_12989_out0;
wire v$G1_12990_out0;
wire v$G1_12991_out0;
wire v$G1_12992_out0;
wire v$G1_12993_out0;
wire v$G1_12994_out0;
wire v$G1_12995_out0;
wire v$G1_12996_out0;
wire v$G1_12997_out0;
wire v$G1_12998_out0;
wire v$G1_12999_out0;
wire v$G1_13000_out0;
wire v$G1_13001_out0;
wire v$G1_13002_out0;
wire v$G1_13003_out0;
wire v$G1_13004_out0;
wire v$G1_13005_out0;
wire v$G1_13006_out0;
wire v$G1_13007_out0;
wire v$G1_13008_out0;
wire v$G1_13009_out0;
wire v$G1_13010_out0;
wire v$G1_13011_out0;
wire v$G1_13012_out0;
wire v$G1_13013_out0;
wire v$G1_13014_out0;
wire v$G1_13015_out0;
wire v$G1_13016_out0;
wire v$G1_13017_out0;
wire v$G1_13018_out0;
wire v$G1_13019_out0;
wire v$G1_13020_out0;
wire v$G1_13021_out0;
wire v$G1_13022_out0;
wire v$G1_13023_out0;
wire v$G1_13024_out0;
wire v$G1_13025_out0;
wire v$G1_13026_out0;
wire v$G1_13027_out0;
wire v$G1_13028_out0;
wire v$G1_13029_out0;
wire v$G1_13030_out0;
wire v$G1_13031_out0;
wire v$G1_13032_out0;
wire v$G1_13033_out0;
wire v$G1_13034_out0;
wire v$G1_13035_out0;
wire v$G1_13036_out0;
wire v$G1_13037_out0;
wire v$G1_13038_out0;
wire v$G1_13039_out0;
wire v$G1_13040_out0;
wire v$G1_13041_out0;
wire v$G1_13042_out0;
wire v$G1_13043_out0;
wire v$G1_13044_out0;
wire v$G1_13045_out0;
wire v$G1_1343_out0;
wire v$G1_1344_out0;
wire v$G1_13554_out0;
wire v$G1_13555_out0;
wire v$G1_13556_out0;
wire v$G1_13557_out0;
wire v$G1_13558_out0;
wire v$G1_13559_out0;
wire v$G1_13560_out0;
wire v$G1_13725_out0;
wire v$G1_13726_out0;
wire v$G1_13767_out0;
wire v$G1_13768_out0;
wire v$G1_13769_out0;
wire v$G1_13770_out0;
wire v$G1_1403_out0;
wire v$G1_1404_out0;
wire v$G1_14123_out0;
wire v$G1_14124_out0;
wire v$G1_15015_out0;
wire v$G1_15078_out0;
wire v$G1_15079_out0;
wire v$G1_15191_out0;
wire v$G1_15192_out0;
wire v$G1_15193_out0;
wire v$G1_15194_out0;
wire v$G1_15195_out0;
wire v$G1_15196_out0;
wire v$G1_15197_out0;
wire v$G1_15198_out0;
wire v$G1_15199_out0;
wire v$G1_15200_out0;
wire v$G1_15752_out0;
wire v$G1_15753_out0;
wire v$G1_15877_out0;
wire v$G1_15878_out0;
wire v$G1_16179_out0;
wire v$G1_16180_out0;
wire v$G1_16383_out0;
wire v$G1_16384_out0;
wire v$G1_16643_out0;
wire v$G1_16644_out0;
wire v$G1_16645_out0;
wire v$G1_16646_out0;
wire v$G1_16647_out0;
wire v$G1_16648_out0;
wire v$G1_16649_out0;
wire v$G1_16650_out0;
wire v$G1_166_out0;
wire v$G1_16754_out0;
wire v$G1_16755_out0;
wire v$G1_16756_out0;
wire v$G1_16757_out0;
wire v$G1_167_out0;
wire v$G1_17020_out0;
wire v$G1_17021_out0;
wire v$G1_17122_out0;
wire v$G1_17123_out0;
wire v$G1_1750_out0;
wire v$G1_1751_out0;
wire v$G1_17610_out0;
wire v$G1_17611_out0;
wire v$G1_18090_out0;
wire v$G1_18091_out0;
wire v$G1_18092_out0;
wire v$G1_18093_out0;
wire v$G1_18498_out0;
wire v$G1_18499_out0;
wire v$G1_19257_out0;
wire v$G1_19258_out0;
wire v$G1_2078_out0;
wire v$G1_2079_out0;
wire v$G1_34_out0;
wire v$G1_35_out0;
wire v$G1_4372_out0;
wire v$G1_4373_out0;
wire v$G1_5269_out0;
wire v$G1_5270_out0;
wire v$G1_5271_out0;
wire v$G1_5272_out0;
wire v$G1_5273_out0;
wire v$G1_5274_out0;
wire v$G1_5662_out0;
wire v$G1_5663_out0;
wire v$G1_5763_out0;
wire v$G1_5764_out0;
wire v$G1_5765_out0;
wire v$G1_5766_out0;
wire v$G1_5767_out0;
wire v$G1_5768_out0;
wire v$G1_5769_out0;
wire v$G1_5770_out0;
wire v$G1_5771_out0;
wire v$G1_5772_out0;
wire v$G1_5773_out0;
wire v$G1_5774_out0;
wire v$G1_5775_out0;
wire v$G1_5776_out0;
wire v$G1_5777_out0;
wire v$G1_5778_out0;
wire v$G1_5779_out0;
wire v$G1_5780_out0;
wire v$G1_5781_out0;
wire v$G1_5782_out0;
wire v$G1_5783_out0;
wire v$G1_5784_out0;
wire v$G1_5785_out0;
wire v$G1_5786_out0;
wire v$G1_5787_out0;
wire v$G1_5788_out0;
wire v$G1_5789_out0;
wire v$G1_5790_out0;
wire v$G1_5791_out0;
wire v$G1_5792_out0;
wire v$G1_5793_out0;
wire v$G1_5794_out0;
wire v$G1_5795_out0;
wire v$G1_5796_out0;
wire v$G1_5797_out0;
wire v$G1_5798_out0;
wire v$G1_5799_out0;
wire v$G1_5800_out0;
wire v$G1_5801_out0;
wire v$G1_5802_out0;
wire v$G1_5803_out0;
wire v$G1_5804_out0;
wire v$G1_5805_out0;
wire v$G1_5806_out0;
wire v$G1_5807_out0;
wire v$G1_5808_out0;
wire v$G1_5809_out0;
wire v$G1_5810_out0;
wire v$G1_5811_out0;
wire v$G1_5812_out0;
wire v$G1_5813_out0;
wire v$G1_5814_out0;
wire v$G1_5815_out0;
wire v$G1_5816_out0;
wire v$G1_5817_out0;
wire v$G1_5818_out0;
wire v$G1_5819_out0;
wire v$G1_5820_out0;
wire v$G1_5821_out0;
wire v$G1_5822_out0;
wire v$G1_5823_out0;
wire v$G1_5824_out0;
wire v$G1_5825_out0;
wire v$G1_5826_out0;
wire v$G1_5827_out0;
wire v$G1_5828_out0;
wire v$G1_5829_out0;
wire v$G1_5830_out0;
wire v$G1_5831_out0;
wire v$G1_5832_out0;
wire v$G1_5833_out0;
wire v$G1_5834_out0;
wire v$G1_5835_out0;
wire v$G1_5836_out0;
wire v$G1_5837_out0;
wire v$G1_5838_out0;
wire v$G1_5839_out0;
wire v$G1_5840_out0;
wire v$G1_5841_out0;
wire v$G1_5842_out0;
wire v$G1_5843_out0;
wire v$G1_5844_out0;
wire v$G1_5845_out0;
wire v$G1_5846_out0;
wire v$G1_5847_out0;
wire v$G1_5848_out0;
wire v$G1_5849_out0;
wire v$G1_5850_out0;
wire v$G1_5851_out0;
wire v$G1_5852_out0;
wire v$G1_5853_out0;
wire v$G1_5854_out0;
wire v$G1_5855_out0;
wire v$G1_5856_out0;
wire v$G1_5857_out0;
wire v$G1_5858_out0;
wire v$G1_5859_out0;
wire v$G1_5860_out0;
wire v$G1_5861_out0;
wire v$G1_5862_out0;
wire v$G1_5863_out0;
wire v$G1_5864_out0;
wire v$G1_5865_out0;
wire v$G1_5866_out0;
wire v$G1_5867_out0;
wire v$G1_5868_out0;
wire v$G1_5869_out0;
wire v$G1_5870_out0;
wire v$G1_5871_out0;
wire v$G1_5872_out0;
wire v$G1_5873_out0;
wire v$G1_5874_out0;
wire v$G1_5875_out0;
wire v$G1_5876_out0;
wire v$G1_5877_out0;
wire v$G1_5878_out0;
wire v$G1_5879_out0;
wire v$G1_5880_out0;
wire v$G1_5881_out0;
wire v$G1_5882_out0;
wire v$G1_5883_out0;
wire v$G1_5884_out0;
wire v$G1_5885_out0;
wire v$G1_5886_out0;
wire v$G1_5887_out0;
wire v$G1_5888_out0;
wire v$G1_5889_out0;
wire v$G1_5890_out0;
wire v$G1_5891_out0;
wire v$G1_5892_out0;
wire v$G1_5893_out0;
wire v$G1_5894_out0;
wire v$G1_5895_out0;
wire v$G1_5896_out0;
wire v$G1_5897_out0;
wire v$G1_5898_out0;
wire v$G1_5899_out0;
wire v$G1_5900_out0;
wire v$G1_5901_out0;
wire v$G1_5902_out0;
wire v$G1_5903_out0;
wire v$G1_5904_out0;
wire v$G1_5905_out0;
wire v$G1_5906_out0;
wire v$G1_5907_out0;
wire v$G1_5908_out0;
wire v$G1_5909_out0;
wire v$G1_5910_out0;
wire v$G1_5911_out0;
wire v$G1_5912_out0;
wire v$G1_5913_out0;
wire v$G1_5914_out0;
wire v$G1_5915_out0;
wire v$G1_5916_out0;
wire v$G1_5917_out0;
wire v$G1_5918_out0;
wire v$G1_5919_out0;
wire v$G1_5920_out0;
wire v$G1_5921_out0;
wire v$G1_5922_out0;
wire v$G1_5923_out0;
wire v$G1_5924_out0;
wire v$G1_5925_out0;
wire v$G1_5926_out0;
wire v$G1_5927_out0;
wire v$G1_5928_out0;
wire v$G1_5929_out0;
wire v$G1_5930_out0;
wire v$G1_5931_out0;
wire v$G1_5932_out0;
wire v$G1_5933_out0;
wire v$G1_5934_out0;
wire v$G1_5935_out0;
wire v$G1_5936_out0;
wire v$G1_5937_out0;
wire v$G1_5938_out0;
wire v$G1_5939_out0;
wire v$G1_5940_out0;
wire v$G1_5941_out0;
wire v$G1_5942_out0;
wire v$G1_5943_out0;
wire v$G1_5944_out0;
wire v$G1_5945_out0;
wire v$G1_5946_out0;
wire v$G1_5947_out0;
wire v$G1_5948_out0;
wire v$G1_5949_out0;
wire v$G1_5950_out0;
wire v$G1_5951_out0;
wire v$G1_5952_out0;
wire v$G1_5953_out0;
wire v$G1_5954_out0;
wire v$G1_5955_out0;
wire v$G1_5956_out0;
wire v$G1_5957_out0;
wire v$G1_5958_out0;
wire v$G1_5959_out0;
wire v$G1_5960_out0;
wire v$G1_5961_out0;
wire v$G1_5962_out0;
wire v$G1_5963_out0;
wire v$G1_5964_out0;
wire v$G1_5965_out0;
wire v$G1_5966_out0;
wire v$G1_5967_out0;
wire v$G1_5968_out0;
wire v$G1_5969_out0;
wire v$G1_5970_out0;
wire v$G1_5971_out0;
wire v$G1_5972_out0;
wire v$G1_5973_out0;
wire v$G1_5974_out0;
wire v$G1_5975_out0;
wire v$G1_5976_out0;
wire v$G1_5977_out0;
wire v$G1_5978_out0;
wire v$G1_5979_out0;
wire v$G1_5980_out0;
wire v$G1_5981_out0;
wire v$G1_5982_out0;
wire v$G1_5983_out0;
wire v$G1_5984_out0;
wire v$G1_5985_out0;
wire v$G1_5986_out0;
wire v$G1_5987_out0;
wire v$G1_5988_out0;
wire v$G1_5989_out0;
wire v$G1_5990_out0;
wire v$G1_5991_out0;
wire v$G1_5992_out0;
wire v$G1_5993_out0;
wire v$G1_5994_out0;
wire v$G1_5995_out0;
wire v$G1_5996_out0;
wire v$G1_5997_out0;
wire v$G1_5998_out0;
wire v$G1_5999_out0;
wire v$G1_6000_out0;
wire v$G1_6001_out0;
wire v$G1_6002_out0;
wire v$G1_6003_out0;
wire v$G1_6004_out0;
wire v$G1_6005_out0;
wire v$G1_6006_out0;
wire v$G1_6007_out0;
wire v$G1_6008_out0;
wire v$G1_7537_out0;
wire v$G1_7538_out0;
wire v$G1_7643_out0;
wire v$G1_7644_out0;
wire v$G1_7651_out0;
wire v$G1_9137_out0;
wire v$G1_9138_out0;
wire v$G1_9139_out0;
wire v$G1_9140_out0;
wire v$G1_9759_out0;
wire v$G1_9760_out0;
wire v$G1_9761_out0;
wire v$G1_9762_out0;
wire v$G1_9763_out0;
wire v$G1_9764_out0;
wire v$G1_9765_out0;
wire v$G1_9766_out0;
wire v$G20_10303_out0;
wire v$G20_10304_out0;
wire v$G20_10305_out0;
wire v$G20_10306_out0;
wire v$G20_10307_out0;
wire v$G20_10308_out0;
wire v$G20_10309_out0;
wire v$G20_10310_out0;
wire v$G20_10311_out0;
wire v$G20_10312_out0;
wire v$G20_10313_out0;
wire v$G20_10314_out0;
wire v$G20_10315_out0;
wire v$G20_10316_out0;
wire v$G20_10317_out0;
wire v$G20_10318_out0;
wire v$G20_10319_out0;
wire v$G20_10320_out0;
wire v$G20_10321_out0;
wire v$G20_10322_out0;
wire v$G20_10323_out0;
wire v$G20_10324_out0;
wire v$G20_10325_out0;
wire v$G20_10326_out0;
wire v$G20_12278_out0;
wire v$G20_12279_out0;
wire v$G20_12774_out0;
wire v$G20_12775_out0;
wire v$G20_12859_out0;
wire v$G20_12860_out0;
wire v$G20_13310_out0;
wire v$G20_13311_out0;
wire v$G20_16542_out0;
wire v$G20_16543_out0;
wire v$G20_18885_out0;
wire v$G20_18886_out0;
wire v$G20_2788_out0;
wire v$G20_2789_out0;
wire v$G20_5691_out0;
wire v$G20_5692_out0;
wire v$G20_7717_out0;
wire v$G20_7718_out0;
wire v$G20_8533_out0;
wire v$G20_8534_out0;
wire v$G20_8535_out0;
wire v$G20_8536_out0;
wire v$G20_8537_out0;
wire v$G20_8538_out0;
wire v$G21_12447_out0;
wire v$G21_12448_out0;
wire v$G21_14626_out0;
wire v$G21_14627_out0;
wire v$G21_14628_out0;
wire v$G21_14629_out0;
wire v$G21_14630_out0;
wire v$G21_14631_out0;
wire v$G21_14847_out0;
wire v$G21_14848_out0;
wire v$G21_15317_out0;
wire v$G21_15318_out0;
wire v$G21_15897_out0;
wire v$G21_15898_out0;
wire v$G21_16426_out0;
wire v$G21_16427_out0;
wire v$G21_18276_out0;
wire v$G21_18277_out0;
wire v$G21_19292_out0;
wire v$G21_19293_out0;
wire v$G21_3722_out0;
wire v$G21_3723_out0;
wire v$G21_3724_out0;
wire v$G21_3725_out0;
wire v$G21_3726_out0;
wire v$G21_3727_out0;
wire v$G21_3728_out0;
wire v$G21_3729_out0;
wire v$G21_3730_out0;
wire v$G21_3731_out0;
wire v$G21_3732_out0;
wire v$G21_3733_out0;
wire v$G21_3734_out0;
wire v$G21_3735_out0;
wire v$G21_3736_out0;
wire v$G21_3737_out0;
wire v$G21_3738_out0;
wire v$G21_3739_out0;
wire v$G21_3740_out0;
wire v$G21_3741_out0;
wire v$G21_3742_out0;
wire v$G21_3743_out0;
wire v$G21_3744_out0;
wire v$G21_3745_out0;
wire v$G21_7321_out0;
wire v$G21_7322_out0;
wire v$G21_7802_out0;
wire v$G21_7803_out0;
wire v$G22_13104_out0;
wire v$G22_13105_out0;
wire v$G22_13106_out0;
wire v$G22_13107_out0;
wire v$G22_13108_out0;
wire v$G22_13109_out0;
wire v$G22_13912_out0;
wire v$G22_13913_out0;
wire v$G22_13914_out0;
wire v$G22_13915_out0;
wire v$G22_13916_out0;
wire v$G22_13917_out0;
wire v$G22_13918_out0;
wire v$G22_13919_out0;
wire v$G22_13920_out0;
wire v$G22_13921_out0;
wire v$G22_13922_out0;
wire v$G22_13923_out0;
wire v$G22_13924_out0;
wire v$G22_13925_out0;
wire v$G22_13926_out0;
wire v$G22_13927_out0;
wire v$G22_13928_out0;
wire v$G22_13929_out0;
wire v$G22_13930_out0;
wire v$G22_13931_out0;
wire v$G22_13932_out0;
wire v$G22_13933_out0;
wire v$G22_13934_out0;
wire v$G22_13935_out0;
wire v$G22_15929_out0;
wire v$G22_15930_out0;
wire v$G22_16224_out0;
wire v$G22_16225_out0;
wire v$G22_16456_out0;
wire v$G22_16457_out0;
wire v$G22_4474_out0;
wire v$G22_4475_out0;
wire v$G22_5098_out0;
wire v$G22_5099_out0;
wire v$G22_5701_out0;
wire v$G22_5702_out0;
wire v$G22_7584_out0;
wire v$G22_7585_out0;
wire v$G23_12740_out0;
wire v$G23_12741_out0;
wire v$G23_12742_out0;
wire v$G23_12743_out0;
wire v$G23_12744_out0;
wire v$G23_12745_out0;
wire v$G23_12746_out0;
wire v$G23_12747_out0;
wire v$G23_12748_out0;
wire v$G23_12749_out0;
wire v$G23_12750_out0;
wire v$G23_12751_out0;
wire v$G23_12752_out0;
wire v$G23_12753_out0;
wire v$G23_12754_out0;
wire v$G23_12755_out0;
wire v$G23_12756_out0;
wire v$G23_12757_out0;
wire v$G23_12758_out0;
wire v$G23_12759_out0;
wire v$G23_12760_out0;
wire v$G23_12761_out0;
wire v$G23_12762_out0;
wire v$G23_12763_out0;
wire v$G23_14691_out0;
wire v$G23_14692_out0;
wire v$G23_14920_out0;
wire v$G23_14921_out0;
wire v$G23_14922_out0;
wire v$G23_14923_out0;
wire v$G23_14924_out0;
wire v$G23_14925_out0;
wire v$G23_16554_out0;
wire v$G23_16555_out0;
wire v$G23_17391_out0;
wire v$G23_17392_out0;
wire v$G23_18289_out0;
wire v$G23_18290_out0;
wire v$G23_19263_out0;
wire v$G23_19264_out0;
wire v$G23_2483_out0;
wire v$G23_2484_out0;
wire v$G23_4550_out0;
wire v$G23_4551_out0;
wire v$G23_7274_out0;
wire v$G23_7275_out0;
wire v$G23_9729_out0;
wire v$G23_9730_out0;
wire v$G23_9982_out0;
wire v$G23_9983_out0;
wire v$G24_10000_out0;
wire v$G24_10001_out0;
wire v$G24_10805_out0;
wire v$G24_10806_out0;
wire v$G24_12651_out0;
wire v$G24_12652_out0;
wire v$G24_14443_out0;
wire v$G24_14444_out0;
wire v$G24_16279_out0;
wire v$G24_16280_out0;
wire v$G24_16281_out0;
wire v$G24_16282_out0;
wire v$G24_16283_out0;
wire v$G24_16284_out0;
wire v$G24_16285_out0;
wire v$G24_16286_out0;
wire v$G24_16287_out0;
wire v$G24_16288_out0;
wire v$G24_16289_out0;
wire v$G24_16290_out0;
wire v$G24_16291_out0;
wire v$G24_16292_out0;
wire v$G24_16293_out0;
wire v$G24_16294_out0;
wire v$G24_16295_out0;
wire v$G24_16296_out0;
wire v$G24_16297_out0;
wire v$G24_16298_out0;
wire v$G24_16299_out0;
wire v$G24_16300_out0;
wire v$G24_16301_out0;
wire v$G24_16302_out0;
wire v$G24_17612_out0;
wire v$G24_17613_out0;
wire v$G24_18545_out0;
wire v$G24_18546_out0;
wire v$G24_18994_out0;
wire v$G24_18995_out0;
wire v$G24_249_out0;
wire v$G24_250_out0;
wire v$G24_3609_out0;
wire v$G24_3610_out0;
wire v$G24_734_out0;
wire v$G24_735_out0;
wire v$G24_8223_out0;
wire v$G24_8224_out0;
wire v$G25_10727_out0;
wire v$G25_10728_out0;
wire v$G25_11439_out0;
wire v$G25_11440_out0;
wire v$G25_11441_out0;
wire v$G25_11442_out0;
wire v$G25_11443_out0;
wire v$G25_11444_out0;
wire v$G25_11445_out0;
wire v$G25_11446_out0;
wire v$G25_11447_out0;
wire v$G25_11448_out0;
wire v$G25_11449_out0;
wire v$G25_11450_out0;
wire v$G25_11451_out0;
wire v$G25_11452_out0;
wire v$G25_11453_out0;
wire v$G25_11454_out0;
wire v$G25_11455_out0;
wire v$G25_11456_out0;
wire v$G25_11457_out0;
wire v$G25_11458_out0;
wire v$G25_11459_out0;
wire v$G25_11460_out0;
wire v$G25_11461_out0;
wire v$G25_11462_out0;
wire v$G25_13323_out0;
wire v$G25_13324_out0;
wire v$G25_13587_out0;
wire v$G25_13588_out0;
wire v$G25_14641_out0;
wire v$G25_14642_out0;
wire v$G25_1470_out0;
wire v$G25_1471_out0;
wire v$G25_15179_out0;
wire v$G25_15180_out0;
wire v$G25_15262_out0;
wire v$G25_15263_out0;
wire v$G25_16715_out0;
wire v$G25_16716_out0;
wire v$G25_18703_out0;
wire v$G25_18704_out0;
wire v$G25_2658_out0;
wire v$G25_2659_out0;
wire v$G25_3750_out0;
wire v$G25_3751_out0;
wire v$G26_10775_out0;
wire v$G26_10776_out0;
wire v$G26_11896_out0;
wire v$G26_11897_out0;
wire v$G26_11898_out0;
wire v$G26_11899_out0;
wire v$G26_13237_out0;
wire v$G26_13238_out0;
wire v$G26_13755_out0;
wire v$G26_13756_out0;
wire v$G26_14220_out0;
wire v$G26_14221_out0;
wire v$G26_15513_out0;
wire v$G26_15514_out0;
wire v$G26_16633_out0;
wire v$G26_16634_out0;
wire v$G26_16639_out0;
wire v$G26_16640_out0;
wire v$G26_18725_out0;
wire v$G26_18726_out0;
wire v$G26_4254_out0;
wire v$G26_4255_out0;
wire v$G26_5343_out0;
wire v$G26_5344_out0;
wire v$G27_10687_out0;
wire v$G27_10688_out0;
wire v$G27_11224_out0;
wire v$G27_11225_out0;
wire v$G27_12274_out0;
wire v$G27_12275_out0;
wire v$G27_12276_out0;
wire v$G27_12277_out0;
wire v$G27_17148_out0;
wire v$G27_17149_out0;
wire v$G27_19099_out0;
wire v$G27_19100_out0;
wire v$G27_269_out0;
wire v$G27_2708_out0;
wire v$G27_2709_out0;
wire v$G27_270_out0;
wire v$G27_4064_out0;
wire v$G27_4065_out0;
wire v$G27_4989_out0;
wire v$G27_4990_out0;
wire v$G27_4991_out0;
wire v$G27_4992_out0;
wire v$G27_4993_out0;
wire v$G27_4994_out0;
wire v$G27_4995_out0;
wire v$G27_4996_out0;
wire v$G27_4997_out0;
wire v$G27_4998_out0;
wire v$G27_4999_out0;
wire v$G27_5000_out0;
wire v$G27_5001_out0;
wire v$G27_5002_out0;
wire v$G27_5003_out0;
wire v$G27_5004_out0;
wire v$G27_5005_out0;
wire v$G27_5006_out0;
wire v$G27_5007_out0;
wire v$G27_5008_out0;
wire v$G27_5009_out0;
wire v$G27_5010_out0;
wire v$G27_5011_out0;
wire v$G27_5012_out0;
wire v$G28_11298_out0;
wire v$G28_11299_out0;
wire v$G28_12513_out0;
wire v$G28_12514_out0;
wire v$G28_13591_out0;
wire v$G28_13592_out0;
wire v$G28_13593_out0;
wire v$G28_13594_out0;
wire v$G28_13595_out0;
wire v$G28_13596_out0;
wire v$G28_13597_out0;
wire v$G28_13598_out0;
wire v$G28_13599_out0;
wire v$G28_13600_out0;
wire v$G28_13601_out0;
wire v$G28_13602_out0;
wire v$G28_13603_out0;
wire v$G28_13604_out0;
wire v$G28_13605_out0;
wire v$G28_13606_out0;
wire v$G28_13607_out0;
wire v$G28_13608_out0;
wire v$G28_13609_out0;
wire v$G28_13610_out0;
wire v$G28_13611_out0;
wire v$G28_13612_out0;
wire v$G28_13613_out0;
wire v$G28_13614_out0;
wire v$G28_14373_out0;
wire v$G28_14374_out0;
wire v$G28_15272_out0;
wire v$G28_15273_out0;
wire v$G28_15972_out0;
wire v$G28_15973_out0;
wire v$G28_16226_out0;
wire v$G28_16227_out0;
wire v$G28_19161_out0;
wire v$G28_19162_out0;
wire v$G28_3387_out0;
wire v$G28_3388_out0;
wire v$G28_3947_out0;
wire v$G28_3948_out0;
wire v$G28_9040_out0;
wire v$G28_9041_out0;
wire v$G29_10753_out0;
wire v$G29_10754_out0;
wire v$G29_10755_out0;
wire v$G29_10756_out0;
wire v$G29_11326_out0;
wire v$G29_11327_out0;
wire v$G29_14601_out0;
wire v$G29_14602_out0;
wire v$G29_16375_out0;
wire v$G29_16376_out0;
wire v$G29_3814_out0;
wire v$G29_3815_out0;
wire v$G29_5727_out0;
wire v$G29_5728_out0;
wire v$G29_744_out0;
wire v$G29_745_out0;
wire v$G29_7784_out0;
wire v$G29_7785_out0;
wire v$G29_8174_out0;
wire v$G29_8175_out0;
wire v$G2_10851_out0;
wire v$G2_10852_out0;
wire v$G2_10853_out0;
wire v$G2_10854_out0;
wire v$G2_12265_out0;
wire v$G2_12476_out0;
wire v$G2_12477_out0;
wire v$G2_12478_out0;
wire v$G2_12479_out0;
wire v$G2_13475_out0;
wire v$G2_13476_out0;
wire v$G2_13477_out0;
wire v$G2_13478_out0;
wire v$G2_13479_out0;
wire v$G2_13480_out0;
wire v$G2_13481_out0;
wire v$G2_13482_out0;
wire v$G2_14274_out0;
wire v$G2_14275_out0;
wire v$G2_1447_out0;
wire v$G2_1448_out0;
wire v$G2_15098_out0;
wire v$G2_15099_out0;
wire v$G2_15651_out0;
wire v$G2_15652_out0;
wire v$G2_15653_out0;
wire v$G2_15654_out0;
wire v$G2_15655_out0;
wire v$G2_15656_out0;
wire v$G2_15657_out0;
wire v$G2_15658_out0;
wire v$G2_15659_out0;
wire v$G2_15660_out0;
wire v$G2_15661_out0;
wire v$G2_15662_out0;
wire v$G2_16133_out0;
wire v$G2_16134_out0;
wire v$G2_16361_out0;
wire v$G2_16362_out0;
wire v$G2_16466_out0;
wire v$G2_16467_out0;
wire v$G2_16568_out0;
wire v$G2_16569_out0;
wire v$G2_16570_out0;
wire v$G2_16571_out0;
wire v$G2_16572_out0;
wire v$G2_16573_out0;
wire v$G2_17128_out0;
wire v$G2_17129_out0;
wire v$G2_17660_out0;
wire v$G2_17661_out0;
wire v$G2_18054_out0;
wire v$G2_18055_out0;
wire v$G2_18056_out0;
wire v$G2_18057_out0;
wire v$G2_18058_out0;
wire v$G2_18059_out0;
wire v$G2_18060_out0;
wire v$G2_18061_out0;
wire v$G2_18263_out0;
wire v$G2_18264_out0;
wire v$G2_18840_out0;
wire v$G2_18841_out0;
wire v$G2_18842_out0;
wire v$G2_18843_out0;
wire v$G2_19037_out0;
wire v$G2_19038_out0;
wire v$G2_19310_out0;
wire v$G2_19311_out0;
wire v$G2_2058_out0;
wire v$G2_2059_out0;
wire v$G2_2620_out0;
wire v$G2_2621_out0;
wire v$G2_3905_out0;
wire v$G2_3906_out0;
wire v$G2_4246_out0;
wire v$G2_4247_out0;
wire v$G2_5263_out0;
wire v$G2_5264_out0;
wire v$G2_5471_out0;
wire v$G2_5472_out0;
wire v$G2_5478_out0;
wire v$G2_5479_out0;
wire v$G2_5480_out0;
wire v$G2_5481_out0;
wire v$G2_5482_out0;
wire v$G2_5483_out0;
wire v$G2_5484_out0;
wire v$G2_5485_out0;
wire v$G2_5486_out0;
wire v$G2_5487_out0;
wire v$G2_5488_out0;
wire v$G2_5489_out0;
wire v$G2_5490_out0;
wire v$G2_5491_out0;
wire v$G2_5492_out0;
wire v$G2_5493_out0;
wire v$G2_5494_out0;
wire v$G2_5495_out0;
wire v$G2_5496_out0;
wire v$G2_5497_out0;
wire v$G2_5498_out0;
wire v$G2_5499_out0;
wire v$G2_5500_out0;
wire v$G2_5501_out0;
wire v$G2_5502_out0;
wire v$G2_5503_out0;
wire v$G2_5504_out0;
wire v$G2_5505_out0;
wire v$G2_5506_out0;
wire v$G2_5507_out0;
wire v$G2_5508_out0;
wire v$G2_5509_out0;
wire v$G2_5510_out0;
wire v$G2_5511_out0;
wire v$G2_5512_out0;
wire v$G2_5513_out0;
wire v$G2_5514_out0;
wire v$G2_5515_out0;
wire v$G2_5516_out0;
wire v$G2_5517_out0;
wire v$G2_5518_out0;
wire v$G2_5519_out0;
wire v$G2_5520_out0;
wire v$G2_5521_out0;
wire v$G2_5522_out0;
wire v$G2_5523_out0;
wire v$G2_5524_out0;
wire v$G2_5525_out0;
wire v$G2_5526_out0;
wire v$G2_5527_out0;
wire v$G2_5528_out0;
wire v$G2_5529_out0;
wire v$G2_5530_out0;
wire v$G2_5531_out0;
wire v$G2_5532_out0;
wire v$G2_5533_out0;
wire v$G2_5534_out0;
wire v$G2_5535_out0;
wire v$G2_5536_out0;
wire v$G2_5537_out0;
wire v$G2_5538_out0;
wire v$G2_5539_out0;
wire v$G2_5540_out0;
wire v$G2_5541_out0;
wire v$G2_5542_out0;
wire v$G2_5543_out0;
wire v$G2_5544_out0;
wire v$G2_5545_out0;
wire v$G2_5546_out0;
wire v$G2_5547_out0;
wire v$G2_5548_out0;
wire v$G2_5549_out0;
wire v$G2_5550_out0;
wire v$G2_5551_out0;
wire v$G2_5552_out0;
wire v$G2_5553_out0;
wire v$G2_5554_out0;
wire v$G2_5555_out0;
wire v$G2_5556_out0;
wire v$G2_5557_out0;
wire v$G2_5558_out0;
wire v$G2_5559_out0;
wire v$G2_5560_out0;
wire v$G2_5561_out0;
wire v$G2_5562_out0;
wire v$G2_5563_out0;
wire v$G2_5564_out0;
wire v$G2_5565_out0;
wire v$G2_5566_out0;
wire v$G2_5567_out0;
wire v$G2_5568_out0;
wire v$G2_5569_out0;
wire v$G2_5570_out0;
wire v$G2_5571_out0;
wire v$G2_5572_out0;
wire v$G2_5573_out0;
wire v$G2_5574_out0;
wire v$G2_5575_out0;
wire v$G2_5576_out0;
wire v$G2_5577_out0;
wire v$G2_5578_out0;
wire v$G2_5579_out0;
wire v$G2_5580_out0;
wire v$G2_5581_out0;
wire v$G2_5582_out0;
wire v$G2_5583_out0;
wire v$G2_5584_out0;
wire v$G2_5585_out0;
wire v$G2_5586_out0;
wire v$G2_5587_out0;
wire v$G2_5588_out0;
wire v$G2_5589_out0;
wire v$G2_5590_out0;
wire v$G2_5591_out0;
wire v$G2_5592_out0;
wire v$G2_5593_out0;
wire v$G2_5594_out0;
wire v$G2_5595_out0;
wire v$G2_5596_out0;
wire v$G2_5597_out0;
wire v$G2_5598_out0;
wire v$G2_5599_out0;
wire v$G2_5600_out0;
wire v$G2_5601_out0;
wire v$G2_5602_out0;
wire v$G2_5603_out0;
wire v$G2_5604_out0;
wire v$G2_5605_out0;
wire v$G2_5606_out0;
wire v$G2_5607_out0;
wire v$G2_5608_out0;
wire v$G2_5609_out0;
wire v$G2_5610_out0;
wire v$G2_5611_out0;
wire v$G2_5612_out0;
wire v$G2_5613_out0;
wire v$G2_5614_out0;
wire v$G2_5615_out0;
wire v$G2_5616_out0;
wire v$G2_5617_out0;
wire v$G2_5618_out0;
wire v$G2_5619_out0;
wire v$G2_5620_out0;
wire v$G2_5621_out0;
wire v$G2_5670_out0;
wire v$G2_5671_out0;
wire v$G2_66_out0;
wire v$G2_67_out0;
wire v$G2_7886_out0;
wire v$G2_7899_out0;
wire v$G2_7900_out0;
wire v$G2_7901_out0;
wire v$G2_7902_out0;
wire v$G2_7903_out0;
wire v$G2_7904_out0;
wire v$G2_7905_out0;
wire v$G2_8098_out0;
wire v$G2_8099_out0;
wire v$G2_8434_out0;
wire v$G2_8647_out0;
wire v$G2_8648_out0;
wire v$G2_9406_out0;
wire v$G2_9407_out0;
wire v$G30_16506_out0;
wire v$G30_16507_out0;
wire v$G30_1877_out0;
wire v$G30_1878_out0;
wire v$G30_19215_out0;
wire v$G30_19216_out0;
wire v$G30_1930_out0;
wire v$G30_1931_out0;
wire v$G30_1932_out0;
wire v$G30_1933_out0;
wire v$G30_1934_out0;
wire v$G30_1935_out0;
wire v$G30_1936_out0;
wire v$G30_1937_out0;
wire v$G30_1938_out0;
wire v$G30_1939_out0;
wire v$G30_1940_out0;
wire v$G30_1941_out0;
wire v$G30_1942_out0;
wire v$G30_1943_out0;
wire v$G30_1944_out0;
wire v$G30_1945_out0;
wire v$G30_1946_out0;
wire v$G30_1947_out0;
wire v$G30_1948_out0;
wire v$G30_1949_out0;
wire v$G30_1950_out0;
wire v$G30_1951_out0;
wire v$G30_1952_out0;
wire v$G30_1953_out0;
wire v$G30_2660_out0;
wire v$G30_2661_out0;
wire v$G30_3945_out0;
wire v$G30_3946_out0;
wire v$G30_5138_out0;
wire v$G30_5139_out0;
wire v$G31_10014_out0;
wire v$G31_10015_out0;
wire v$G31_11288_out0;
wire v$G31_11289_out0;
wire v$G31_16097_out0;
wire v$G31_16098_out0;
wire v$G31_16099_out0;
wire v$G31_16100_out0;
wire v$G31_16101_out0;
wire v$G31_16102_out0;
wire v$G31_16103_out0;
wire v$G31_16104_out0;
wire v$G31_16105_out0;
wire v$G31_16106_out0;
wire v$G31_16107_out0;
wire v$G31_16108_out0;
wire v$G31_16109_out0;
wire v$G31_16110_out0;
wire v$G31_16111_out0;
wire v$G31_16112_out0;
wire v$G31_16113_out0;
wire v$G31_16114_out0;
wire v$G31_16115_out0;
wire v$G31_16116_out0;
wire v$G31_16117_out0;
wire v$G31_16118_out0;
wire v$G31_16119_out0;
wire v$G31_16120_out0;
wire v$G31_19245_out0;
wire v$G31_19246_out0;
wire v$G31_1983_out0;
wire v$G31_1984_out0;
wire v$G31_2537_out0;
wire v$G31_2538_out0;
wire v$G32_12457_out0;
wire v$G32_12458_out0;
wire v$G32_14802_out0;
wire v$G32_14803_out0;
wire v$G32_16950_out0;
wire v$G32_16951_out0;
wire v$G32_16952_out0;
wire v$G32_16953_out0;
wire v$G32_17032_out0;
wire v$G32_17033_out0;
wire v$G32_1987_out0;
wire v$G32_1988_out0;
wire v$G32_411_out0;
wire v$G32_412_out0;
wire v$G32_413_out0;
wire v$G32_414_out0;
wire v$G32_415_out0;
wire v$G32_416_out0;
wire v$G32_417_out0;
wire v$G32_418_out0;
wire v$G32_419_out0;
wire v$G32_420_out0;
wire v$G32_421_out0;
wire v$G32_422_out0;
wire v$G32_423_out0;
wire v$G32_424_out0;
wire v$G32_425_out0;
wire v$G32_426_out0;
wire v$G32_427_out0;
wire v$G32_428_out0;
wire v$G32_429_out0;
wire v$G32_430_out0;
wire v$G32_431_out0;
wire v$G32_432_out0;
wire v$G32_433_out0;
wire v$G32_434_out0;
wire v$G32_9441_out0;
wire v$G32_9442_out0;
wire v$G33_11239_out0;
wire v$G33_11240_out0;
wire v$G33_13675_out0;
wire v$G33_13676_out0;
wire v$G33_13677_out0;
wire v$G33_13678_out0;
wire v$G33_13679_out0;
wire v$G33_13680_out0;
wire v$G33_13681_out0;
wire v$G33_13682_out0;
wire v$G33_13683_out0;
wire v$G33_13684_out0;
wire v$G33_13685_out0;
wire v$G33_13686_out0;
wire v$G33_13687_out0;
wire v$G33_13688_out0;
wire v$G33_13689_out0;
wire v$G33_13690_out0;
wire v$G33_13691_out0;
wire v$G33_13692_out0;
wire v$G33_13693_out0;
wire v$G33_13694_out0;
wire v$G33_13695_out0;
wire v$G33_13696_out0;
wire v$G33_13697_out0;
wire v$G33_13698_out0;
wire v$G33_1384_out0;
wire v$G33_1385_out0;
wire v$G33_19227_out0;
wire v$G33_19228_out0;
wire v$G33_338_out0;
wire v$G33_339_out0;
wire v$G33_5348_out0;
wire v$G33_5349_out0;
wire v$G34_1727_out0;
wire v$G34_1728_out0;
wire v$G34_17931_out0;
wire v$G34_17932_out0;
wire v$G34_17933_out0;
wire v$G34_17934_out0;
wire v$G34_17935_out0;
wire v$G34_17936_out0;
wire v$G34_17937_out0;
wire v$G34_17938_out0;
wire v$G34_17939_out0;
wire v$G34_17940_out0;
wire v$G34_17941_out0;
wire v$G34_17942_out0;
wire v$G34_17943_out0;
wire v$G34_17944_out0;
wire v$G34_17945_out0;
wire v$G34_17946_out0;
wire v$G34_17947_out0;
wire v$G34_17948_out0;
wire v$G34_17949_out0;
wire v$G34_17950_out0;
wire v$G34_17951_out0;
wire v$G34_17952_out0;
wire v$G34_17953_out0;
wire v$G34_17954_out0;
wire v$G34_5096_out0;
wire v$G34_5097_out0;
wire v$G34_5132_out0;
wire v$G34_5133_out0;
wire v$G35_10777_out0;
wire v$G35_10778_out0;
wire v$G35_1289_out0;
wire v$G35_1290_out0;
wire v$G35_13219_out0;
wire v$G35_13220_out0;
wire v$G35_15122_out0;
wire v$G35_15123_out0;
wire v$G35_15124_out0;
wire v$G35_15125_out0;
wire v$G35_15126_out0;
wire v$G35_15127_out0;
wire v$G35_15128_out0;
wire v$G35_15129_out0;
wire v$G35_15130_out0;
wire v$G35_15131_out0;
wire v$G35_15132_out0;
wire v$G35_15133_out0;
wire v$G35_15134_out0;
wire v$G35_15135_out0;
wire v$G35_15136_out0;
wire v$G35_15137_out0;
wire v$G35_15138_out0;
wire v$G35_15139_out0;
wire v$G35_15140_out0;
wire v$G35_15141_out0;
wire v$G35_15142_out0;
wire v$G35_15143_out0;
wire v$G35_15144_out0;
wire v$G35_15145_out0;
wire v$G35_19105_out0;
wire v$G35_19106_out0;
wire v$G35_4476_out0;
wire v$G35_4477_out0;
wire v$G36_11364_out0;
wire v$G36_11365_out0;
wire v$G36_14715_out0;
wire v$G36_14716_out0;
wire v$G36_17318_out0;
wire v$G36_17991_out0;
wire v$G36_17992_out0;
wire v$G36_6184_out0;
wire v$G36_6185_out0;
wire v$G36_6186_out0;
wire v$G36_6187_out0;
wire v$G36_6188_out0;
wire v$G36_6189_out0;
wire v$G36_6190_out0;
wire v$G36_6191_out0;
wire v$G36_6192_out0;
wire v$G36_6193_out0;
wire v$G36_6194_out0;
wire v$G36_6195_out0;
wire v$G36_6196_out0;
wire v$G36_6197_out0;
wire v$G36_6198_out0;
wire v$G36_6199_out0;
wire v$G36_6200_out0;
wire v$G36_6201_out0;
wire v$G36_6202_out0;
wire v$G36_6203_out0;
wire v$G36_6204_out0;
wire v$G36_6205_out0;
wire v$G36_6206_out0;
wire v$G36_6207_out0;
wire v$G36_8364_out0;
wire v$G36_8365_out0;
wire v$G37_14699_out0;
wire v$G37_14700_out0;
wire v$G37_1523_out0;
wire v$G37_1524_out0;
wire v$G37_1671_out0;
wire v$G37_1672_out0;
wire v$G37_1673_out0;
wire v$G37_1674_out0;
wire v$G37_19073_out0;
wire v$G37_19074_out0;
wire v$G37_748_out0;
wire v$G37_749_out0;
wire v$G38_10705_out0;
wire v$G38_10706_out0;
wire v$G38_7609_out0;
wire v$G38_7610_out0;
wire v$G38_7611_out0;
wire v$G38_7612_out0;
wire v$G38_7613_out0;
wire v$G38_7614_out0;
wire v$G38_7615_out0;
wire v$G38_7616_out0;
wire v$G38_7617_out0;
wire v$G38_7618_out0;
wire v$G38_7619_out0;
wire v$G38_7620_out0;
wire v$G38_7621_out0;
wire v$G38_7622_out0;
wire v$G38_7623_out0;
wire v$G38_7624_out0;
wire v$G38_7625_out0;
wire v$G38_7626_out0;
wire v$G38_7627_out0;
wire v$G38_7628_out0;
wire v$G38_7629_out0;
wire v$G38_7630_out0;
wire v$G38_7631_out0;
wire v$G38_7632_out0;
wire v$G39_17501_out0;
wire v$G39_17502_out0;
wire v$G39_18001_out0;
wire v$G39_18002_out0;
wire v$G39_18003_out0;
wire v$G39_18004_out0;
wire v$G39_6326_out0;
wire v$G39_6327_out0;
wire v$G3_0_out0;
wire v$G3_10364_out0;
wire v$G3_10365_out0;
wire v$G3_10685_out0;
wire v$G3_10686_out0;
wire v$G3_11496_out0;
wire v$G3_11497_out0;
wire v$G3_11602_out0;
wire v$G3_11603_out0;
wire v$G3_11604_out0;
wire v$G3_11605_out0;
wire v$G3_11606_out0;
wire v$G3_11607_out0;
wire v$G3_13244_out0;
wire v$G3_13245_out0;
wire v$G3_13246_out0;
wire v$G3_13247_out0;
wire v$G3_13248_out0;
wire v$G3_13249_out0;
wire v$G3_13250_out0;
wire v$G3_13251_out0;
wire v$G3_13252_out0;
wire v$G3_13253_out0;
wire v$G3_13254_out0;
wire v$G3_13255_out0;
wire v$G3_13256_out0;
wire v$G3_13257_out0;
wire v$G3_13258_out0;
wire v$G3_13259_out0;
wire v$G3_13260_out0;
wire v$G3_13261_out0;
wire v$G3_13262_out0;
wire v$G3_13263_out0;
wire v$G3_13264_out0;
wire v$G3_13265_out0;
wire v$G3_13266_out0;
wire v$G3_13267_out0;
wire v$G3_13268_out0;
wire v$G3_13269_out0;
wire v$G3_13270_out0;
wire v$G3_13271_out0;
wire v$G3_13272_out0;
wire v$G3_13273_out0;
wire v$G3_13274_out0;
wire v$G3_13275_out0;
wire v$G3_13276_out0;
wire v$G3_13277_out0;
wire v$G3_13278_out0;
wire v$G3_13279_out0;
wire v$G3_13520_out0;
wire v$G3_13521_out0;
wire v$G3_13637_out0;
wire v$G3_13638_out0;
wire v$G3_13639_out0;
wire v$G3_13640_out0;
wire v$G3_14794_out0;
wire v$G3_14795_out0;
wire v$G3_16441_out0;
wire v$G3_16442_out0;
wire v$G3_16620_out0;
wire v$G3_16621_out0;
wire v$G3_16702_out0;
wire v$G3_18094_out0;
wire v$G3_18095_out0;
wire v$G3_18293_out0;
wire v$G3_18294_out0;
wire v$G3_18295_out0;
wire v$G3_18296_out0;
wire v$G3_18297_out0;
wire v$G3_18298_out0;
wire v$G3_18299_out0;
wire v$G3_19021_out0;
wire v$G3_19022_out0;
wire v$G3_1_out0;
wire v$G3_20_out0;
wire v$G3_21_out0;
wire v$G3_2634_out0;
wire v$G3_2635_out0;
wire v$G3_2800_out0;
wire v$G3_2801_out0;
wire v$G3_2802_out0;
wire v$G3_2803_out0;
wire v$G3_2804_out0;
wire v$G3_2805_out0;
wire v$G3_2806_out0;
wire v$G3_2807_out0;
wire v$G3_2868_out0;
wire v$G3_2869_out0;
wire v$G3_3187_out0;
wire v$G3_4110_out0;
wire v$G3_4111_out0;
wire v$G3_4120_out0;
wire v$G3_4121_out0;
wire v$G3_4262_out0;
wire v$G3_4263_out0;
wire v$G3_4935_out0;
wire v$G3_4936_out0;
wire v$G3_5216_out0;
wire v$G3_7804_out0;
wire v$G3_7805_out0;
wire v$G3_7806_out0;
wire v$G3_7807_out0;
wire v$G3_7838_out0;
wire v$G3_7839_out0;
wire v$G3_7926_out0;
wire v$G3_7927_out0;
wire v$G3_8354_out0;
wire v$G3_8355_out0;
wire v$G3_9159_out0;
wire v$G3_9160_out0;
wire v$G3_9161_out0;
wire v$G3_9162_out0;
wire v$G3_9163_out0;
wire v$G3_9164_out0;
wire v$G3_9165_out0;
wire v$G3_9166_out0;
wire v$G3_9167_out0;
wire v$G3_9168_out0;
wire v$G3_9809_out0;
wire v$G3_9810_out0;
wire v$G40_13945_out0;
wire v$G40_13946_out0;
wire v$G40_13947_out0;
wire v$G40_13948_out0;
wire v$G40_13949_out0;
wire v$G40_13950_out0;
wire v$G40_13951_out0;
wire v$G40_13952_out0;
wire v$G40_13953_out0;
wire v$G40_13954_out0;
wire v$G40_13955_out0;
wire v$G40_13956_out0;
wire v$G40_13957_out0;
wire v$G40_13958_out0;
wire v$G40_13959_out0;
wire v$G40_13960_out0;
wire v$G40_13961_out0;
wire v$G40_13962_out0;
wire v$G40_13963_out0;
wire v$G40_13964_out0;
wire v$G40_13965_out0;
wire v$G40_13966_out0;
wire v$G40_13967_out0;
wire v$G40_13968_out0;
wire v$G40_14259_out0;
wire v$G40_14260_out0;
wire v$G40_15739_out0;
wire v$G40_15740_out0;
wire v$G41_11374_out0;
wire v$G41_11375_out0;
wire v$G41_11376_out0;
wire v$G41_11377_out0;
wire v$G41_11378_out0;
wire v$G41_11379_out0;
wire v$G41_11380_out0;
wire v$G41_11381_out0;
wire v$G41_11382_out0;
wire v$G41_11383_out0;
wire v$G41_11384_out0;
wire v$G41_11385_out0;
wire v$G41_11386_out0;
wire v$G41_11387_out0;
wire v$G41_11388_out0;
wire v$G41_11389_out0;
wire v$G41_11390_out0;
wire v$G41_11391_out0;
wire v$G41_11392_out0;
wire v$G41_11393_out0;
wire v$G41_11394_out0;
wire v$G41_11395_out0;
wire v$G41_11396_out0;
wire v$G41_11397_out0;
wire v$G41_19089_out0;
wire v$G41_19090_out0;
wire v$G42_19085_out0;
wire v$G42_19086_out0;
wire v$G42_9958_out0;
wire v$G42_9959_out0;
wire v$G43_409_out0;
wire v$G43_410_out0;
wire v$G43_7337_out0;
wire v$G43_7338_out0;
wire v$G44_8561_out0;
wire v$G45_15949_out0;
wire v$G45_17511_out0;
wire v$G45_17512_out0;
wire v$G46_11405_out0;
wire v$G46_11406_out0;
wire v$G46_16729_out0;
wire v$G46_16730_out0;
wire v$G47_1685_out0;
wire v$G47_1686_out0;
wire v$G47_5660_out0;
wire v$G47_5661_out0;
wire v$G48_19127_out0;
wire v$G48_19128_out0;
wire v$G48_2487_out0;
wire v$G48_2488_out0;
wire v$G48_5092_out0;
wire v$G48_5093_out0;
wire v$G49_10904_out0;
wire v$G49_10905_out0;
wire v$G49_11564_out0;
wire v$G49_11565_out0;
wire v$G49_5461_out0;
wire v$G49_5462_out0;
wire v$G4_11610_out0;
wire v$G4_11611_out0;
wire v$G4_11612_out0;
wire v$G4_11613_out0;
wire v$G4_11614_out0;
wire v$G4_11615_out0;
wire v$G4_11616_out0;
wire v$G4_11617_out0;
wire v$G4_11618_out0;
wire v$G4_11619_out0;
wire v$G4_11620_out0;
wire v$G4_11621_out0;
wire v$G4_11622_out0;
wire v$G4_11623_out0;
wire v$G4_11624_out0;
wire v$G4_11625_out0;
wire v$G4_11626_out0;
wire v$G4_11627_out0;
wire v$G4_11628_out0;
wire v$G4_11629_out0;
wire v$G4_11630_out0;
wire v$G4_11631_out0;
wire v$G4_11632_out0;
wire v$G4_11633_out0;
wire v$G4_11634_out0;
wire v$G4_11635_out0;
wire v$G4_11636_out0;
wire v$G4_11637_out0;
wire v$G4_11638_out0;
wire v$G4_11639_out0;
wire v$G4_11640_out0;
wire v$G4_11641_out0;
wire v$G4_11642_out0;
wire v$G4_11643_out0;
wire v$G4_11644_out0;
wire v$G4_11645_out0;
wire v$G4_11646_out0;
wire v$G4_11647_out0;
wire v$G4_11648_out0;
wire v$G4_11649_out0;
wire v$G4_11650_out0;
wire v$G4_11651_out0;
wire v$G4_11652_out0;
wire v$G4_11653_out0;
wire v$G4_11654_out0;
wire v$G4_11655_out0;
wire v$G4_11656_out0;
wire v$G4_11657_out0;
wire v$G4_11658_out0;
wire v$G4_11659_out0;
wire v$G4_11660_out0;
wire v$G4_11661_out0;
wire v$G4_11662_out0;
wire v$G4_11663_out0;
wire v$G4_11664_out0;
wire v$G4_11665_out0;
wire v$G4_11666_out0;
wire v$G4_11667_out0;
wire v$G4_11668_out0;
wire v$G4_11669_out0;
wire v$G4_11670_out0;
wire v$G4_11671_out0;
wire v$G4_11672_out0;
wire v$G4_11673_out0;
wire v$G4_11674_out0;
wire v$G4_11675_out0;
wire v$G4_11676_out0;
wire v$G4_11677_out0;
wire v$G4_11678_out0;
wire v$G4_11679_out0;
wire v$G4_11680_out0;
wire v$G4_11681_out0;
wire v$G4_11682_out0;
wire v$G4_11683_out0;
wire v$G4_11684_out0;
wire v$G4_11685_out0;
wire v$G4_11686_out0;
wire v$G4_11687_out0;
wire v$G4_11688_out0;
wire v$G4_11689_out0;
wire v$G4_11690_out0;
wire v$G4_11691_out0;
wire v$G4_11692_out0;
wire v$G4_11693_out0;
wire v$G4_11694_out0;
wire v$G4_11695_out0;
wire v$G4_11696_out0;
wire v$G4_11697_out0;
wire v$G4_11698_out0;
wire v$G4_11699_out0;
wire v$G4_11700_out0;
wire v$G4_11701_out0;
wire v$G4_11702_out0;
wire v$G4_11703_out0;
wire v$G4_11704_out0;
wire v$G4_11705_out0;
wire v$G4_11706_out0;
wire v$G4_11707_out0;
wire v$G4_11708_out0;
wire v$G4_11709_out0;
wire v$G4_11710_out0;
wire v$G4_11711_out0;
wire v$G4_11712_out0;
wire v$G4_11713_out0;
wire v$G4_11714_out0;
wire v$G4_11715_out0;
wire v$G4_11716_out0;
wire v$G4_11717_out0;
wire v$G4_11718_out0;
wire v$G4_11719_out0;
wire v$G4_11720_out0;
wire v$G4_11721_out0;
wire v$G4_11722_out0;
wire v$G4_11723_out0;
wire v$G4_11724_out0;
wire v$G4_11725_out0;
wire v$G4_11726_out0;
wire v$G4_11727_out0;
wire v$G4_11728_out0;
wire v$G4_11729_out0;
wire v$G4_11730_out0;
wire v$G4_11731_out0;
wire v$G4_11732_out0;
wire v$G4_11733_out0;
wire v$G4_11734_out0;
wire v$G4_11735_out0;
wire v$G4_11736_out0;
wire v$G4_11737_out0;
wire v$G4_11738_out0;
wire v$G4_11739_out0;
wire v$G4_11740_out0;
wire v$G4_11741_out0;
wire v$G4_11742_out0;
wire v$G4_11743_out0;
wire v$G4_11744_out0;
wire v$G4_11745_out0;
wire v$G4_11746_out0;
wire v$G4_11747_out0;
wire v$G4_11748_out0;
wire v$G4_11749_out0;
wire v$G4_11750_out0;
wire v$G4_11751_out0;
wire v$G4_11752_out0;
wire v$G4_11753_out0;
wire v$G4_11754_out0;
wire v$G4_11755_out0;
wire v$G4_11756_out0;
wire v$G4_11757_out0;
wire v$G4_11758_out0;
wire v$G4_11759_out0;
wire v$G4_11760_out0;
wire v$G4_11761_out0;
wire v$G4_11762_out0;
wire v$G4_11763_out0;
wire v$G4_11764_out0;
wire v$G4_11765_out0;
wire v$G4_11766_out0;
wire v$G4_11767_out0;
wire v$G4_11768_out0;
wire v$G4_11769_out0;
wire v$G4_11770_out0;
wire v$G4_11771_out0;
wire v$G4_11772_out0;
wire v$G4_11773_out0;
wire v$G4_11774_out0;
wire v$G4_11775_out0;
wire v$G4_11776_out0;
wire v$G4_11777_out0;
wire v$G4_11778_out0;
wire v$G4_11779_out0;
wire v$G4_11780_out0;
wire v$G4_11781_out0;
wire v$G4_11782_out0;
wire v$G4_11783_out0;
wire v$G4_11784_out0;
wire v$G4_11785_out0;
wire v$G4_11786_out0;
wire v$G4_11787_out0;
wire v$G4_11788_out0;
wire v$G4_11789_out0;
wire v$G4_11790_out0;
wire v$G4_11791_out0;
wire v$G4_11792_out0;
wire v$G4_11793_out0;
wire v$G4_11794_out0;
wire v$G4_11795_out0;
wire v$G4_11796_out0;
wire v$G4_11797_out0;
wire v$G4_11798_out0;
wire v$G4_11799_out0;
wire v$G4_11800_out0;
wire v$G4_11801_out0;
wire v$G4_11802_out0;
wire v$G4_11803_out0;
wire v$G4_11804_out0;
wire v$G4_11805_out0;
wire v$G4_11806_out0;
wire v$G4_11807_out0;
wire v$G4_11808_out0;
wire v$G4_11809_out0;
wire v$G4_11810_out0;
wire v$G4_11811_out0;
wire v$G4_11812_out0;
wire v$G4_11813_out0;
wire v$G4_11814_out0;
wire v$G4_11815_out0;
wire v$G4_11816_out0;
wire v$G4_11817_out0;
wire v$G4_11818_out0;
wire v$G4_11819_out0;
wire v$G4_11820_out0;
wire v$G4_11821_out0;
wire v$G4_11822_out0;
wire v$G4_11823_out0;
wire v$G4_11824_out0;
wire v$G4_11825_out0;
wire v$G4_11826_out0;
wire v$G4_11827_out0;
wire v$G4_11828_out0;
wire v$G4_11829_out0;
wire v$G4_11830_out0;
wire v$G4_11831_out0;
wire v$G4_11832_out0;
wire v$G4_11833_out0;
wire v$G4_11834_out0;
wire v$G4_11835_out0;
wire v$G4_11836_out0;
wire v$G4_11837_out0;
wire v$G4_11838_out0;
wire v$G4_11839_out0;
wire v$G4_11840_out0;
wire v$G4_11841_out0;
wire v$G4_11842_out0;
wire v$G4_11843_out0;
wire v$G4_11844_out0;
wire v$G4_11845_out0;
wire v$G4_11846_out0;
wire v$G4_11847_out0;
wire v$G4_11848_out0;
wire v$G4_11849_out0;
wire v$G4_11850_out0;
wire v$G4_11851_out0;
wire v$G4_11852_out0;
wire v$G4_11853_out0;
wire v$G4_11854_out0;
wire v$G4_11855_out0;
wire v$G4_12405_out0;
wire v$G4_12406_out0;
wire v$G4_12407_out0;
wire v$G4_12408_out0;
wire v$G4_12409_out0;
wire v$G4_12410_out0;
wire v$G4_12411_out0;
wire v$G4_12412_out0;
wire v$G4_12413_out0;
wire v$G4_12414_out0;
wire v$G4_12443_out0;
wire v$G4_12444_out0;
wire v$G4_12565_out0;
wire v$G4_12566_out0;
wire v$G4_13766_out0;
wire v$G4_14607_out0;
wire v$G4_14608_out0;
wire v$G4_14816_out0;
wire v$G4_14817_out0;
wire v$G4_1491_out0;
wire v$G4_1492_out0;
wire v$G4_15100_out0;
wire v$G4_15101_out0;
wire v$G4_15287_out0;
wire v$G4_15288_out0;
wire v$G4_15735_out0;
wire v$G4_15736_out0;
wire v$G4_15927_out0;
wire v$G4_15928_out0;
wire v$G4_16044_out0;
wire v$G4_16045_out0;
wire v$G4_16135_out0;
wire v$G4_16136_out0;
wire v$G4_16428_out0;
wire v$G4_16429_out0;
wire v$G4_18158_out0;
wire v$G4_18159_out0;
wire v$G4_18160_out0;
wire v$G4_18161_out0;
wire v$G4_18162_out0;
wire v$G4_18163_out0;
wire v$G4_18164_out0;
wire v$G4_18165_out0;
wire v$G4_18166_out0;
wire v$G4_18167_out0;
wire v$G4_18168_out0;
wire v$G4_18169_out0;
wire v$G4_18170_out0;
wire v$G4_18171_out0;
wire v$G4_18172_out0;
wire v$G4_18173_out0;
wire v$G4_18174_out0;
wire v$G4_18175_out0;
wire v$G4_18176_out0;
wire v$G4_18177_out0;
wire v$G4_18178_out0;
wire v$G4_18179_out0;
wire v$G4_18180_out0;
wire v$G4_18181_out0;
wire v$G4_18182_out0;
wire v$G4_18183_out0;
wire v$G4_18184_out0;
wire v$G4_18185_out0;
wire v$G4_18186_out0;
wire v$G4_18187_out0;
wire v$G4_18188_out0;
wire v$G4_18189_out0;
wire v$G4_18190_out0;
wire v$G4_18191_out0;
wire v$G4_18192_out0;
wire v$G4_18193_out0;
wire v$G4_18209_out0;
wire v$G4_18210_out0;
wire v$G4_18881_out0;
wire v$G4_18882_out0;
wire v$G4_3096_out0;
wire v$G4_3097_out0;
wire v$G4_4186_out0;
wire v$G4_4187_out0;
wire v$G4_4188_out0;
wire v$G4_4189_out0;
wire v$G4_4190_out0;
wire v$G4_4191_out0;
wire v$G4_4192_out0;
wire v$G4_4193_out0;
wire v$G4_5116_out0;
wire v$G4_5117_out0;
wire v$G4_6019_out0;
wire v$G4_6020_out0;
wire v$G4_6021_out0;
wire v$G4_6022_out0;
wire v$G4_6023_out0;
wire v$G4_6024_out0;
wire v$G4_6334_out0;
wire v$G4_6335_out0;
wire v$G4_6336_out0;
wire v$G4_6337_out0;
wire v$G4_6660_out0;
wire v$G4_7870_out0;
wire v$G4_7871_out0;
wire v$G4_8057_out0;
wire v$G4_8058_out0;
wire v$G50_13791_out0;
wire v$G50_13792_out0;
wire v$G50_13889_out0;
wire v$G50_16979_out0;
wire v$G50_16980_out0;
wire v$G50_17963_out0;
wire v$G50_17964_out0;
wire v$G51_14624_out0;
wire v$G51_14625_out0;
wire v$G51_19373_out0;
wire v$G51_3076_out0;
wire v$G51_3077_out0;
wire v$G51_3675_out0;
wire v$G51_3676_out0;
wire v$G52_16544_out0;
wire v$G52_16545_out0;
wire v$G52_3181_out0;
wire v$G52_3182_out0;
wire v$G52_8213_out0;
wire v$G53_13284_out0;
wire v$G53_13285_out0;
wire v$G53_16434_out0;
wire v$G53_16435_out0;
wire v$G53_18133_out0;
wire v$G54_13869_out0;
wire v$G54_14798_out0;
wire v$G54_14799_out0;
wire v$G54_2064_out0;
wire v$G54_2065_out0;
wire v$G54_8437_out0;
wire v$G54_8438_out0;
wire v$G55_14278_out0;
wire v$G55_17278_out0;
wire v$G55_17279_out0;
wire v$G55_18799_out0;
wire v$G55_18800_out0;
wire v$G55_5265_out0;
wire v$G55_5266_out0;
wire v$G56_18278_out0;
wire v$G56_3361_out0;
wire v$G56_3362_out0;
wire v$G56_708_out0;
wire v$G56_709_out0;
wire v$G57_12214_out0;
wire v$G57_12215_out0;
wire v$G57_14037_out0;
wire v$G57_14038_out0;
wire v$G57_18569_out0;
wire v$G57_9305_out0;
wire v$G57_9306_out0;
wire v$G58_168_out0;
wire v$G58_169_out0;
wire v$G58_2714_out0;
wire v$G58_2715_out0;
wire v$G58_7333_out0;
wire v$G58_7334_out0;
wire v$G59_15731_out0;
wire v$G59_15732_out0;
wire v$G59_2763_out0;
wire v$G59_4024_out0;
wire v$G59_4025_out0;
wire v$G5_11170_out0;
wire v$G5_11171_out0;
wire v$G5_11172_out0;
wire v$G5_11173_out0;
wire v$G5_11174_out0;
wire v$G5_11175_out0;
wire v$G5_11186_out0;
wire v$G5_11187_out0;
wire v$G5_1267_out0;
wire v$G5_1268_out0;
wire v$G5_1269_out0;
wire v$G5_1270_out0;
wire v$G5_1271_out0;
wire v$G5_1272_out0;
wire v$G5_1273_out0;
wire v$G5_1274_out0;
wire v$G5_1275_out0;
wire v$G5_1276_out0;
wire v$G5_13317_out0;
wire v$G5_13318_out0;
wire v$G5_14126_out0;
wire v$G5_14127_out0;
wire v$G5_15253_out0;
wire v$G5_15254_out0;
wire v$G5_15257_out0;
wire v$G5_15258_out0;
wire v$G5_15815_out0;
wire v$G5_15816_out0;
wire v$G5_16393_out0;
wire v$G5_16394_out0;
wire v$G5_16731_out0;
wire v$G5_16732_out0;
wire v$G5_16764_out0;
wire v$G5_16765_out0;
wire v$G5_17176_out0;
wire v$G5_17177_out0;
wire v$G5_18148_out0;
wire v$G5_18149_out0;
wire v$G5_18150_out0;
wire v$G5_18151_out0;
wire v$G5_18490_out0;
wire v$G5_18491_out0;
wire v$G5_2440_out0;
wire v$G5_2441_out0;
wire v$G5_2865_out0;
wire v$G5_4689_out0;
wire v$G5_4690_out0;
wire v$G5_4691_out0;
wire v$G5_4692_out0;
wire v$G5_4693_out0;
wire v$G5_4694_out0;
wire v$G5_4695_out0;
wire v$G5_4696_out0;
wire v$G5_4697_out0;
wire v$G5_4698_out0;
wire v$G5_4699_out0;
wire v$G5_4700_out0;
wire v$G5_4701_out0;
wire v$G5_4702_out0;
wire v$G5_4703_out0;
wire v$G5_4704_out0;
wire v$G5_4705_out0;
wire v$G5_4706_out0;
wire v$G5_4707_out0;
wire v$G5_4708_out0;
wire v$G5_4709_out0;
wire v$G5_4710_out0;
wire v$G5_4711_out0;
wire v$G5_4712_out0;
wire v$G5_4713_out0;
wire v$G5_4714_out0;
wire v$G5_4715_out0;
wire v$G5_4716_out0;
wire v$G5_4717_out0;
wire v$G5_4718_out0;
wire v$G5_4719_out0;
wire v$G5_4720_out0;
wire v$G5_4721_out0;
wire v$G5_4722_out0;
wire v$G5_4723_out0;
wire v$G5_4724_out0;
wire v$G5_4725_out0;
wire v$G5_4726_out0;
wire v$G5_4727_out0;
wire v$G5_4728_out0;
wire v$G5_4729_out0;
wire v$G5_4730_out0;
wire v$G5_4731_out0;
wire v$G5_4732_out0;
wire v$G5_4733_out0;
wire v$G5_4734_out0;
wire v$G5_4735_out0;
wire v$G5_4736_out0;
wire v$G5_4737_out0;
wire v$G5_4738_out0;
wire v$G5_4739_out0;
wire v$G5_4740_out0;
wire v$G5_4741_out0;
wire v$G5_4742_out0;
wire v$G5_4743_out0;
wire v$G5_4744_out0;
wire v$G5_4745_out0;
wire v$G5_4746_out0;
wire v$G5_4747_out0;
wire v$G5_4748_out0;
wire v$G5_4749_out0;
wire v$G5_4750_out0;
wire v$G5_4751_out0;
wire v$G5_4752_out0;
wire v$G5_4753_out0;
wire v$G5_4754_out0;
wire v$G5_4755_out0;
wire v$G5_4756_out0;
wire v$G5_4757_out0;
wire v$G5_4758_out0;
wire v$G5_4759_out0;
wire v$G5_4760_out0;
wire v$G5_4761_out0;
wire v$G5_4762_out0;
wire v$G5_4763_out0;
wire v$G5_4764_out0;
wire v$G5_4765_out0;
wire v$G5_4766_out0;
wire v$G5_4767_out0;
wire v$G5_4768_out0;
wire v$G5_4769_out0;
wire v$G5_4770_out0;
wire v$G5_4771_out0;
wire v$G5_4772_out0;
wire v$G5_4773_out0;
wire v$G5_4774_out0;
wire v$G5_4775_out0;
wire v$G5_4776_out0;
wire v$G5_4777_out0;
wire v$G5_4778_out0;
wire v$G5_4779_out0;
wire v$G5_4780_out0;
wire v$G5_4781_out0;
wire v$G5_4782_out0;
wire v$G5_4783_out0;
wire v$G5_4784_out0;
wire v$G5_4785_out0;
wire v$G5_4786_out0;
wire v$G5_4787_out0;
wire v$G5_4788_out0;
wire v$G5_4789_out0;
wire v$G5_4790_out0;
wire v$G5_4791_out0;
wire v$G5_4792_out0;
wire v$G5_4793_out0;
wire v$G5_4794_out0;
wire v$G5_4795_out0;
wire v$G5_4796_out0;
wire v$G5_4797_out0;
wire v$G5_4798_out0;
wire v$G5_4799_out0;
wire v$G5_4800_out0;
wire v$G5_4801_out0;
wire v$G5_4802_out0;
wire v$G5_4803_out0;
wire v$G5_4804_out0;
wire v$G5_4805_out0;
wire v$G5_4806_out0;
wire v$G5_4807_out0;
wire v$G5_4808_out0;
wire v$G5_4809_out0;
wire v$G5_4810_out0;
wire v$G5_4811_out0;
wire v$G5_4812_out0;
wire v$G5_4813_out0;
wire v$G5_4814_out0;
wire v$G5_4815_out0;
wire v$G5_4816_out0;
wire v$G5_4817_out0;
wire v$G5_4818_out0;
wire v$G5_4819_out0;
wire v$G5_4820_out0;
wire v$G5_4821_out0;
wire v$G5_4822_out0;
wire v$G5_4823_out0;
wire v$G5_4824_out0;
wire v$G5_4825_out0;
wire v$G5_4826_out0;
wire v$G5_4827_out0;
wire v$G5_4828_out0;
wire v$G5_4829_out0;
wire v$G5_4830_out0;
wire v$G5_4831_out0;
wire v$G5_4832_out0;
wire v$G5_4833_out0;
wire v$G5_4834_out0;
wire v$G5_4835_out0;
wire v$G5_4836_out0;
wire v$G5_4837_out0;
wire v$G5_4838_out0;
wire v$G5_4839_out0;
wire v$G5_4840_out0;
wire v$G5_4841_out0;
wire v$G5_4842_out0;
wire v$G5_4843_out0;
wire v$G5_4844_out0;
wire v$G5_4845_out0;
wire v$G5_4846_out0;
wire v$G5_4847_out0;
wire v$G5_4848_out0;
wire v$G5_4849_out0;
wire v$G5_4850_out0;
wire v$G5_4851_out0;
wire v$G5_4852_out0;
wire v$G5_4853_out0;
wire v$G5_4854_out0;
wire v$G5_4855_out0;
wire v$G5_4856_out0;
wire v$G5_4857_out0;
wire v$G5_4858_out0;
wire v$G5_4859_out0;
wire v$G5_4860_out0;
wire v$G5_4861_out0;
wire v$G5_4862_out0;
wire v$G5_4863_out0;
wire v$G5_4864_out0;
wire v$G5_4865_out0;
wire v$G5_4866_out0;
wire v$G5_4867_out0;
wire v$G5_4868_out0;
wire v$G5_4869_out0;
wire v$G5_4870_out0;
wire v$G5_4871_out0;
wire v$G5_4872_out0;
wire v$G5_4873_out0;
wire v$G5_4874_out0;
wire v$G5_4875_out0;
wire v$G5_4876_out0;
wire v$G5_4877_out0;
wire v$G5_4878_out0;
wire v$G5_4879_out0;
wire v$G5_4880_out0;
wire v$G5_4881_out0;
wire v$G5_4882_out0;
wire v$G5_4883_out0;
wire v$G5_4884_out0;
wire v$G5_4885_out0;
wire v$G5_4886_out0;
wire v$G5_4887_out0;
wire v$G5_4888_out0;
wire v$G5_4889_out0;
wire v$G5_4890_out0;
wire v$G5_4891_out0;
wire v$G5_4892_out0;
wire v$G5_4893_out0;
wire v$G5_4894_out0;
wire v$G5_4895_out0;
wire v$G5_4896_out0;
wire v$G5_4897_out0;
wire v$G5_4898_out0;
wire v$G5_4899_out0;
wire v$G5_4900_out0;
wire v$G5_4901_out0;
wire v$G5_4902_out0;
wire v$G5_4903_out0;
wire v$G5_4904_out0;
wire v$G5_4905_out0;
wire v$G5_4906_out0;
wire v$G5_4907_out0;
wire v$G5_4908_out0;
wire v$G5_4909_out0;
wire v$G5_4910_out0;
wire v$G5_4911_out0;
wire v$G5_4912_out0;
wire v$G5_4913_out0;
wire v$G5_4914_out0;
wire v$G5_4915_out0;
wire v$G5_4916_out0;
wire v$G5_4917_out0;
wire v$G5_4918_out0;
wire v$G5_4919_out0;
wire v$G5_4920_out0;
wire v$G5_4921_out0;
wire v$G5_4922_out0;
wire v$G5_4923_out0;
wire v$G5_4924_out0;
wire v$G5_4925_out0;
wire v$G5_4926_out0;
wire v$G5_4927_out0;
wire v$G5_4928_out0;
wire v$G5_4929_out0;
wire v$G5_4930_out0;
wire v$G5_4931_out0;
wire v$G5_4932_out0;
wire v$G5_4933_out0;
wire v$G5_4934_out0;
wire v$G5_6084_out0;
wire v$G5_6119_out0;
wire v$G5_6120_out0;
wire v$G5_6121_out0;
wire v$G5_6122_out0;
wire v$G5_6123_out0;
wire v$G5_6124_out0;
wire v$G5_6125_out0;
wire v$G5_6126_out0;
wire v$G5_6127_out0;
wire v$G5_6128_out0;
wire v$G5_6129_out0;
wire v$G5_6130_out0;
wire v$G5_6131_out0;
wire v$G5_6132_out0;
wire v$G5_6133_out0;
wire v$G5_6134_out0;
wire v$G5_6135_out0;
wire v$G5_6136_out0;
wire v$G5_6137_out0;
wire v$G5_6138_out0;
wire v$G5_6139_out0;
wire v$G5_6140_out0;
wire v$G5_6141_out0;
wire v$G5_6142_out0;
wire v$G5_6143_out0;
wire v$G5_6144_out0;
wire v$G5_6145_out0;
wire v$G5_6146_out0;
wire v$G5_6147_out0;
wire v$G5_6148_out0;
wire v$G5_6149_out0;
wire v$G5_6150_out0;
wire v$G5_6151_out0;
wire v$G5_6152_out0;
wire v$G5_6153_out0;
wire v$G5_6154_out0;
wire v$G5_6460_out0;
wire v$G5_6461_out0;
wire v$G5_7215_out0;
wire v$G5_7216_out0;
wire v$G5_7217_out0;
wire v$G5_7218_out0;
wire v$G5_7219_out0;
wire v$G5_7220_out0;
wire v$G5_7221_out0;
wire v$G5_7222_out0;
wire v$G5_7223_out0;
wire v$G5_7224_out0;
wire v$G5_7225_out0;
wire v$G5_7226_out0;
wire v$G5_7227_out0;
wire v$G5_7228_out0;
wire v$G5_7229_out0;
wire v$G5_7230_out0;
wire v$G5_7231_out0;
wire v$G5_7232_out0;
wire v$G5_7233_out0;
wire v$G5_7234_out0;
wire v$G5_7235_out0;
wire v$G5_7236_out0;
wire v$G5_7237_out0;
wire v$G5_7238_out0;
wire v$G5_7910_out0;
wire v$G5_7911_out0;
wire v$G5_8754_out0;
wire v$G5_8755_out0;
wire v$G60_19369_out0;
wire v$G60_19370_out0;
wire v$G60_9841_out0;
wire v$G60_9842_out0;
wire v$G61_12174_out0;
wire v$G61_12175_out0;
wire v$G61_17069_out0;
wire v$G61_17070_out0;
wire v$G61_8592_out0;
wire v$G61_8593_out0;
wire v$G62_12324_out0;
wire v$G62_12325_out0;
wire v$G62_12543_out0;
wire v$G62_15602_out0;
wire v$G62_15603_out0;
wire v$G63_10444_out0;
wire v$G63_10445_out0;
wire v$G63_14258_out0;
wire v$G63_17433_out0;
wire v$G63_17434_out0;
wire v$G64_15843_out0;
wire v$G64_15844_out0;
wire v$G64_6638_out0;
wire v$G64_6639_out0;
wire v$G64_6675_out0;
wire v$G64_8104_out0;
wire v$G64_8105_out0;
wire v$G65_14732_out0;
wire v$G65_14733_out0;
wire v$G65_18812_out0;
wire v$G65_18813_out0;
wire v$G65_2654_out0;
wire v$G65_2655_out0;
wire v$G65_9154_out0;
wire v$G66_15853_out0;
wire v$G66_15854_out0;
wire v$G66_17456_out0;
wire v$G66_17457_out0;
wire v$G66_9020_out0;
wire v$G66_9021_out0;
wire v$G66_9263_out0;
wire v$G67_11571_out0;
wire v$G67_11572_out0;
wire v$G67_14340_out0;
wire v$G67_14719_out0;
wire v$G67_14720_out0;
wire v$G68_15429_out0;
wire v$G68_15784_out0;
wire v$G68_15785_out0;
wire v$G68_18717_out0;
wire v$G68_18718_out0;
wire v$G69_1355_out0;
wire v$G69_1356_out0;
wire v$G69_16415_out0;
wire v$G69_8519_out0;
wire v$G69_8520_out0;
wire v$G6_12509_out0;
wire v$G6_12510_out0;
wire v$G6_12692_out0;
wire v$G6_12693_out0;
wire v$G6_13585_out0;
wire v$G6_13586_out0;
wire v$G6_14205_out0;
wire v$G6_14206_out0;
wire v$G6_16151_out0;
wire v$G6_16152_out0;
wire v$G6_16153_out0;
wire v$G6_16154_out0;
wire v$G6_16155_out0;
wire v$G6_16156_out0;
wire v$G6_16157_out0;
wire v$G6_16158_out0;
wire v$G6_16159_out0;
wire v$G6_16160_out0;
wire v$G6_16161_out0;
wire v$G6_16162_out0;
wire v$G6_16163_out0;
wire v$G6_16164_out0;
wire v$G6_16165_out0;
wire v$G6_16166_out0;
wire v$G6_16167_out0;
wire v$G6_16168_out0;
wire v$G6_16169_out0;
wire v$G6_16170_out0;
wire v$G6_16171_out0;
wire v$G6_16172_out0;
wire v$G6_16970_out0;
wire v$G6_16971_out0;
wire v$G6_16972_out0;
wire v$G6_16973_out0;
wire v$G6_16974_out0;
wire v$G6_16975_out0;
wire v$G6_17432_out0;
wire v$G6_18041_out0;
wire v$G6_2452_out0;
wire v$G6_2453_out0;
wire v$G6_279_out0;
wire v$G6_280_out0;
wire v$G6_3383_out0;
wire v$G6_3384_out0;
wire v$G6_3580_out0;
wire v$G6_3581_out0;
wire v$G6_3703_out0;
wire v$G6_3756_out0;
wire v$G6_3757_out0;
wire v$G6_3758_out0;
wire v$G6_3759_out0;
wire v$G6_3760_out0;
wire v$G6_3761_out0;
wire v$G6_3762_out0;
wire v$G6_3763_out0;
wire v$G6_3764_out0;
wire v$G6_3765_out0;
wire v$G6_3766_out0;
wire v$G6_3767_out0;
wire v$G6_3768_out0;
wire v$G6_3769_out0;
wire v$G6_3770_out0;
wire v$G6_3771_out0;
wire v$G6_3772_out0;
wire v$G6_3773_out0;
wire v$G6_3774_out0;
wire v$G6_3775_out0;
wire v$G6_3776_out0;
wire v$G6_3777_out0;
wire v$G6_3778_out0;
wire v$G6_3779_out0;
wire v$G6_3780_out0;
wire v$G6_3781_out0;
wire v$G6_3782_out0;
wire v$G6_3783_out0;
wire v$G6_3784_out0;
wire v$G6_3785_out0;
wire v$G6_3786_out0;
wire v$G6_3787_out0;
wire v$G6_3788_out0;
wire v$G6_3789_out0;
wire v$G6_3790_out0;
wire v$G6_3791_out0;
wire v$G6_452_out0;
wire v$G6_453_out0;
wire v$G6_454_out0;
wire v$G6_455_out0;
wire v$G6_456_out0;
wire v$G6_457_out0;
wire v$G6_458_out0;
wire v$G6_459_out0;
wire v$G6_460_out0;
wire v$G6_461_out0;
wire v$G6_462_out0;
wire v$G6_463_out0;
wire v$G6_464_out0;
wire v$G6_465_out0;
wire v$G6_466_out0;
wire v$G6_467_out0;
wire v$G6_468_out0;
wire v$G6_469_out0;
wire v$G6_470_out0;
wire v$G6_471_out0;
wire v$G6_472_out0;
wire v$G6_473_out0;
wire v$G6_474_out0;
wire v$G6_475_out0;
wire v$G6_476_out0;
wire v$G6_477_out0;
wire v$G6_478_out0;
wire v$G6_479_out0;
wire v$G6_480_out0;
wire v$G6_481_out0;
wire v$G6_482_out0;
wire v$G6_483_out0;
wire v$G6_484_out0;
wire v$G6_485_out0;
wire v$G6_486_out0;
wire v$G6_487_out0;
wire v$G6_488_out0;
wire v$G6_489_out0;
wire v$G6_490_out0;
wire v$G6_491_out0;
wire v$G6_492_out0;
wire v$G6_493_out0;
wire v$G6_494_out0;
wire v$G6_495_out0;
wire v$G6_496_out0;
wire v$G6_497_out0;
wire v$G6_498_out0;
wire v$G6_499_out0;
wire v$G6_500_out0;
wire v$G6_501_out0;
wire v$G6_502_out0;
wire v$G6_503_out0;
wire v$G6_504_out0;
wire v$G6_505_out0;
wire v$G6_506_out0;
wire v$G6_507_out0;
wire v$G6_508_out0;
wire v$G6_509_out0;
wire v$G6_510_out0;
wire v$G6_511_out0;
wire v$G6_512_out0;
wire v$G6_513_out0;
wire v$G6_514_out0;
wire v$G6_515_out0;
wire v$G6_516_out0;
wire v$G6_517_out0;
wire v$G6_518_out0;
wire v$G6_519_out0;
wire v$G6_520_out0;
wire v$G6_521_out0;
wire v$G6_522_out0;
wire v$G6_523_out0;
wire v$G6_524_out0;
wire v$G6_525_out0;
wire v$G6_526_out0;
wire v$G6_527_out0;
wire v$G6_528_out0;
wire v$G6_529_out0;
wire v$G6_530_out0;
wire v$G6_531_out0;
wire v$G6_532_out0;
wire v$G6_533_out0;
wire v$G6_534_out0;
wire v$G6_535_out0;
wire v$G6_536_out0;
wire v$G6_537_out0;
wire v$G6_538_out0;
wire v$G6_539_out0;
wire v$G6_540_out0;
wire v$G6_541_out0;
wire v$G6_542_out0;
wire v$G6_543_out0;
wire v$G6_544_out0;
wire v$G6_545_out0;
wire v$G6_546_out0;
wire v$G6_547_out0;
wire v$G6_548_out0;
wire v$G6_549_out0;
wire v$G6_550_out0;
wire v$G6_551_out0;
wire v$G6_552_out0;
wire v$G6_553_out0;
wire v$G6_554_out0;
wire v$G6_555_out0;
wire v$G6_556_out0;
wire v$G6_557_out0;
wire v$G6_558_out0;
wire v$G6_559_out0;
wire v$G6_560_out0;
wire v$G6_561_out0;
wire v$G6_562_out0;
wire v$G6_563_out0;
wire v$G6_564_out0;
wire v$G6_565_out0;
wire v$G6_566_out0;
wire v$G6_567_out0;
wire v$G6_568_out0;
wire v$G6_569_out0;
wire v$G6_5703_out0;
wire v$G6_5704_out0;
wire v$G6_570_out0;
wire v$G6_571_out0;
wire v$G6_572_out0;
wire v$G6_573_out0;
wire v$G6_574_out0;
wire v$G6_575_out0;
wire v$G6_576_out0;
wire v$G6_577_out0;
wire v$G6_578_out0;
wire v$G6_579_out0;
wire v$G6_580_out0;
wire v$G6_581_out0;
wire v$G6_582_out0;
wire v$G6_583_out0;
wire v$G6_584_out0;
wire v$G6_585_out0;
wire v$G6_586_out0;
wire v$G6_587_out0;
wire v$G6_588_out0;
wire v$G6_589_out0;
wire v$G6_590_out0;
wire v$G6_591_out0;
wire v$G6_592_out0;
wire v$G6_593_out0;
wire v$G6_594_out0;
wire v$G6_595_out0;
wire v$G6_596_out0;
wire v$G6_597_out0;
wire v$G6_598_out0;
wire v$G6_599_out0;
wire v$G6_600_out0;
wire v$G6_601_out0;
wire v$G6_602_out0;
wire v$G6_603_out0;
wire v$G6_604_out0;
wire v$G6_605_out0;
wire v$G6_606_out0;
wire v$G6_607_out0;
wire v$G6_608_out0;
wire v$G6_609_out0;
wire v$G6_610_out0;
wire v$G6_611_out0;
wire v$G6_612_out0;
wire v$G6_613_out0;
wire v$G6_614_out0;
wire v$G6_615_out0;
wire v$G6_616_out0;
wire v$G6_617_out0;
wire v$G6_618_out0;
wire v$G6_619_out0;
wire v$G6_620_out0;
wire v$G6_621_out0;
wire v$G6_6224_out0;
wire v$G6_6225_out0;
wire v$G6_622_out0;
wire v$G6_623_out0;
wire v$G6_624_out0;
wire v$G6_625_out0;
wire v$G6_626_out0;
wire v$G6_627_out0;
wire v$G6_628_out0;
wire v$G6_629_out0;
wire v$G6_630_out0;
wire v$G6_631_out0;
wire v$G6_632_out0;
wire v$G6_633_out0;
wire v$G6_634_out0;
wire v$G6_635_out0;
wire v$G6_636_out0;
wire v$G6_637_out0;
wire v$G6_638_out0;
wire v$G6_639_out0;
wire v$G6_640_out0;
wire v$G6_641_out0;
wire v$G6_6428_out0;
wire v$G6_6429_out0;
wire v$G6_642_out0;
wire v$G6_6434_out0;
wire v$G6_6435_out0;
wire v$G6_6436_out0;
wire v$G6_6437_out0;
wire v$G6_6438_out0;
wire v$G6_6439_out0;
wire v$G6_643_out0;
wire v$G6_6440_out0;
wire v$G6_6441_out0;
wire v$G6_644_out0;
wire v$G6_645_out0;
wire v$G6_646_out0;
wire v$G6_647_out0;
wire v$G6_648_out0;
wire v$G6_649_out0;
wire v$G6_650_out0;
wire v$G6_651_out0;
wire v$G6_652_out0;
wire v$G6_653_out0;
wire v$G6_654_out0;
wire v$G6_655_out0;
wire v$G6_656_out0;
wire v$G6_657_out0;
wire v$G6_658_out0;
wire v$G6_659_out0;
wire v$G6_660_out0;
wire v$G6_661_out0;
wire v$G6_662_out0;
wire v$G6_663_out0;
wire v$G6_664_out0;
wire v$G6_665_out0;
wire v$G6_666_out0;
wire v$G6_667_out0;
wire v$G6_668_out0;
wire v$G6_669_out0;
wire v$G6_670_out0;
wire v$G6_671_out0;
wire v$G6_672_out0;
wire v$G6_673_out0;
wire v$G6_674_out0;
wire v$G6_675_out0;
wire v$G6_676_out0;
wire v$G6_677_out0;
wire v$G6_6783_out0;
wire v$G6_6784_out0;
wire v$G6_6785_out0;
wire v$G6_6786_out0;
wire v$G6_6787_out0;
wire v$G6_6788_out0;
wire v$G6_6789_out0;
wire v$G6_678_out0;
wire v$G6_6790_out0;
wire v$G6_6791_out0;
wire v$G6_6792_out0;
wire v$G6_6793_out0;
wire v$G6_6794_out0;
wire v$G6_6795_out0;
wire v$G6_6796_out0;
wire v$G6_6797_out0;
wire v$G6_6798_out0;
wire v$G6_6799_out0;
wire v$G6_679_out0;
wire v$G6_6800_out0;
wire v$G6_6801_out0;
wire v$G6_6802_out0;
wire v$G6_6803_out0;
wire v$G6_6804_out0;
wire v$G6_6805_out0;
wire v$G6_6806_out0;
wire v$G6_680_out0;
wire v$G6_681_out0;
wire v$G6_682_out0;
wire v$G6_683_out0;
wire v$G6_684_out0;
wire v$G6_685_out0;
wire v$G6_686_out0;
wire v$G6_687_out0;
wire v$G6_688_out0;
wire v$G6_689_out0;
wire v$G6_690_out0;
wire v$G6_691_out0;
wire v$G6_692_out0;
wire v$G6_693_out0;
wire v$G6_694_out0;
wire v$G6_695_out0;
wire v$G6_696_out0;
wire v$G6_697_out0;
wire v$G6_730_out0;
wire v$G6_731_out0;
wire v$G6_7798_out0;
wire v$G6_7799_out0;
wire v$G6_8265_out0;
wire v$G6_8266_out0;
wire v$G6_9404_out0;
wire v$G6_9405_out0;
wire v$G70_10735_out0;
wire v$G70_10736_out0;
wire v$G70_14638_out0;
wire v$G71_15857_out0;
wire v$G71_15858_out0;
wire v$G72_6179_out0;
wire v$G74_16338_out0;
wire v$G77_18811_out0;
wire v$G78_7386_out0;
wire v$G79_13307_out0;
wire v$G7_10017_out0;
wire v$G7_10018_out0;
wire v$G7_10019_out0;
wire v$G7_10020_out0;
wire v$G7_10021_out0;
wire v$G7_10022_out0;
wire v$G7_10023_out0;
wire v$G7_10024_out0;
wire v$G7_10025_out0;
wire v$G7_10026_out0;
wire v$G7_10027_out0;
wire v$G7_10028_out0;
wire v$G7_10029_out0;
wire v$G7_10030_out0;
wire v$G7_10031_out0;
wire v$G7_10032_out0;
wire v$G7_10033_out0;
wire v$G7_10034_out0;
wire v$G7_10035_out0;
wire v$G7_10036_out0;
wire v$G7_10037_out0;
wire v$G7_10038_out0;
wire v$G7_10039_out0;
wire v$G7_10040_out0;
wire v$G7_10041_out0;
wire v$G7_10042_out0;
wire v$G7_10043_out0;
wire v$G7_10044_out0;
wire v$G7_10045_out0;
wire v$G7_10046_out0;
wire v$G7_10047_out0;
wire v$G7_10048_out0;
wire v$G7_10049_out0;
wire v$G7_10050_out0;
wire v$G7_10051_out0;
wire v$G7_10052_out0;
wire v$G7_10053_out0;
wire v$G7_10054_out0;
wire v$G7_10055_out0;
wire v$G7_10056_out0;
wire v$G7_10057_out0;
wire v$G7_10058_out0;
wire v$G7_10059_out0;
wire v$G7_10060_out0;
wire v$G7_10061_out0;
wire v$G7_10062_out0;
wire v$G7_10063_out0;
wire v$G7_10064_out0;
wire v$G7_10065_out0;
wire v$G7_10066_out0;
wire v$G7_10067_out0;
wire v$G7_10068_out0;
wire v$G7_10069_out0;
wire v$G7_10070_out0;
wire v$G7_10071_out0;
wire v$G7_10072_out0;
wire v$G7_10073_out0;
wire v$G7_10074_out0;
wire v$G7_10075_out0;
wire v$G7_10076_out0;
wire v$G7_10077_out0;
wire v$G7_10078_out0;
wire v$G7_10079_out0;
wire v$G7_10080_out0;
wire v$G7_10081_out0;
wire v$G7_10082_out0;
wire v$G7_10083_out0;
wire v$G7_10084_out0;
wire v$G7_10085_out0;
wire v$G7_10086_out0;
wire v$G7_10087_out0;
wire v$G7_10088_out0;
wire v$G7_10089_out0;
wire v$G7_10090_out0;
wire v$G7_10091_out0;
wire v$G7_10092_out0;
wire v$G7_10093_out0;
wire v$G7_10094_out0;
wire v$G7_10095_out0;
wire v$G7_10096_out0;
wire v$G7_10097_out0;
wire v$G7_10098_out0;
wire v$G7_10099_out0;
wire v$G7_10100_out0;
wire v$G7_10101_out0;
wire v$G7_10102_out0;
wire v$G7_10103_out0;
wire v$G7_10104_out0;
wire v$G7_10105_out0;
wire v$G7_10106_out0;
wire v$G7_10107_out0;
wire v$G7_10108_out0;
wire v$G7_10109_out0;
wire v$G7_10110_out0;
wire v$G7_10111_out0;
wire v$G7_10112_out0;
wire v$G7_10113_out0;
wire v$G7_10114_out0;
wire v$G7_10115_out0;
wire v$G7_10116_out0;
wire v$G7_10117_out0;
wire v$G7_10118_out0;
wire v$G7_10119_out0;
wire v$G7_10120_out0;
wire v$G7_10121_out0;
wire v$G7_10122_out0;
wire v$G7_10123_out0;
wire v$G7_10124_out0;
wire v$G7_10125_out0;
wire v$G7_10126_out0;
wire v$G7_10127_out0;
wire v$G7_10128_out0;
wire v$G7_10129_out0;
wire v$G7_10130_out0;
wire v$G7_10131_out0;
wire v$G7_10132_out0;
wire v$G7_10133_out0;
wire v$G7_10134_out0;
wire v$G7_10135_out0;
wire v$G7_10136_out0;
wire v$G7_10137_out0;
wire v$G7_10138_out0;
wire v$G7_10139_out0;
wire v$G7_10140_out0;
wire v$G7_10141_out0;
wire v$G7_10142_out0;
wire v$G7_10143_out0;
wire v$G7_10144_out0;
wire v$G7_10145_out0;
wire v$G7_10146_out0;
wire v$G7_10147_out0;
wire v$G7_10148_out0;
wire v$G7_10149_out0;
wire v$G7_10150_out0;
wire v$G7_10151_out0;
wire v$G7_10152_out0;
wire v$G7_10153_out0;
wire v$G7_10154_out0;
wire v$G7_10155_out0;
wire v$G7_10156_out0;
wire v$G7_10157_out0;
wire v$G7_10158_out0;
wire v$G7_10159_out0;
wire v$G7_10160_out0;
wire v$G7_10161_out0;
wire v$G7_10162_out0;
wire v$G7_10163_out0;
wire v$G7_10164_out0;
wire v$G7_10165_out0;
wire v$G7_10166_out0;
wire v$G7_10167_out0;
wire v$G7_10168_out0;
wire v$G7_10169_out0;
wire v$G7_10170_out0;
wire v$G7_10171_out0;
wire v$G7_10172_out0;
wire v$G7_10173_out0;
wire v$G7_10174_out0;
wire v$G7_10175_out0;
wire v$G7_10176_out0;
wire v$G7_10177_out0;
wire v$G7_10178_out0;
wire v$G7_10179_out0;
wire v$G7_10180_out0;
wire v$G7_10181_out0;
wire v$G7_10182_out0;
wire v$G7_10183_out0;
wire v$G7_10184_out0;
wire v$G7_10185_out0;
wire v$G7_10186_out0;
wire v$G7_10187_out0;
wire v$G7_10188_out0;
wire v$G7_10189_out0;
wire v$G7_10190_out0;
wire v$G7_10191_out0;
wire v$G7_10192_out0;
wire v$G7_10193_out0;
wire v$G7_10194_out0;
wire v$G7_10195_out0;
wire v$G7_10196_out0;
wire v$G7_10197_out0;
wire v$G7_10198_out0;
wire v$G7_10199_out0;
wire v$G7_10200_out0;
wire v$G7_10201_out0;
wire v$G7_10202_out0;
wire v$G7_10203_out0;
wire v$G7_10204_out0;
wire v$G7_10205_out0;
wire v$G7_10206_out0;
wire v$G7_10207_out0;
wire v$G7_10208_out0;
wire v$G7_10209_out0;
wire v$G7_10210_out0;
wire v$G7_10211_out0;
wire v$G7_10212_out0;
wire v$G7_10213_out0;
wire v$G7_10214_out0;
wire v$G7_10215_out0;
wire v$G7_10216_out0;
wire v$G7_10217_out0;
wire v$G7_10218_out0;
wire v$G7_10219_out0;
wire v$G7_10220_out0;
wire v$G7_10221_out0;
wire v$G7_10222_out0;
wire v$G7_10223_out0;
wire v$G7_10224_out0;
wire v$G7_10225_out0;
wire v$G7_10226_out0;
wire v$G7_10227_out0;
wire v$G7_10228_out0;
wire v$G7_10229_out0;
wire v$G7_10230_out0;
wire v$G7_10231_out0;
wire v$G7_10232_out0;
wire v$G7_10233_out0;
wire v$G7_10234_out0;
wire v$G7_10235_out0;
wire v$G7_10236_out0;
wire v$G7_10237_out0;
wire v$G7_10238_out0;
wire v$G7_10239_out0;
wire v$G7_10240_out0;
wire v$G7_10241_out0;
wire v$G7_10242_out0;
wire v$G7_10243_out0;
wire v$G7_10244_out0;
wire v$G7_10245_out0;
wire v$G7_10246_out0;
wire v$G7_10247_out0;
wire v$G7_10248_out0;
wire v$G7_10249_out0;
wire v$G7_10250_out0;
wire v$G7_10251_out0;
wire v$G7_10252_out0;
wire v$G7_10253_out0;
wire v$G7_10254_out0;
wire v$G7_10255_out0;
wire v$G7_10256_out0;
wire v$G7_10257_out0;
wire v$G7_10258_out0;
wire v$G7_10259_out0;
wire v$G7_10260_out0;
wire v$G7_10261_out0;
wire v$G7_10262_out0;
wire v$G7_10275_out0;
wire v$G7_10276_out0;
wire v$G7_10277_out0;
wire v$G7_10278_out0;
wire v$G7_10295_out0;
wire v$G7_10362_out0;
wire v$G7_10363_out0;
wire v$G7_11473_out0;
wire v$G7_11474_out0;
wire v$G7_12368_out0;
wire v$G7_12369_out0;
wire v$G7_12768_out0;
wire v$G7_12769_out0;
wire v$G7_13231_out0;
wire v$G7_13232_out0;
wire v$G7_14015_out0;
wire v$G7_14016_out0;
wire v$G7_14136_out0;
wire v$G7_14137_out0;
wire v$G7_14734_out0;
wire v$G7_14735_out0;
wire v$G7_14736_out0;
wire v$G7_14737_out0;
wire v$G7_14738_out0;
wire v$G7_14739_out0;
wire v$G7_14740_out0;
wire v$G7_14741_out0;
wire v$G7_14742_out0;
wire v$G7_14743_out0;
wire v$G7_14744_out0;
wire v$G7_14745_out0;
wire v$G7_14914_out0;
wire v$G7_14915_out0;
wire v$G7_15277_out0;
wire v$G7_15278_out0;
wire v$G7_15414_out0;
wire v$G7_1653_out0;
wire v$G7_1654_out0;
wire v$G7_18265_out0;
wire v$G7_1849_out0;
wire v$G7_1850_out0;
wire v$G7_1851_out0;
wire v$G7_1852_out0;
wire v$G7_1853_out0;
wire v$G7_1854_out0;
wire v$G7_18741_out0;
wire v$G7_18742_out0;
wire v$G7_18743_out0;
wire v$G7_18744_out0;
wire v$G7_18745_out0;
wire v$G7_18746_out0;
wire v$G7_18747_out0;
wire v$G7_18748_out0;
wire v$G7_18749_out0;
wire v$G7_18750_out0;
wire v$G7_18751_out0;
wire v$G7_18752_out0;
wire v$G7_18753_out0;
wire v$G7_18754_out0;
wire v$G7_18755_out0;
wire v$G7_18756_out0;
wire v$G7_18757_out0;
wire v$G7_18758_out0;
wire v$G7_18759_out0;
wire v$G7_18760_out0;
wire v$G7_18761_out0;
wire v$G7_18762_out0;
wire v$G7_18763_out0;
wire v$G7_18764_out0;
wire v$G7_18765_out0;
wire v$G7_18766_out0;
wire v$G7_18767_out0;
wire v$G7_18768_out0;
wire v$G7_18769_out0;
wire v$G7_18770_out0;
wire v$G7_18771_out0;
wire v$G7_18772_out0;
wire v$G7_18773_out0;
wire v$G7_18774_out0;
wire v$G7_18775_out0;
wire v$G7_18776_out0;
wire v$G7_19251_out0;
wire v$G7_19252_out0;
wire v$G7_1991_out0;
wire v$G7_1992_out0;
wire v$G7_2442_out0;
wire v$G7_2443_out0;
wire v$G7_2444_out0;
wire v$G7_2445_out0;
wire v$G7_3377_out0;
wire v$G7_3378_out0;
wire v$G7_8043_out0;
wire v$G7_8044_out0;
wire v$G7_8168_out0;
wire v$G7_8169_out0;
wire v$G83_447_out0;
wire v$G84_1386_out0;
wire v$G85_6462_out0;
wire v$G86_14102_out0;
wire v$G87_5362_out0;
wire v$G88_7716_out0;
wire v$G89_18384_out0;
wire v$G8_11581_out0;
wire v$G8_11582_out0;
wire v$G8_11925_out0;
wire v$G8_11926_out0;
wire v$G8_11927_out0;
wire v$G8_11928_out0;
wire v$G8_11929_out0;
wire v$G8_11930_out0;
wire v$G8_11931_out0;
wire v$G8_11932_out0;
wire v$G8_11933_out0;
wire v$G8_11934_out0;
wire v$G8_11935_out0;
wire v$G8_11936_out0;
wire v$G8_11937_out0;
wire v$G8_11938_out0;
wire v$G8_11939_out0;
wire v$G8_11940_out0;
wire v$G8_11941_out0;
wire v$G8_11942_out0;
wire v$G8_11943_out0;
wire v$G8_11944_out0;
wire v$G8_11945_out0;
wire v$G8_11946_out0;
wire v$G8_11947_out0;
wire v$G8_11948_out0;
wire v$G8_11949_out0;
wire v$G8_11950_out0;
wire v$G8_11951_out0;
wire v$G8_11952_out0;
wire v$G8_11953_out0;
wire v$G8_11954_out0;
wire v$G8_11955_out0;
wire v$G8_11956_out0;
wire v$G8_11957_out0;
wire v$G8_11958_out0;
wire v$G8_11959_out0;
wire v$G8_11960_out0;
wire v$G8_11961_out0;
wire v$G8_11962_out0;
wire v$G8_11963_out0;
wire v$G8_11964_out0;
wire v$G8_11965_out0;
wire v$G8_11966_out0;
wire v$G8_11967_out0;
wire v$G8_11968_out0;
wire v$G8_11969_out0;
wire v$G8_11970_out0;
wire v$G8_11971_out0;
wire v$G8_11972_out0;
wire v$G8_11973_out0;
wire v$G8_11974_out0;
wire v$G8_11975_out0;
wire v$G8_11976_out0;
wire v$G8_11977_out0;
wire v$G8_11978_out0;
wire v$G8_11979_out0;
wire v$G8_11980_out0;
wire v$G8_11981_out0;
wire v$G8_11982_out0;
wire v$G8_11983_out0;
wire v$G8_11984_out0;
wire v$G8_11985_out0;
wire v$G8_11986_out0;
wire v$G8_11987_out0;
wire v$G8_11988_out0;
wire v$G8_11989_out0;
wire v$G8_11990_out0;
wire v$G8_11991_out0;
wire v$G8_11992_out0;
wire v$G8_11993_out0;
wire v$G8_11994_out0;
wire v$G8_11995_out0;
wire v$G8_11996_out0;
wire v$G8_11997_out0;
wire v$G8_11998_out0;
wire v$G8_11999_out0;
wire v$G8_12000_out0;
wire v$G8_12001_out0;
wire v$G8_12002_out0;
wire v$G8_12003_out0;
wire v$G8_12004_out0;
wire v$G8_12005_out0;
wire v$G8_12006_out0;
wire v$G8_12007_out0;
wire v$G8_12008_out0;
wire v$G8_12009_out0;
wire v$G8_12010_out0;
wire v$G8_12011_out0;
wire v$G8_12012_out0;
wire v$G8_12013_out0;
wire v$G8_12014_out0;
wire v$G8_12015_out0;
wire v$G8_12016_out0;
wire v$G8_12017_out0;
wire v$G8_12018_out0;
wire v$G8_12019_out0;
wire v$G8_12020_out0;
wire v$G8_12021_out0;
wire v$G8_12022_out0;
wire v$G8_12023_out0;
wire v$G8_12024_out0;
wire v$G8_12025_out0;
wire v$G8_12026_out0;
wire v$G8_12027_out0;
wire v$G8_12028_out0;
wire v$G8_12029_out0;
wire v$G8_12030_out0;
wire v$G8_12031_out0;
wire v$G8_12032_out0;
wire v$G8_12033_out0;
wire v$G8_12034_out0;
wire v$G8_12035_out0;
wire v$G8_12036_out0;
wire v$G8_12037_out0;
wire v$G8_12038_out0;
wire v$G8_12039_out0;
wire v$G8_12040_out0;
wire v$G8_12041_out0;
wire v$G8_12042_out0;
wire v$G8_12043_out0;
wire v$G8_12044_out0;
wire v$G8_12045_out0;
wire v$G8_12046_out0;
wire v$G8_12047_out0;
wire v$G8_12048_out0;
wire v$G8_12049_out0;
wire v$G8_12050_out0;
wire v$G8_12051_out0;
wire v$G8_12052_out0;
wire v$G8_12053_out0;
wire v$G8_12054_out0;
wire v$G8_12055_out0;
wire v$G8_12056_out0;
wire v$G8_12057_out0;
wire v$G8_12058_out0;
wire v$G8_12059_out0;
wire v$G8_12060_out0;
wire v$G8_12061_out0;
wire v$G8_12062_out0;
wire v$G8_12063_out0;
wire v$G8_12064_out0;
wire v$G8_12065_out0;
wire v$G8_12066_out0;
wire v$G8_12067_out0;
wire v$G8_12068_out0;
wire v$G8_12069_out0;
wire v$G8_12070_out0;
wire v$G8_12071_out0;
wire v$G8_12072_out0;
wire v$G8_12073_out0;
wire v$G8_12074_out0;
wire v$G8_12075_out0;
wire v$G8_12076_out0;
wire v$G8_12077_out0;
wire v$G8_12078_out0;
wire v$G8_12079_out0;
wire v$G8_12080_out0;
wire v$G8_12081_out0;
wire v$G8_12082_out0;
wire v$G8_12083_out0;
wire v$G8_12084_out0;
wire v$G8_12085_out0;
wire v$G8_12086_out0;
wire v$G8_12087_out0;
wire v$G8_12088_out0;
wire v$G8_12089_out0;
wire v$G8_12090_out0;
wire v$G8_12091_out0;
wire v$G8_12092_out0;
wire v$G8_12093_out0;
wire v$G8_12094_out0;
wire v$G8_12095_out0;
wire v$G8_12096_out0;
wire v$G8_12097_out0;
wire v$G8_12098_out0;
wire v$G8_12099_out0;
wire v$G8_12100_out0;
wire v$G8_12101_out0;
wire v$G8_12102_out0;
wire v$G8_12103_out0;
wire v$G8_12104_out0;
wire v$G8_12105_out0;
wire v$G8_12106_out0;
wire v$G8_12107_out0;
wire v$G8_12108_out0;
wire v$G8_12109_out0;
wire v$G8_12110_out0;
wire v$G8_12111_out0;
wire v$G8_12112_out0;
wire v$G8_12113_out0;
wire v$G8_12114_out0;
wire v$G8_12115_out0;
wire v$G8_12116_out0;
wire v$G8_12117_out0;
wire v$G8_12118_out0;
wire v$G8_12119_out0;
wire v$G8_12120_out0;
wire v$G8_12121_out0;
wire v$G8_12122_out0;
wire v$G8_12123_out0;
wire v$G8_12124_out0;
wire v$G8_12125_out0;
wire v$G8_12126_out0;
wire v$G8_12127_out0;
wire v$G8_12128_out0;
wire v$G8_12129_out0;
wire v$G8_12130_out0;
wire v$G8_12131_out0;
wire v$G8_12132_out0;
wire v$G8_12133_out0;
wire v$G8_12134_out0;
wire v$G8_12135_out0;
wire v$G8_12136_out0;
wire v$G8_12137_out0;
wire v$G8_12138_out0;
wire v$G8_12139_out0;
wire v$G8_12140_out0;
wire v$G8_12141_out0;
wire v$G8_12142_out0;
wire v$G8_12143_out0;
wire v$G8_12144_out0;
wire v$G8_12145_out0;
wire v$G8_12146_out0;
wire v$G8_12147_out0;
wire v$G8_12148_out0;
wire v$G8_12149_out0;
wire v$G8_12150_out0;
wire v$G8_12151_out0;
wire v$G8_12152_out0;
wire v$G8_12153_out0;
wire v$G8_12154_out0;
wire v$G8_12155_out0;
wire v$G8_12156_out0;
wire v$G8_12157_out0;
wire v$G8_12158_out0;
wire v$G8_12159_out0;
wire v$G8_12160_out0;
wire v$G8_12161_out0;
wire v$G8_12162_out0;
wire v$G8_12163_out0;
wire v$G8_12164_out0;
wire v$G8_12165_out0;
wire v$G8_12166_out0;
wire v$G8_12167_out0;
wire v$G8_12168_out0;
wire v$G8_12169_out0;
wire v$G8_12170_out0;
wire v$G8_12567_out0;
wire v$G8_12568_out0;
wire v$G8_12569_out0;
wire v$G8_12570_out0;
wire v$G8_12571_out0;
wire v$G8_12572_out0;
wire v$G8_12573_out0;
wire v$G8_12574_out0;
wire v$G8_12575_out0;
wire v$G8_12576_out0;
wire v$G8_12577_out0;
wire v$G8_12578_out0;
wire v$G8_12579_out0;
wire v$G8_12580_out0;
wire v$G8_12581_out0;
wire v$G8_12582_out0;
wire v$G8_12583_out0;
wire v$G8_12584_out0;
wire v$G8_12585_out0;
wire v$G8_12586_out0;
wire v$G8_12587_out0;
wire v$G8_12588_out0;
wire v$G8_12589_out0;
wire v$G8_12590_out0;
wire v$G8_12591_out0;
wire v$G8_12592_out0;
wire v$G8_12593_out0;
wire v$G8_12594_out0;
wire v$G8_12595_out0;
wire v$G8_12596_out0;
wire v$G8_12597_out0;
wire v$G8_12598_out0;
wire v$G8_12599_out0;
wire v$G8_12600_out0;
wire v$G8_12601_out0;
wire v$G8_12602_out0;
wire v$G8_12863_out0;
wire v$G8_12864_out0;
wire v$G8_13076_out0;
wire v$G8_13077_out0;
wire v$G8_13988_out0;
wire v$G8_13989_out0;
wire v$G8_1401_out0;
wire v$G8_1402_out0;
wire v$G8_14859_out0;
wire v$G8_14860_out0;
wire v$G8_14861_out0;
wire v$G8_14862_out0;
wire v$G8_14863_out0;
wire v$G8_14864_out0;
wire v$G8_14865_out0;
wire v$G8_14866_out0;
wire v$G8_14867_out0;
wire v$G8_14868_out0;
wire v$G8_14869_out0;
wire v$G8_14870_out0;
wire v$G8_16068_out0;
wire v$G8_16069_out0;
wire v$G8_16329_out0;
wire v$G8_18510_out0;
wire v$G8_18511_out0;
wire v$G8_19390_out0;
wire v$G8_19391_out0;
wire v$G8_2050_out0;
wire v$G8_2051_out0;
wire v$G8_2052_out0;
wire v$G8_2053_out0;
wire v$G8_2054_out0;
wire v$G8_2055_out0;
wire v$G8_2056_out0;
wire v$G8_2057_out0;
wire v$G8_2448_out0;
wire v$G8_2449_out0;
wire v$G8_2473_out0;
wire v$G8_2474_out0;
wire v$G8_255_out0;
wire v$G8_256_out0;
wire v$G8_2607_out0;
wire v$G8_2608_out0;
wire v$G8_2770_out0;
wire v$G8_2771_out0;
wire v$G8_2772_out0;
wire v$G8_2773_out0;
wire v$G8_2774_out0;
wire v$G8_2775_out0;
wire v$G8_3907_out0;
wire v$G8_3908_out0;
wire v$G8_3909_out0;
wire v$G8_3910_out0;
wire v$G8_3911_out0;
wire v$G8_3912_out0;
wire v$G8_3913_out0;
wire v$G8_3914_out0;
wire v$G8_3915_out0;
wire v$G8_3916_out0;
wire v$G8_3917_out0;
wire v$G8_3918_out0;
wire v$G8_3919_out0;
wire v$G8_3920_out0;
wire v$G8_3921_out0;
wire v$G8_3922_out0;
wire v$G8_3923_out0;
wire v$G8_3924_out0;
wire v$G8_3925_out0;
wire v$G8_3926_out0;
wire v$G8_3927_out0;
wire v$G8_3928_out0;
wire v$G8_3929_out0;
wire v$G8_3930_out0;
wire v$G8_5032_out0;
wire v$G8_5033_out0;
wire v$G8_6328_out0;
wire v$G8_6329_out0;
wire v$G8_6340_out0;
wire v$G8_6341_out0;
wire v$G8_9410_out0;
wire v$G8_9411_out0;
wire v$G8_9881_out0;
wire v$G8_9882_out0;
wire v$G90_8368_out0;
wire v$G9_1331_out0;
wire v$G9_1332_out0;
wire v$G9_14031_out0;
wire v$G9_14032_out0;
wire v$G9_15733_out0;
wire v$G9_15734_out0;
wire v$G9_15797_out0;
wire v$G9_15798_out0;
wire v$G9_15799_out0;
wire v$G9_15800_out0;
wire v$G9_15801_out0;
wire v$G9_15802_out0;
wire v$G9_15803_out0;
wire v$G9_15804_out0;
wire v$G9_16121_out0;
wire v$G9_16122_out0;
wire v$G9_16183_out0;
wire v$G9_16184_out0;
wire v$G9_16651_out0;
wire v$G9_16652_out0;
wire v$G9_17120_out0;
wire v$G9_17121_out0;
wire v$G9_17527_out0;
wire v$G9_17528_out0;
wire v$G9_17559_out0;
wire v$G9_17560_out0;
wire v$G9_17602_out0;
wire v$G9_17603_out0;
wire v$G9_18211_out0;
wire v$G9_18212_out0;
wire v$G9_18213_out0;
wire v$G9_18214_out0;
wire v$G9_18215_out0;
wire v$G9_18216_out0;
wire v$G9_18217_out0;
wire v$G9_18218_out0;
wire v$G9_18219_out0;
wire v$G9_18220_out0;
wire v$G9_18221_out0;
wire v$G9_18222_out0;
wire v$G9_18223_out0;
wire v$G9_18224_out0;
wire v$G9_18225_out0;
wire v$G9_18226_out0;
wire v$G9_18227_out0;
wire v$G9_18228_out0;
wire v$G9_18229_out0;
wire v$G9_18230_out0;
wire v$G9_18231_out0;
wire v$G9_18232_out0;
wire v$G9_18233_out0;
wire v$G9_18234_out0;
wire v$G9_18235_out0;
wire v$G9_18236_out0;
wire v$G9_18237_out0;
wire v$G9_18238_out0;
wire v$G9_18239_out0;
wire v$G9_18240_out0;
wire v$G9_18241_out0;
wire v$G9_18242_out0;
wire v$G9_18243_out0;
wire v$G9_18244_out0;
wire v$G9_18245_out0;
wire v$G9_18246_out0;
wire v$G9_18316_out0;
wire v$G9_18317_out0;
wire v$G9_2724_out0;
wire v$G9_2725_out0;
wire v$G9_3651_out0;
wire v$G9_3652_out0;
wire v$G9_6085_out0;
wire v$G9_6086_out0;
wire v$G9_6490_out0;
wire v$G9_6491_out0;
wire v$G9_6588_out0;
wire v$G9_6589_out0;
wire v$G9_9018_out0;
wire v$G9_9019_out0;
wire v$G9_9255_out0;
wire v$G9_9256_out0;
wire v$G9_9257_out0;
wire v$G9_9258_out0;
wire v$G9_9259_out0;
wire v$G9_9260_out0;
wire v$GATE1_720_out0;
wire v$GATE1_721_out0;
wire v$GATE1_722_out0;
wire v$GATE1_723_out0;
wire v$GATE1_724_out0;
wire v$GATE1_725_out0;
wire v$GATE2_16355_out0;
wire v$GATE2_16356_out0;
wire v$GATE2_16357_out0;
wire v$GATE2_16358_out0;
wire v$GATE2_16359_out0;
wire v$GATE2_16360_out0;
wire v$G_10482_out0;
wire v$G_10483_out0;
wire v$G_10484_out0;
wire v$G_10485_out0;
wire v$G_10486_out0;
wire v$G_10487_out0;
wire v$G_10488_out0;
wire v$G_10489_out0;
wire v$G_10490_out0;
wire v$G_10491_out0;
wire v$G_10492_out0;
wire v$G_10493_out0;
wire v$G_10494_out0;
wire v$G_10495_out0;
wire v$G_10496_out0;
wire v$G_10497_out0;
wire v$G_10498_out0;
wire v$G_10499_out0;
wire v$G_10500_out0;
wire v$G_10501_out0;
wire v$G_10502_out0;
wire v$G_10503_out0;
wire v$G_10504_out0;
wire v$G_10505_out0;
wire v$G_10506_out0;
wire v$G_10507_out0;
wire v$G_10508_out0;
wire v$G_10509_out0;
wire v$G_10510_out0;
wire v$G_10511_out0;
wire v$G_10512_out0;
wire v$G_10513_out0;
wire v$G_10514_out0;
wire v$G_10515_out0;
wire v$G_10516_out0;
wire v$G_10517_out0;
wire v$G_10518_out0;
wire v$G_10519_out0;
wire v$G_10520_out0;
wire v$G_10521_out0;
wire v$G_10522_out0;
wire v$G_10523_out0;
wire v$G_10524_out0;
wire v$G_10525_out0;
wire v$G_10526_out0;
wire v$G_10527_out0;
wire v$G_10528_out0;
wire v$G_10529_out0;
wire v$G_10530_out0;
wire v$G_10531_out0;
wire v$G_10532_out0;
wire v$G_10533_out0;
wire v$G_10534_out0;
wire v$G_10535_out0;
wire v$G_10536_out0;
wire v$G_10537_out0;
wire v$G_10538_out0;
wire v$G_10539_out0;
wire v$G_10540_out0;
wire v$G_10541_out0;
wire v$G_10542_out0;
wire v$G_10543_out0;
wire v$G_10544_out0;
wire v$G_10545_out0;
wire v$G_10546_out0;
wire v$G_10547_out0;
wire v$G_10548_out0;
wire v$G_10549_out0;
wire v$G_10550_out0;
wire v$G_10551_out0;
wire v$G_10552_out0;
wire v$G_10553_out0;
wire v$G_10554_out0;
wire v$G_10555_out0;
wire v$G_10556_out0;
wire v$G_10557_out0;
wire v$G_10558_out0;
wire v$G_10559_out0;
wire v$G_10560_out0;
wire v$G_10561_out0;
wire v$G_10562_out0;
wire v$G_10563_out0;
wire v$G_10564_out0;
wire v$G_10565_out0;
wire v$G_10566_out0;
wire v$G_10567_out0;
wire v$G_10568_out0;
wire v$G_10569_out0;
wire v$G_10570_out0;
wire v$G_10571_out0;
wire v$G_10572_out0;
wire v$G_10573_out0;
wire v$G_10574_out0;
wire v$G_10575_out0;
wire v$G_10576_out0;
wire v$G_10577_out0;
wire v$G_10578_out0;
wire v$G_10579_out0;
wire v$G_10580_out0;
wire v$G_10581_out0;
wire v$G_10582_out0;
wire v$G_10583_out0;
wire v$G_10584_out0;
wire v$G_10585_out0;
wire v$G_10586_out0;
wire v$G_10587_out0;
wire v$G_10588_out0;
wire v$G_10589_out0;
wire v$G_10590_out0;
wire v$G_10591_out0;
wire v$G_10592_out0;
wire v$G_10593_out0;
wire v$G_10594_out0;
wire v$G_10595_out0;
wire v$G_10596_out0;
wire v$G_10597_out0;
wire v$G_10598_out0;
wire v$G_10599_out0;
wire v$G_10600_out0;
wire v$G_10601_out0;
wire v$G_10602_out0;
wire v$G_10603_out0;
wire v$G_10604_out0;
wire v$G_10605_out0;
wire v$G_10606_out0;
wire v$G_10607_out0;
wire v$G_10608_out0;
wire v$G_10609_out0;
wire v$G_10610_out0;
wire v$G_10611_out0;
wire v$G_10612_out0;
wire v$G_10613_out0;
wire v$G_10614_out0;
wire v$G_10615_out0;
wire v$G_10616_out0;
wire v$G_10617_out0;
wire v$G_10618_out0;
wire v$G_10619_out0;
wire v$G_10620_out0;
wire v$G_10621_out0;
wire v$G_10622_out0;
wire v$G_10623_out0;
wire v$G_10624_out0;
wire v$G_10625_out0;
wire v$HALT$PREV$PREV$PREV_8049_out0;
wire v$HALT$PREV$PREV$PREV_8050_out0;
wire v$HALT$PREV$PREV_18681_out0;
wire v$HALT$PREV$PREV_18682_out0;
wire v$HALT$PREV_10837_out0;
wire v$HALT$PREV_10838_out0;
wire v$HALT0_12252_out0;
wire v$HALT0_14750_out0;
wire v$HALT0_380_out0;
wire v$HALT0_6091_out0;
wire v$HALT1_18913_out0;
wire v$HALT1_3317_out0;
wire v$HALT1_4317_out0;
wire v$HALT1_7543_out0;
wire v$HALTED_12399_out0;
wire v$HALTED_12400_out0;
wire v$HALTSEL_15349_out0;
wire v$HALTVALID_13870_out0;
wire v$HALTVALID_8061_out0;
wire v$HALT_13471_out0;
wire v$HALT_13472_out0;
wire v$HALT_1449_out0;
wire v$HALT_16989_out0;
wire v$HALT_18283_out0;
wire v$HALT_18284_out0;
wire v$HALT_3106_out0;
wire v$HALT_3107_out0;
wire v$HALT_7897_out0;
wire v$HALT_7898_out0;
wire v$HIGHER$OUT_4011_out0;
wire v$HIGHER$OUT_4012_out0;
wire v$HIGHER$OUT_4013_out0;
wire v$HIGHER$OUT_4014_out0;
wire v$HIGHER$OUT_4015_out0;
wire v$HIGHER$OUT_4016_out0;
wire v$HIGHER$OUT_4017_out0;
wire v$HIGHER$OUT_4018_out0;
wire v$HIGHER$OUT_8106_out0;
wire v$HIGHER$OUT_8107_out0;
wire v$HIGHER$OUT_8108_out0;
wire v$HIGHER$OUT_8109_out0;
wire v$HIGHER$SAME_15638_out0;
wire v$HIGHER$SAME_15639_out0;
wire v$HIGHER$SAME_15640_out0;
wire v$HIGHER$SAME_15641_out0;
wire v$HIGHER$SAME_15642_out0;
wire v$HIGHER$SAME_15643_out0;
wire v$HIGHER$SAME_15644_out0;
wire v$HIGHER$SAME_15645_out0;
wire v$HIGHER$SAME_9460_out0;
wire v$HIGHER$SAME_9461_out0;
wire v$HIGHER$SAME_9462_out0;
wire v$HIGHER$SAME_9463_out0;
wire v$I0EN_8356_out0;
wire v$I0EN_8357_out0;
wire v$I0P_10763_out0;
wire v$I0P_10764_out0;
wire v$I0P_2632_out0;
wire v$I0P_2633_out0;
wire v$I0P_4512_out0;
wire v$I0P_4513_out0;
wire v$I0REGISTERWRITE_3578_out0;
wire v$I0REGISTERWRITE_3579_out0;
wire v$I0_19117_out0;
wire v$I0_19118_out0;
wire v$I1EN_19009_out0;
wire v$I1EN_19010_out0;
wire v$I1P_15425_out0;
wire v$I1P_15426_out0;
wire v$I1P_2710_out0;
wire v$I1P_2711_out0;
wire v$I1P_6684_out0;
wire v$I1P_6685_out0;
wire v$I1REGISTERWRITE_3139_out0;
wire v$I1REGISTERWRITE_3140_out0;
wire v$I1_5106_out0;
wire v$I1_5107_out0;
wire v$I2EN_16345_out0;
wire v$I2EN_16346_out0;
wire v$I2P_2465_out0;
wire v$I2P_2466_out0;
wire v$I2P_6676_out0;
wire v$I2P_6677_out0;
wire v$I2P_7810_out0;
wire v$I2P_7811_out0;
wire v$I2REGISTERWRITE_12504_out0;
wire v$I2REGISTERWRITE_12505_out0;
wire v$I2_15092_out0;
wire v$I2_15093_out0;
wire v$I3EN_18387_out0;
wire v$I3EN_18388_out0;
wire v$I3P_11324_out0;
wire v$I3P_11325_out0;
wire v$I3P_14197_out0;
wire v$I3P_14198_out0;
wire v$I3P_9295_out0;
wire v$I3P_9296_out0;
wire v$I3REGISTERWRITE_1419_out0;
wire v$I3REGISTERWRITE_1420_out0;
wire v$I3_5036_out0;
wire v$I3_5037_out0;
wire v$IGNORE_12272_out0;
wire v$IGNORE_12273_out0;
wire v$IGNORE_17180_out0;
wire v$IGNORE_17181_out0;
wire v$IGNORE_5650_out0;
wire v$IGNORE_5651_out0;
wire v$IGNORE_8594_out0;
wire v$INCOMINGINTERRUPT_2066_out0;
wire v$INCOMINGINTERRUPT_2067_out0;
wire v$ININTERRUPT_1277_out0;
wire v$ININTERRUPT_1278_out0;
wire v$ININT_16052_out0;
wire v$ININT_16053_out0;
wire v$INITIAL$FETCH$OCCURRED_1691_out0;
wire v$INITIAL$FETCH$OCCURRED_1692_out0;
wire v$INIT_11241_out0;
wire v$INIT_11242_out0;
wire v$INT2_3379_out0;
wire v$INT2_3380_out0;
wire v$INT2_5648_out0;
wire v$INT2_5649_out0;
wire v$INT3_14645_out0;
wire v$INT3_14646_out0;
wire v$INT3_18737_out0;
wire v$INT3_18738_out0;
wire v$INTCAPTURE0_14107_out0;
wire v$INTCAPTURE0_14108_out0;
wire v$INTCLEAR_8096_out0;
wire v$INTCLEAR_8097_out0;
wire v$INTCLR_220_out0;
wire v$INTCLR_221_out0;
wire v$INTCOUNT_7792_out0;
wire v$INTCOUNT_7793_out0;
wire v$INTDISABLE_2882_out0;
wire v$INTDISABLE_2883_out0;
wire v$INTDISABLE_5214_out0;
wire v$INTDISABLE_5215_out0;
wire v$INTENABLE_18046_out0;
wire v$INTENABLE_18047_out0;
wire v$INTENABLE_3148_out0;
wire v$INTENABLE_3149_out0;
wire v$INTERRUPT0_12268_out0;
wire v$INTERRUPT0_12269_out0;
wire v$INTERRUPT0_1967_out0;
wire v$INTERRUPT0_1968_out0;
wire v$INTERRUPT1_18306_out0;
wire v$INTERRUPT1_18307_out0;
wire v$INTERRUPT1_8595_out0;
wire v$INTERRUPT1_8596_out0;
wire v$INTERRUPT2_1821_out0;
wire v$INTERRUPT2_1822_out0;
wire v$INTERRUPT2_4034_out0;
wire v$INTERRUPT2_4035_out0;
wire v$INTERRUPT3_3040_out0;
wire v$INTERRUPT3_3041_out0;
wire v$INTERRUPT3_3708_out0;
wire v$INTERRUPT3_3709_out0;
wire v$INTERRUPTOVERFLOW_15719_out0;
wire v$INTERRUPTOVERFLOW_15720_out0;
wire v$INTERRUPTOVERFLOW_2438_out0;
wire v$INTERRUPTOVERFLOW_2439_out0;
wire v$INTERRUPTSENABLED_10002_out0;
wire v$INTERRUPTSENABLED_10003_out0;
wire v$INTOVERFLOW_16653_out0;
wire v$INTOVERFLOW_16654_out0;
wire v$IR1$15_6043_out0;
wire v$IR1$15_6044_out0;
wire v$IR1$32$BITS_8191_out0;
wire v$IR1$32$BITS_8192_out0;
wire v$IR1$C$L_10480_out0;
wire v$IR1$C$L_10481_out0;
wire v$IR1$IS$FPU$ARITHMETIC_1533_out0;
wire v$IR1$IS$FPU$ARITHMETIC_1534_out0;
wire v$IR1$IS$FPU$LOAD$STORE_9261_out0;
wire v$IR1$IS$FPU$LOAD$STORE_9262_out0;
wire v$IR1$IS$LDST_13783_out0;
wire v$IR1$IS$LDST_13784_out0;
wire v$IR1$IS$STORE_4631_out0;
wire v$IR1$IS$STORE_4632_out0;
wire v$IR1$LS_17045_out0;
wire v$IR1$LS_17046_out0;
wire v$IR1$L_5356_out0;
wire v$IR1$L_5357_out0;
wire v$IR1$P_3871_out0;
wire v$IR1$P_3872_out0;
wire v$IR1$S$WB_336_out0;
wire v$IR1$S$WB_337_out0;
wire v$IR1$S_8164_out0;
wire v$IR1$S_8165_out0;
wire v$IR1$U_15384_out0;
wire v$IR1$U_15385_out0;
wire v$IR1$VALID$VIEWER_1769_out0;
wire v$IR1$VALID$VIEWER_1770_out0;
wire v$IR1$VALID_14622_out0;
wire v$IR1$VALID_14623_out0;
wire v$IR1$VALID_18403_out0;
wire v$IR1$VALID_18404_out0;
wire v$IR1$VALID_19035_out0;
wire v$IR1$VALID_19036_out0;
wire v$IR1$VALID_4028_out0;
wire v$IR1$VALID_4029_out0;
wire v$IR1$VALID_6037_out0;
wire v$IR1$VALID_6038_out0;
wire v$IR1$VALID_62_out0;
wire v$IR1$VALID_63_out0;
wire v$IR1$VALID_9829_out0;
wire v$IR1$VALID_9830_out0;
wire v$IR1$W_17168_out0;
wire v$IR1$W_17169_out0;
wire v$IR15_11184_out0;
wire v$IR15_11185_out0;
wire v$IR15_11494_out0;
wire v$IR15_11495_out0;
wire v$IR2$15_7754_out0;
wire v$IR2$15_7755_out0;
wire v$IR2$FPU$32BIT_12372_out0;
wire v$IR2$FPU$32BIT_12373_out0;
wire v$IR2$FPU$LOADA_15851_out0;
wire v$IR2$FPU$LOADA_15852_out0;
wire v$IR2$FPU$LOAD_4390_out0;
wire v$IR2$FPU$LOAD_4391_out0;
wire v$IR2$FPU$L_11232_out0;
wire v$IR2$FPU$L_11233_out0;
wire v$IR2$IS$FPU_12415_out0;
wire v$IR2$IS$FPU_12416_out0;
wire v$IR2$IS$FPU_3137_out0;
wire v$IR2$IS$FPU_3138_out0;
wire v$IR2$IS$FPU_7335_out0;
wire v$IR2$IS$FPU_7336_out0;
wire v$IR2$IS$LDST_4560_out0;
wire v$IR2$IS$LDST_4561_out0;
wire v$IR2$LS_16436_out0;
wire v$IR2$LS_16437_out0;
wire v$IR2$L_13058_out0;
wire v$IR2$L_13059_out0;
wire v$IR2$P_17955_out0;
wire v$IR2$P_17956_out0;
wire v$IR2$REG$IMMEDIATE_6456_out0;
wire v$IR2$REG$IMMEDIATE_6457_out0;
wire v$IR2$S$WB_18080_out0;
wire v$IR2$S$WB_18081_out0;
wire v$IR2$S_1315_out0;
wire v$IR2$S_1316_out0;
wire v$IR2$U_6182_out0;
wire v$IR2$U_6183_out0;
wire v$IR2$VALID$AND$NOT$FLOAD_5094_out0;
wire v$IR2$VALID$AND$NOT$FLOAD_5095_out0;
wire v$IR2$VALID$AND$NOT$FLOAD_7603_out0;
wire v$IR2$VALID$AND$NOT$FLOAD_7604_out0;
wire v$IR2$VALID$VIEWER_6087_out0;
wire v$IR2$VALID$VIEWER_6088_out0;
wire v$IR2$VALID_11160_out0;
wire v$IR2$VALID_11161_out0;
wire v$IR2$VALID_12366_out0;
wire v$IR2$VALID_12367_out0;
wire v$IR2$VALID_13833_out0;
wire v$IR2$VALID_13834_out0;
wire v$IR2$VALID_15430_out0;
wire v$IR2$VALID_15431_out0;
wire v$IR2$VALID_16482_out0;
wire v$IR2$VALID_16483_out0;
wire v$IR2$VALID_19367_out0;
wire v$IR2$VALID_19368_out0;
wire v$IR2$VALID_4376_out0;
wire v$IR2$VALID_4377_out0;
wire v$IR2$VALID_6701_out0;
wire v$IR2$VALID_6702_out0;
wire v$IR2$VALID_7739_out0;
wire v$IR2$VALID_7740_out0;
wire v$IR2$W_15717_out0;
wire v$IR2$W_15718_out0;
wire v$IS$32$BIT$FPU$ADDER_15580_out0;
wire v$IS$32$BIT$FPU$ADDER_15581_out0;
wire v$IS$32$BITS$VIEWER_1387_out0;
wire v$IS$32$BITS$VIEWER_1388_out0;
wire v$IS$32$BITS_14649_out0;
wire v$IS$32$BITS_14650_out0;
wire v$IS$32$BITS_18206_out0;
wire v$IS$32$BITS_18207_out0;
wire v$IS$32$BITS_3203_out0;
wire v$IS$32$BITS_3204_out0;
wire v$IS$32$BITS_4307_out0;
wire v$IS$32$BITS_4308_out0;
wire v$IS$32$BIT_11362_out0;
wire v$IS$32$BIT_11363_out0;
wire v$IS$32$BIT_11513_out0;
wire v$IS$32$BIT_11514_out0;
wire v$IS$A$LARGER_10896_out0;
wire v$IS$A$LARGER_10897_out0;
wire v$IS$A$LARGER_15264_out0;
wire v$IS$A$LARGER_15265_out0;
wire v$IS$A$LARGER_16598_out0;
wire v$IS$A$LARGER_16599_out0;
wire v$IS$A$LARGER_17444_out0;
wire v$IS$A$LARGER_17445_out0;
wire v$IS$A$LARGER_7361_out0;
wire v$IS$A$LARGER_7362_out0;
wire v$IS$FPU$HAZARD_358_out0;
wire v$IS$FPU$HAZARD_359_out0;
wire v$IS$IR1$FMUL_15879_out0;
wire v$IS$IR1$FMUL_15880_out0;
wire v$IS$IR1$FMUL_3174_out0;
wire v$IS$IR1$FMUL_3175_out0;
wire v$IS$IR2$DATA$PROCESSING_10368_out0;
wire v$IS$IR2$DATA$PROCESSING_10369_out0;
wire v$IS$SUB$MANTISA$ADDER_3389_out0;
wire v$IS$SUB$MANTISA$ADDER_3390_out0;
wire v$IS$SUB$VIEW_235_out0;
wire v$IS$SUB$VIEW_236_out0;
wire v$IS$SUB_13643_out0;
wire v$IS$SUB_13644_out0;
wire v$IS$SUB_16036_out0;
wire v$IS$SUB_16037_out0;
wire v$IS$SUB_4611_out0;
wire v$IS$SUB_4612_out0;
wire v$IS$SUM$0_1000_out0;
wire v$IS$SUM$0_1001_out0;
wire v$IS$SUM$0_16216_out0;
wire v$IS$SUM$0_16217_out0;
wire v$IS$SUM$0_16276_out0;
wire v$IS$SUM$0_16277_out0;
wire v$ISINTERRUPTED_12429_out0;
wire v$ISINTERRUPTED_12430_out0;
wire v$ISINTERRUPTED_12544_out0;
wire v$ISINTERRUPTED_12545_out0;
wire v$ISMOV_13213_out0;
wire v$ISMOV_13214_out0;
wire v$ISMOV_4234_out0;
wire v$ISMOV_4235_out0;
wire v$ISMOV_6907_out0;
wire v$ISMOV_6908_out0;
wire v$ISMOV_9117_out0;
wire v$ISMOV_9118_out0;
wire v$JEQ_1833_out0;
wire v$JEQ_1834_out0;
wire v$JEQ_18641_out0;
wire v$JEQ_18642_out0;
wire v$JLO_15598_out0;
wire v$JLO_15599_out0;
wire v$JLO_8424_out0;
wire v$JLO_8425_out0;
wire v$JLS_17065_out0;
wire v$JLS_17066_out0;
wire v$JLS_2120_out0;
wire v$JLS_2121_out0;
wire v$JMI_13727_out0;
wire v$JMI_13728_out0;
wire v$JMI_72_out0;
wire v$JMI_73_out0;
wire v$JMP_1825_out0;
wire v$JMP_1826_out0;
wire v$JMP_4500_out0;
wire v$JMP_4501_out0;
wire v$LASTQ_12664_out0;
wire v$LASTQ_12665_out0;
wire v$LASTQ_12666_out0;
wire v$LASTQ_12667_out0;
wire v$LASTQ_12668_out0;
wire v$LASTQ_12669_out0;
wire v$LASTQ_12670_out0;
wire v$LASTQ_12671_out0;
wire v$LASTQ_12672_out0;
wire v$LASTQ_12673_out0;
wire v$LASTQ_12674_out0;
wire v$LASTQ_12675_out0;
wire v$LASTQ_12676_out0;
wire v$LASTQ_12677_out0;
wire v$LASTQ_12678_out0;
wire v$LASTQ_12679_out0;
wire v$LASTQ_12680_out0;
wire v$LASTQ_12681_out0;
wire v$LASTQ_12682_out0;
wire v$LASTQ_12683_out0;
wire v$LASTQ_12684_out0;
wire v$LASTQ_12685_out0;
wire v$LDMAINPC_14212_out0;
wire v$LDMAINPC_14213_out0;
wire v$LDMAIN_14395_out0;
wire v$LDMAIN_14396_out0;
wire v$LDMAIN_3427_out0;
wire v$LDMAIN_3428_out0;
wire v$LDSTRAMMUX_16752_out0;
wire v$LDSTRAMMUX_16753_out0;
wire v$LEFT$SHIFT_13403_out0;
wire v$LEFT$SHIFT_13404_out0;
wire v$LEFT$SHIFT_13405_out0;
wire v$LEFT$SHIFT_13406_out0;
wire v$LEFT$SHIFT_13407_out0;
wire v$LEFT$SHIFT_13408_out0;
wire v$LEFT$SHIFT_13409_out0;
wire v$LEFT$SHIFT_13410_out0;
wire v$LEFT$SHIFT_9143_out0;
wire v$LEFT$SHIFT_9144_out0;
wire v$LEFT$SHIFT_9145_out0;
wire v$LEFT$SHIFT_9146_out0;
wire v$LEFT$SHIFT_9147_out0;
wire v$LEFT$SHIFT_9148_out0;
wire v$LEFT$SHIFT_9149_out0;
wire v$LEFT$SHIFT_9150_out0;
wire v$LEFT$SHIT_3255_out0;
wire v$LEFT$SHIT_3256_out0;
wire v$LEFT$SHIT_3257_out0;
wire v$LEFT$SHIT_3258_out0;
wire v$LEFT$SHIT_3259_out0;
wire v$LEFT$SHIT_3260_out0;
wire v$LEFT$SHIT_3261_out0;
wire v$LEFT$SHIT_3262_out0;
wire v$LEFT$SHIT_3263_out0;
wire v$LEFT$SHIT_3264_out0;
wire v$LEFT$SHIT_3265_out0;
wire v$LEFT$SHIT_3266_out0;
wire v$LEFT$SHIT_3267_out0;
wire v$LEFT$SHIT_3268_out0;
wire v$LEFT$SHIT_3269_out0;
wire v$LEFT$SHIT_3270_out0;
wire v$LEFT$SHIT_3271_out0;
wire v$LEFT$SHIT_3272_out0;
wire v$LEFT$SHIT_3273_out0;
wire v$LEFT$SHIT_3274_out0;
wire v$LEFT$SHIT_3275_out0;
wire v$LEFT$SHIT_3276_out0;
wire v$LEFT$SHIT_3277_out0;
wire v$LEFT$SHIT_3278_out0;
wire v$LEFT$SHIT_3279_out0;
wire v$LEFT$SHIT_3280_out0;
wire v$LEFT$SHIT_3281_out0;
wire v$LEFT$SHIT_3282_out0;
wire v$LEFT$SHIT_3283_out0;
wire v$LEFT$SHIT_3284_out0;
wire v$LEFT$SHIT_3285_out0;
wire v$LEFT$SHIT_3286_out0;
wire v$LEFT$SHIT_3287_out0;
wire v$LEFT$SHIT_3288_out0;
wire v$LEFT$SHIT_3289_out0;
wire v$LEFT$SHIT_3290_out0;
wire v$LEFT$SHIT_3291_out0;
wire v$LEFT$SHIT_3292_out0;
wire v$LEFT$SHIT_3293_out0;
wire v$LEFT$SHIT_3294_out0;
wire v$LEFT$SHIT_3295_out0;
wire v$LEFT$SHIT_3296_out0;
wire v$LEFT$SHIT_3297_out0;
wire v$LEFT$SHIT_3298_out0;
wire v$LEFT$SHIT_3299_out0;
wire v$LEFT$SHIT_3300_out0;
wire v$LEFT$SHIT_3301_out0;
wire v$LEFT$SHIT_3302_out0;
wire v$LEFT$SHIT_3303_out0;
wire v$LEFT$SHIT_3304_out0;
wire v$LEFT$SHIT_3305_out0;
wire v$LEFT$SHIT_3306_out0;
wire v$LEFT$SHIT_3307_out0;
wire v$LEFT$SHIT_3308_out0;
wire v$LEFT$SHIT_3309_out0;
wire v$LEFT$SHIT_3310_out0;
wire v$LEFT$SHIT_3311_out0;
wire v$LEFT$SHIT_3312_out0;
wire v$LEFT$SHIT_3313_out0;
wire v$LEFT$SHIT_3314_out0;
wire v$LEFT$SHIT_3315_out0;
wire v$LEFT$SHIT_3316_out0;
wire v$LOADA_5295_out0;
wire v$LOADA_5296_out0;
wire v$LOADA_5363_out0;
wire v$LOADA_5364_out0;
wire v$LOAD_12270_out0;
wire v$LOAD_12271_out0;
wire v$LOAD_6451_out0;
wire v$LOAD_6452_out0;
wire v$LOWER$OUT_4380_out0;
wire v$LOWER$OUT_4381_out0;
wire v$LOWER$OUT_4382_out0;
wire v$LOWER$OUT_4383_out0;
wire v$LOWER$OUT_4384_out0;
wire v$LOWER$OUT_4385_out0;
wire v$LOWER$OUT_4386_out0;
wire v$LOWER$OUT_4387_out0;
wire v$LOWER$OUT_6665_out0;
wire v$LOWER$OUT_6666_out0;
wire v$LOWER$OUT_6667_out0;
wire v$LOWER$OUT_6668_out0;
wire v$LOWER$PART_6568_out0;
wire v$LOWER$PART_6569_out0;
wire v$LOWER$PART_6570_out0;
wire v$LOWER$PART_6571_out0;
wire v$LOWER$SAME_10633_out0;
wire v$LOWER$SAME_10634_out0;
wire v$LOWER$SAME_10635_out0;
wire v$LOWER$SAME_10636_out0;
wire v$LOWER$SAME_10637_out0;
wire v$LOWER$SAME_10638_out0;
wire v$LOWER$SAME_10639_out0;
wire v$LOWER$SAME_10640_out0;
wire v$LOWER$SAME_3975_out0;
wire v$LOWER$SAME_3976_out0;
wire v$LOWER$SAME_3977_out0;
wire v$LOWER$SAME_3978_out0;
wire v$LSB_8138_out0;
wire v$LSB_8139_out0;
wire v$MANTISA$SAME_2630_out0;
wire v$MANTISA$SAME_2631_out0;
wire v$MEMHALT_18405_out0;
wire v$MEMHALT_18406_out0;
wire v$MI$LDST_17607_out0;
wire v$MI$LDST_17608_out0;
wire v$MI_12451_out0;
wire v$MI_12452_out0;
wire v$MI_12694_out0;
wire v$MI_12695_out0;
wire v$MI_13060_out0;
wire v$MI_13061_out0;
wire v$MI_14969_out0;
wire v$MI_14970_out0;
wire v$MI_2609_out0;
wire v$MI_2610_out0;
wire v$MI_6504_out0;
wire v$MI_6505_out0;
wire v$MI_8756_out0;
wire v$MI_8757_out0;
wire v$MODEEN_15721_out0;
wire v$MODEEN_15722_out0;
wire v$MODEEN_6041_out0;
wire v$MODEEN_6042_out0;
wire v$MODEWRITE_15321_out0;
wire v$MODEWRITE_15322_out0;
wire v$MUL_17628_out0;
wire v$MUL_17629_out0;
wire v$MUX10_16266_out0;
wire v$MUX10_16267_out0;
wire v$MUX10_16268_out0;
wire v$MUX10_16269_out0;
wire v$MUX10_17016_out0;
wire v$MUX10_17017_out0;
wire v$MUX11_1353_out0;
wire v$MUX11_1354_out0;
wire v$MUX11_18547_out0;
wire v$MUX11_18548_out0;
wire v$MUX11_18549_out0;
wire v$MUX11_18550_out0;
wire v$MUX12_18419_out0;
wire v$MUX12_18420_out0;
wire v$MUX12_18421_out0;
wire v$MUX12_18422_out0;
wire v$MUX13_14263_out0;
wire v$MUX13_14264_out0;
wire v$MUX13_14265_out0;
wire v$MUX13_14266_out0;
wire v$MUX14_3166_out0;
wire v$MUX14_3167_out0;
wire v$MUX14_5134_out0;
wire v$MUX14_5135_out0;
wire v$MUX14_5136_out0;
wire v$MUX14_5137_out0;
wire v$MUX15_1479_out0;
wire v$MUX15_1480_out0;
wire v$MUX15_1481_out0;
wire v$MUX15_1482_out0;
wire v$MUX15_16530_out0;
wire v$MUX15_16531_out0;
wire v$MUX15_9777_out0;
wire v$MUX15_9778_out0;
wire v$MUX16_17383_out0;
wire v$MUX16_17384_out0;
wire v$MUX16_17385_out0;
wire v$MUX16_17386_out0;
wire v$MUX17_17156_out0;
wire v$MUX17_17157_out0;
wire v$MUX17_17158_out0;
wire v$MUX17_17159_out0;
wire v$MUX17_6767_out0;
wire v$MUX17_6768_out0;
wire v$MUX18_5072_out0;
wire v$MUX18_5073_out0;
wire v$MUX18_5074_out0;
wire v$MUX18_5075_out0;
wire v$MUX19_6614_out0;
wire v$MUX19_6615_out0;
wire v$MUX19_6616_out0;
wire v$MUX19_6617_out0;
wire v$MUX1_2776_out0;
wire v$MUX1_2777_out0;
wire v$MUX1_2778_out0;
wire v$MUX1_2779_out0;
wire v$MUX1_2780_out0;
wire v$MUX1_2781_out0;
wire v$MUX1_2782_out0;
wire v$MUX1_2783_out0;
wire v$MUX1_2784_out0;
wire v$MUX1_2785_out0;
wire v$MUX1_2786_out0;
wire v$MUX1_2787_out0;
wire v$MUX1_3078_out0;
wire v$MUX1_3079_out0;
wire v$MUX1_3080_out0;
wire v$MUX1_3081_out0;
wire v$MUX1_435_out0;
wire v$MUX1_436_out0;
wire v$MUX1_5229_out0;
wire v$MUX1_5230_out0;
wire v$MUX1_7971_out0;
wire v$MUX1_7972_out0;
wire v$MUX20_11892_out0;
wire v$MUX20_11893_out0;
wire v$MUX20_11894_out0;
wire v$MUX20_11895_out0;
wire v$MUX21_5118_out0;
wire v$MUX21_5119_out0;
wire v$MUX21_5120_out0;
wire v$MUX21_5121_out0;
wire v$MUX22_17090_out0;
wire v$MUX22_17091_out0;
wire v$MUX22_17092_out0;
wire v$MUX22_17093_out0;
wire v$MUX23_16833_out0;
wire v$MUX23_16834_out0;
wire v$MUX23_16835_out0;
wire v$MUX23_16836_out0;
wire v$MUX24_18661_out0;
wire v$MUX24_18662_out0;
wire v$MUX24_18663_out0;
wire v$MUX24_18664_out0;
wire v$MUX25_8708_out0;
wire v$MUX25_8709_out0;
wire v$MUX25_8710_out0;
wire v$MUX25_8711_out0;
wire v$MUX2_12801_out0;
wire v$MUX2_12802_out0;
wire v$MUX2_13871_out0;
wire v$MUX2_13872_out0;
wire v$MUX2_14185_out0;
wire v$MUX2_14186_out0;
wire v$MUX2_14187_out0;
wire v$MUX2_14188_out0;
wire v$MUX2_14407_out0;
wire v$MUX2_14408_out0;
wire v$MUX2_14409_out0;
wire v$MUX2_14410_out0;
wire v$MUX2_14411_out0;
wire v$MUX2_14412_out0;
wire v$MUX2_14413_out0;
wire v$MUX2_14414_out0;
wire v$MUX2_14415_out0;
wire v$MUX2_14416_out0;
wire v$MUX2_14417_out0;
wire v$MUX2_14418_out0;
wire v$MUX2_5066_out0;
wire v$MUX2_5067_out0;
wire v$MUX2_6922_out0;
wire v$MUX2_6923_out0;
wire v$MUX3_10374_out0;
wire v$MUX3_10375_out0;
wire v$MUX3_10376_out0;
wire v$MUX3_10377_out0;
wire v$MUX3_10378_out0;
wire v$MUX3_10379_out0;
wire v$MUX3_10380_out0;
wire v$MUX3_10381_out0;
wire v$MUX3_10382_out0;
wire v$MUX3_10383_out0;
wire v$MUX3_10384_out0;
wire v$MUX3_10385_out0;
wire v$MUX3_1579_out0;
wire v$MUX3_1580_out0;
wire v$MUX3_18332_out0;
wire v$MUX3_18333_out0;
wire v$MUX3_6396_out0;
wire v$MUX3_6397_out0;
wire v$MUX3_7928_out0;
wire v$MUX3_7929_out0;
wire v$MUX3_7930_out0;
wire v$MUX3_7931_out0;
wire v$MUX4_12210_out0;
wire v$MUX4_12211_out0;
wire v$MUX4_13221_out0;
wire v$MUX4_13222_out0;
wire v$MUX4_16228_out0;
wire v$MUX4_16229_out0;
wire v$MUX4_17458_out0;
wire v$MUX4_17459_out0;
wire v$MUX4_17460_out0;
wire v$MUX4_17461_out0;
wire v$MUX4_17462_out0;
wire v$MUX4_17463_out0;
wire v$MUX4_17464_out0;
wire v$MUX4_17465_out0;
wire v$MUX4_17466_out0;
wire v$MUX4_17467_out0;
wire v$MUX4_17468_out0;
wire v$MUX4_17469_out0;
wire v$MUX4_17682_out0;
wire v$MUX4_17683_out0;
wire v$MUX4_8124_out0;
wire v$MUX4_8125_out0;
wire v$MUX4_8126_out0;
wire v$MUX4_8127_out0;
wire v$MUX5_12419_out0;
wire v$MUX5_12420_out0;
wire v$MUX5_16091_out0;
wire v$MUX5_16092_out0;
wire v$MUX5_17662_out0;
wire v$MUX5_17663_out0;
wire v$MUX5_19171_out0;
wire v$MUX5_19172_out0;
wire v$MUX5_7209_out0;
wire v$MUX5_7210_out0;
wire v$MUX5_7211_out0;
wire v$MUX5_7212_out0;
wire v$MUX5_9902_out0;
wire v$MUX5_9903_out0;
wire v$MUX5_9904_out0;
wire v$MUX5_9905_out0;
wire v$MUX5_9906_out0;
wire v$MUX5_9907_out0;
wire v$MUX5_9908_out0;
wire v$MUX5_9909_out0;
wire v$MUX5_9910_out0;
wire v$MUX5_9911_out0;
wire v$MUX5_9912_out0;
wire v$MUX5_9913_out0;
wire v$MUX6_10839_out0;
wire v$MUX6_10840_out0;
wire v$MUX6_10841_out0;
wire v$MUX6_10842_out0;
wire v$MUX6_10843_out0;
wire v$MUX6_10844_out0;
wire v$MUX6_10845_out0;
wire v$MUX6_10846_out0;
wire v$MUX6_10847_out0;
wire v$MUX6_10848_out0;
wire v$MUX6_10849_out0;
wire v$MUX6_10850_out0;
wire v$MUX6_14134_out0;
wire v$MUX6_14135_out0;
wire v$MUX6_14320_out0;
wire v$MUX6_14321_out0;
wire v$MUX6_16898_out0;
wire v$MUX6_16899_out0;
wire v$MUX6_16900_out0;
wire v$MUX6_16901_out0;
wire v$MUX6_9458_out0;
wire v$MUX6_9459_out0;
wire v$MUX7_11471_out0;
wire v$MUX7_11472_out0;
wire v$MUX7_1378_out0;
wire v$MUX7_1379_out0;
wire v$MUX7_1380_out0;
wire v$MUX7_1381_out0;
wire v$MUX7_18517_out0;
wire v$MUX7_18518_out0;
wire v$MUX7_18519_out0;
wire v$MUX7_18520_out0;
wire v$MUX7_18521_out0;
wire v$MUX7_18522_out0;
wire v$MUX7_18523_out0;
wire v$MUX7_18524_out0;
wire v$MUX7_18525_out0;
wire v$MUX7_18526_out0;
wire v$MUX7_18527_out0;
wire v$MUX7_18528_out0;
wire v$MUX7_9855_out0;
wire v$MUX7_9856_out0;
wire v$MUX8$OUT_14009_out0;
wire v$MUX8$OUT_14010_out0;
wire v$MUX8_1651_out0;
wire v$MUX8_1652_out0;
wire v$MUX8_3154_out0;
wire v$MUX8_3155_out0;
wire v$MUX8_3156_out0;
wire v$MUX8_3157_out0;
wire v$MUX8_3792_out0;
wire v$MUX8_3793_out0;
wire v$MUX8_3794_out0;
wire v$MUX8_3795_out0;
wire v$MUX8_3796_out0;
wire v$MUX8_3797_out0;
wire v$MUX8_3798_out0;
wire v$MUX8_3799_out0;
wire v$MUX8_3800_out0;
wire v$MUX8_3801_out0;
wire v$MUX8_3802_out0;
wire v$MUX8_3803_out0;
wire v$MUX8_4514_out0;
wire v$MUX8_4515_out0;
wire v$MUX9_8553_out0;
wire v$MUX9_8554_out0;
wire v$MUX9_8555_out0;
wire v$MUX9_8556_out0;
wire v$ModeRegAdd_4164_out0;
wire v$ModeRegAdd_4165_out0;
wire v$ModeWrite_4621_out0;
wire v$ModeWrite_4622_out0;
wire v$NEED$SHIFT$OP1_5034_out0;
wire v$NEED$SHIFT$OP1_5035_out0;
wire v$NEWINTERRUPT_4598_out0;
wire v$NEWINTERRUPT_4599_out0;
wire v$NEWINTERRUPT_5672_out0;
wire v$NEWINTERRUPT_5673_out0;
wire v$NEWINTERRUPT_7309_out0;
wire v$NEWINTERRUPT_7310_out0;
wire v$NEWINT_18407_out0;
wire v$NEWINT_18408_out0;
wire v$NEXTINTERRUPT_13321_out0;
wire v$NEXTINTERRUPT_13322_out0;
wire v$NEXTINTERRUPT_17397_out0;
wire v$NEXTINTERRUPT_17398_out0;
wire v$NEXTINTERRUPT_19041_out0;
wire v$NEXTINTERRUPT_19042_out0;
wire v$NEXTINTERRUPT_19157_out0;
wire v$NEXTINTERRUPT_19158_out0;
wire v$NEXTINT_7282_out0;
wire v$NEXTINT_7283_out0;
wire v$NEXTSTATE_14110_out0;
wire v$NEXTSTATE_14111_out0;
wire v$NEXTSTATE_14112_out0;
wire v$NEXTSTATE_14113_out0;
wire v$NEXTSTATE_14114_out0;
wire v$NEXTSTATE_14115_out0;
wire v$NEXTSTATE_14116_out0;
wire v$NE_3637_out0;
wire v$NE_3638_out0;
wire v$NF_15164_out0;
wire v$NF_15165_out0;
wire v$NOT$USED$CARRY_19386_out0;
wire v$NOT$USED$CARRY_19387_out0;
wire v$NOT$USED$CARRY_19388_out0;
wire v$NOT$USED$CARRY_19389_out0;
wire v$NOT$USED1_14983_out0;
wire v$NOT$USED1_14984_out0;
wire v$NOT$USED1_14985_out0;
wire v$NOT$USED1_14986_out0;
wire v$NOT$USED1_14987_out0;
wire v$NOT$USED1_14988_out0;
wire v$NOT$USED1_14989_out0;
wire v$NOT$USED1_14990_out0;
wire v$NOT$USED_16558_out0;
wire v$NOT$USED_16559_out0;
wire v$NOT$USED_16560_out0;
wire v$NOT$USED_16561_out0;
wire v$NOT$USED_3098_out0;
wire v$NOT$USED_3099_out0;
wire v$NOT$USED_5689_out0;
wire v$NOT$USED_5690_out0;
wire v$NP_7574_out0;
wire v$NP_7575_out0;
wire v$NQ0_15970_out0;
wire v$NQ0_15971_out0;
wire v$NQ0_16214_out0;
wire v$NQ0_16215_out0;
wire v$NQ0_8120_out0;
wire v$NQ0_8121_out0;
wire v$NQ1_11550_out0;
wire v$NQ1_11551_out0;
wire v$NQ1_17350_out0;
wire v$NQ1_17351_out0;
wire v$NQ1_263_out0;
wire v$NQ1_264_out0;
wire v$NQ2_17316_out0;
wire v$NQ2_17317_out0;
wire v$NQ2_19175_out0;
wire v$NQ2_19176_out0;
wire v$NQ2_3191_out0;
wire v$NQ2_3192_out0;
wire v$NQ3_1645_out0;
wire v$NQ3_1646_out0;
wire v$NQ3_3209_out0;
wire v$NQ3_3210_out0;
wire v$NR_17276_out0;
wire v$NR_17277_out0;
wire v$NS_18801_out0;
wire v$NS_18802_out0;
wire v$ODDPARITY_16534_out0;
wire v$ODDPARITY_16535_out0;
wire v$OFF_4196_out0;
wire v$OFF_4197_out0;
wire v$OUTPUT_10799_out0;
wire v$OUTPUT_10800_out0;
wire v$OUTPUT_10801_out0;
wire v$OUTPUT_10802_out0;
wire v$OUTPUT_10803_out0;
wire v$OUTPUT_10804_out0;
wire v$OUTPUT_19087_out0;
wire v$OUT_14341_out0;
wire v$OUT_14342_out0;
wire v$OUT_14343_out0;
wire v$OUT_14344_out0;
wire v$OUT_14345_out0;
wire v$OUT_14346_out0;
wire v$OUT_14347_out0;
wire v$OUT_14348_out0;
wire v$OUT_4021_out0;
wire v$OUT_4022_out0;
wire v$OUT_4076_out0;
wire v$OUT_4077_out0;
wire v$OUT_4078_out0;
wire v$OUT_4079_out0;
wire v$OUT_4080_out0;
wire v$OUT_4081_out0;
wire v$OUT_4082_out0;
wire v$OUT_4083_out0;
wire v$OUT_4084_out0;
wire v$OUT_4085_out0;
wire v$OUT_4086_out0;
wire v$OUT_4087_out0;
wire v$OUT_4088_out0;
wire v$OUT_4089_out0;
wire v$OUT_4090_out0;
wire v$OUT_4091_out0;
wire v$OUT_4092_out0;
wire v$OUT_4093_out0;
wire v$OUT_4094_out0;
wire v$OUT_4095_out0;
wire v$OUT_4096_out0;
wire v$OUT_4097_out0;
wire v$OUT_4098_out0;
wire v$OUT_4099_out0;
wire v$OUT_4100_out0;
wire v$OUT_4101_out0;
wire v$OUT_4102_out0;
wire v$OUT_4103_out0;
wire v$OUT_4104_out0;
wire v$OUT_4105_out0;
wire v$OUT_4106_out0;
wire v$OUT_4107_out0;
wire v$OUT_9267_out0;
wire v$OUT_9268_out0;
wire v$OUT_9269_out0;
wire v$OUT_9270_out0;
wire v$OUT_9851_out0;
wire v$OUT_9852_out0;
wire v$OUT_9853_out0;
wire v$OUT_9854_out0;
wire v$OVERFLOW_15590_out0;
wire v$OVERFLOW_15591_out0;
wire v$OVERFLOW_19065_out0;
wire v$OVERFLOW_19066_out0;
wire v$OVERFLOW_19137_out0;
wire v$OVERFLOW_19138_out0;
wire v$OVERFLOW_3820_out0;
wire v$OVERFLOW_3821_out0;
wire v$OVERFLOW_445_out0;
wire v$OVERFLOW_446_out0;
wire v$OddParity_11182_out0;
wire v$OddParity_11183_out0;
wire v$P$AB_2164_out0;
wire v$P$AB_2165_out0;
wire v$P$AB_2166_out0;
wire v$P$AB_2167_out0;
wire v$P$AB_2168_out0;
wire v$P$AB_2169_out0;
wire v$P$AB_2170_out0;
wire v$P$AB_2171_out0;
wire v$P$AB_2172_out0;
wire v$P$AB_2173_out0;
wire v$P$AB_2174_out0;
wire v$P$AB_2175_out0;
wire v$P$AB_2176_out0;
wire v$P$AB_2177_out0;
wire v$P$AB_2178_out0;
wire v$P$AB_2179_out0;
wire v$P$AB_2180_out0;
wire v$P$AB_2181_out0;
wire v$P$AB_2182_out0;
wire v$P$AB_2183_out0;
wire v$P$AB_2184_out0;
wire v$P$AB_2185_out0;
wire v$P$AB_2186_out0;
wire v$P$AB_2187_out0;
wire v$P$AB_2188_out0;
wire v$P$AB_2189_out0;
wire v$P$AB_2190_out0;
wire v$P$AB_2191_out0;
wire v$P$AB_2192_out0;
wire v$P$AB_2193_out0;
wire v$P$AB_2194_out0;
wire v$P$AB_2195_out0;
wire v$P$AB_2196_out0;
wire v$P$AB_2197_out0;
wire v$P$AB_2198_out0;
wire v$P$AB_2199_out0;
wire v$P$AB_2200_out0;
wire v$P$AB_2201_out0;
wire v$P$AB_2202_out0;
wire v$P$AB_2203_out0;
wire v$P$AB_2204_out0;
wire v$P$AB_2205_out0;
wire v$P$AB_2206_out0;
wire v$P$AB_2207_out0;
wire v$P$AB_2208_out0;
wire v$P$AB_2209_out0;
wire v$P$AB_2210_out0;
wire v$P$AB_2211_out0;
wire v$P$AB_2212_out0;
wire v$P$AB_2213_out0;
wire v$P$AB_2214_out0;
wire v$P$AB_2215_out0;
wire v$P$AB_2216_out0;
wire v$P$AB_2217_out0;
wire v$P$AB_2218_out0;
wire v$P$AB_2219_out0;
wire v$P$AB_2220_out0;
wire v$P$AB_2221_out0;
wire v$P$AB_2222_out0;
wire v$P$AB_2223_out0;
wire v$P$AB_2224_out0;
wire v$P$AB_2225_out0;
wire v$P$AB_2226_out0;
wire v$P$AB_2227_out0;
wire v$P$AB_2228_out0;
wire v$P$AB_2229_out0;
wire v$P$AB_2230_out0;
wire v$P$AB_2231_out0;
wire v$P$AB_2232_out0;
wire v$P$AB_2233_out0;
wire v$P$AB_2234_out0;
wire v$P$AB_2235_out0;
wire v$P$AB_2236_out0;
wire v$P$AB_2237_out0;
wire v$P$AB_2238_out0;
wire v$P$AB_2239_out0;
wire v$P$AB_2240_out0;
wire v$P$AB_2241_out0;
wire v$P$AB_2242_out0;
wire v$P$AB_2243_out0;
wire v$P$AB_2244_out0;
wire v$P$AB_2245_out0;
wire v$P$AB_2246_out0;
wire v$P$AB_2247_out0;
wire v$P$AB_2248_out0;
wire v$P$AB_2249_out0;
wire v$P$AB_2250_out0;
wire v$P$AB_2251_out0;
wire v$P$AB_2252_out0;
wire v$P$AB_2253_out0;
wire v$P$AB_2254_out0;
wire v$P$AB_2255_out0;
wire v$P$AB_2256_out0;
wire v$P$AB_2257_out0;
wire v$P$AB_2258_out0;
wire v$P$AB_2259_out0;
wire v$P$AB_2260_out0;
wire v$P$AB_2261_out0;
wire v$P$AB_2262_out0;
wire v$P$AB_2263_out0;
wire v$P$AB_2264_out0;
wire v$P$AB_2265_out0;
wire v$P$AB_2266_out0;
wire v$P$AB_2267_out0;
wire v$P$AB_2268_out0;
wire v$P$AB_2269_out0;
wire v$P$AB_2270_out0;
wire v$P$AB_2271_out0;
wire v$P$AB_2272_out0;
wire v$P$AB_2273_out0;
wire v$P$AB_2274_out0;
wire v$P$AB_2275_out0;
wire v$P$AB_2276_out0;
wire v$P$AB_2277_out0;
wire v$P$AB_2278_out0;
wire v$P$AB_2279_out0;
wire v$P$AB_2280_out0;
wire v$P$AB_2281_out0;
wire v$P$AB_2282_out0;
wire v$P$AB_2283_out0;
wire v$P$AB_2284_out0;
wire v$P$AB_2285_out0;
wire v$P$AB_2286_out0;
wire v$P$AB_2287_out0;
wire v$P$AB_2288_out0;
wire v$P$AB_2289_out0;
wire v$P$AB_2290_out0;
wire v$P$AB_2291_out0;
wire v$P$AB_2292_out0;
wire v$P$AB_2293_out0;
wire v$P$AB_2294_out0;
wire v$P$AB_2295_out0;
wire v$P$AB_2296_out0;
wire v$P$AB_2297_out0;
wire v$P$AB_2298_out0;
wire v$P$AB_2299_out0;
wire v$P$AB_2300_out0;
wire v$P$AB_2301_out0;
wire v$P$AB_2302_out0;
wire v$P$AB_2303_out0;
wire v$P$AB_2304_out0;
wire v$P$AB_2305_out0;
wire v$P$AB_2306_out0;
wire v$P$AB_2307_out0;
wire v$P$AB_2308_out0;
wire v$P$AB_2309_out0;
wire v$P$AB_2310_out0;
wire v$P$AB_2311_out0;
wire v$P$AB_2312_out0;
wire v$P$AB_2313_out0;
wire v$P$AB_2314_out0;
wire v$P$AB_2315_out0;
wire v$P$AB_2316_out0;
wire v$P$AB_2317_out0;
wire v$P$AB_2318_out0;
wire v$P$AB_2319_out0;
wire v$P$AB_2320_out0;
wire v$P$AB_2321_out0;
wire v$P$AB_2322_out0;
wire v$P$AB_2323_out0;
wire v$P$AB_2324_out0;
wire v$P$AB_2325_out0;
wire v$P$AB_2326_out0;
wire v$P$AB_2327_out0;
wire v$P$AB_2328_out0;
wire v$P$AB_2329_out0;
wire v$P$AB_2330_out0;
wire v$P$AB_2331_out0;
wire v$P$AB_2332_out0;
wire v$P$AB_2333_out0;
wire v$P$AB_2334_out0;
wire v$P$AB_2335_out0;
wire v$P$AB_2336_out0;
wire v$P$AB_2337_out0;
wire v$P$AB_2338_out0;
wire v$P$AB_2339_out0;
wire v$P$AB_2340_out0;
wire v$P$AB_2341_out0;
wire v$P$AB_2342_out0;
wire v$P$AB_2343_out0;
wire v$P$AB_2344_out0;
wire v$P$AB_2345_out0;
wire v$P$AB_2346_out0;
wire v$P$AB_2347_out0;
wire v$P$AB_2348_out0;
wire v$P$AB_2349_out0;
wire v$P$AB_2350_out0;
wire v$P$AB_2351_out0;
wire v$P$AB_2352_out0;
wire v$P$AB_2353_out0;
wire v$P$AB_2354_out0;
wire v$P$AB_2355_out0;
wire v$P$AB_2356_out0;
wire v$P$AB_2357_out0;
wire v$P$AB_2358_out0;
wire v$P$AB_2359_out0;
wire v$P$AB_2360_out0;
wire v$P$AB_2361_out0;
wire v$P$AB_2362_out0;
wire v$P$AB_2363_out0;
wire v$P$AB_2364_out0;
wire v$P$AB_2365_out0;
wire v$P$AB_2366_out0;
wire v$P$AB_2367_out0;
wire v$P$AB_2368_out0;
wire v$P$AB_2369_out0;
wire v$P$AB_2370_out0;
wire v$P$AB_2371_out0;
wire v$P$AB_2372_out0;
wire v$P$AB_2373_out0;
wire v$P$AB_2374_out0;
wire v$P$AB_2375_out0;
wire v$P$AB_2376_out0;
wire v$P$AB_2377_out0;
wire v$P$AB_2378_out0;
wire v$P$AB_2379_out0;
wire v$P$AB_2380_out0;
wire v$P$AB_2381_out0;
wire v$P$AB_2382_out0;
wire v$P$AB_2383_out0;
wire v$P$AB_2384_out0;
wire v$P$AB_2385_out0;
wire v$P$AB_2386_out0;
wire v$P$AB_2387_out0;
wire v$P$AB_2388_out0;
wire v$P$AB_2389_out0;
wire v$P$AB_2390_out0;
wire v$P$AB_2391_out0;
wire v$P$AB_2392_out0;
wire v$P$AB_2393_out0;
wire v$P$AB_2394_out0;
wire v$P$AB_2395_out0;
wire v$P$AB_2396_out0;
wire v$P$AB_2397_out0;
wire v$P$AB_2398_out0;
wire v$P$AB_2399_out0;
wire v$P$AB_2400_out0;
wire v$P$AB_2401_out0;
wire v$P$AB_2402_out0;
wire v$P$AB_2403_out0;
wire v$P$AB_2404_out0;
wire v$P$AB_2405_out0;
wire v$P$AB_2406_out0;
wire v$P$AB_2407_out0;
wire v$P$AB_2408_out0;
wire v$P$AB_2409_out0;
wire v$P$AD_750_out0;
wire v$P$AD_751_out0;
wire v$P$AD_752_out0;
wire v$P$AD_753_out0;
wire v$P$AD_754_out0;
wire v$P$AD_755_out0;
wire v$P$AD_756_out0;
wire v$P$AD_757_out0;
wire v$P$AD_758_out0;
wire v$P$AD_759_out0;
wire v$P$AD_760_out0;
wire v$P$AD_761_out0;
wire v$P$AD_762_out0;
wire v$P$AD_763_out0;
wire v$P$AD_764_out0;
wire v$P$AD_765_out0;
wire v$P$AD_766_out0;
wire v$P$AD_767_out0;
wire v$P$AD_768_out0;
wire v$P$AD_769_out0;
wire v$P$AD_770_out0;
wire v$P$AD_771_out0;
wire v$P$AD_772_out0;
wire v$P$AD_773_out0;
wire v$P$AD_774_out0;
wire v$P$AD_775_out0;
wire v$P$AD_776_out0;
wire v$P$AD_777_out0;
wire v$P$AD_778_out0;
wire v$P$AD_779_out0;
wire v$P$AD_780_out0;
wire v$P$AD_781_out0;
wire v$P$AD_782_out0;
wire v$P$AD_783_out0;
wire v$P$AD_784_out0;
wire v$P$AD_785_out0;
wire v$P$AD_786_out0;
wire v$P$AD_787_out0;
wire v$P$AD_788_out0;
wire v$P$AD_789_out0;
wire v$P$AD_790_out0;
wire v$P$AD_791_out0;
wire v$P$AD_792_out0;
wire v$P$AD_793_out0;
wire v$P$AD_794_out0;
wire v$P$AD_795_out0;
wire v$P$AD_796_out0;
wire v$P$AD_797_out0;
wire v$P$AD_798_out0;
wire v$P$AD_799_out0;
wire v$P$AD_800_out0;
wire v$P$AD_801_out0;
wire v$P$AD_802_out0;
wire v$P$AD_803_out0;
wire v$P$AD_804_out0;
wire v$P$AD_805_out0;
wire v$P$AD_806_out0;
wire v$P$AD_807_out0;
wire v$P$AD_808_out0;
wire v$P$AD_809_out0;
wire v$P$AD_810_out0;
wire v$P$AD_811_out0;
wire v$P$AD_812_out0;
wire v$P$AD_813_out0;
wire v$P$AD_814_out0;
wire v$P$AD_815_out0;
wire v$P$AD_816_out0;
wire v$P$AD_817_out0;
wire v$P$AD_818_out0;
wire v$P$AD_819_out0;
wire v$P$AD_820_out0;
wire v$P$AD_821_out0;
wire v$P$AD_822_out0;
wire v$P$AD_823_out0;
wire v$P$AD_824_out0;
wire v$P$AD_825_out0;
wire v$P$AD_826_out0;
wire v$P$AD_827_out0;
wire v$P$AD_828_out0;
wire v$P$AD_829_out0;
wire v$P$AD_830_out0;
wire v$P$AD_831_out0;
wire v$P$AD_832_out0;
wire v$P$AD_833_out0;
wire v$P$AD_834_out0;
wire v$P$AD_835_out0;
wire v$P$AD_836_out0;
wire v$P$AD_837_out0;
wire v$P$AD_838_out0;
wire v$P$AD_839_out0;
wire v$P$AD_840_out0;
wire v$P$AD_841_out0;
wire v$P$AD_842_out0;
wire v$P$AD_843_out0;
wire v$P$AD_844_out0;
wire v$P$AD_845_out0;
wire v$P$AD_846_out0;
wire v$P$AD_847_out0;
wire v$P$AD_848_out0;
wire v$P$AD_849_out0;
wire v$P$AD_850_out0;
wire v$P$AD_851_out0;
wire v$P$AD_852_out0;
wire v$P$AD_853_out0;
wire v$P$AD_854_out0;
wire v$P$AD_855_out0;
wire v$P$AD_856_out0;
wire v$P$AD_857_out0;
wire v$P$AD_858_out0;
wire v$P$AD_859_out0;
wire v$P$AD_860_out0;
wire v$P$AD_861_out0;
wire v$P$AD_862_out0;
wire v$P$AD_863_out0;
wire v$P$AD_864_out0;
wire v$P$AD_865_out0;
wire v$P$AD_866_out0;
wire v$P$AD_867_out0;
wire v$P$AD_868_out0;
wire v$P$AD_869_out0;
wire v$P$AD_870_out0;
wire v$P$AD_871_out0;
wire v$P$AD_872_out0;
wire v$P$AD_873_out0;
wire v$P$AD_874_out0;
wire v$P$AD_875_out0;
wire v$P$AD_876_out0;
wire v$P$AD_877_out0;
wire v$P$AD_878_out0;
wire v$P$AD_879_out0;
wire v$P$AD_880_out0;
wire v$P$AD_881_out0;
wire v$P$AD_882_out0;
wire v$P$AD_883_out0;
wire v$P$AD_884_out0;
wire v$P$AD_885_out0;
wire v$P$AD_886_out0;
wire v$P$AD_887_out0;
wire v$P$AD_888_out0;
wire v$P$AD_889_out0;
wire v$P$AD_890_out0;
wire v$P$AD_891_out0;
wire v$P$AD_892_out0;
wire v$P$AD_893_out0;
wire v$P$AD_894_out0;
wire v$P$AD_895_out0;
wire v$P$AD_896_out0;
wire v$P$AD_897_out0;
wire v$P$AD_898_out0;
wire v$P$AD_899_out0;
wire v$P$AD_900_out0;
wire v$P$AD_901_out0;
wire v$P$AD_902_out0;
wire v$P$AD_903_out0;
wire v$P$AD_904_out0;
wire v$P$AD_905_out0;
wire v$P$AD_906_out0;
wire v$P$AD_907_out0;
wire v$P$AD_908_out0;
wire v$P$AD_909_out0;
wire v$P$AD_910_out0;
wire v$P$AD_911_out0;
wire v$P$AD_912_out0;
wire v$P$AD_913_out0;
wire v$P$AD_914_out0;
wire v$P$AD_915_out0;
wire v$P$AD_916_out0;
wire v$P$AD_917_out0;
wire v$P$AD_918_out0;
wire v$P$AD_919_out0;
wire v$P$AD_920_out0;
wire v$P$AD_921_out0;
wire v$P$AD_922_out0;
wire v$P$AD_923_out0;
wire v$P$AD_924_out0;
wire v$P$AD_925_out0;
wire v$P$AD_926_out0;
wire v$P$AD_927_out0;
wire v$P$AD_928_out0;
wire v$P$AD_929_out0;
wire v$P$AD_930_out0;
wire v$P$AD_931_out0;
wire v$P$AD_932_out0;
wire v$P$AD_933_out0;
wire v$P$AD_934_out0;
wire v$P$AD_935_out0;
wire v$P$AD_936_out0;
wire v$P$AD_937_out0;
wire v$P$AD_938_out0;
wire v$P$AD_939_out0;
wire v$P$AD_940_out0;
wire v$P$AD_941_out0;
wire v$P$AD_942_out0;
wire v$P$AD_943_out0;
wire v$P$AD_944_out0;
wire v$P$AD_945_out0;
wire v$P$AD_946_out0;
wire v$P$AD_947_out0;
wire v$P$AD_948_out0;
wire v$P$AD_949_out0;
wire v$P$AD_950_out0;
wire v$P$AD_951_out0;
wire v$P$AD_952_out0;
wire v$P$AD_953_out0;
wire v$P$AD_954_out0;
wire v$P$AD_955_out0;
wire v$P$AD_956_out0;
wire v$P$AD_957_out0;
wire v$P$AD_958_out0;
wire v$P$AD_959_out0;
wire v$P$AD_960_out0;
wire v$P$AD_961_out0;
wire v$P$AD_962_out0;
wire v$P$AD_963_out0;
wire v$P$AD_964_out0;
wire v$P$AD_965_out0;
wire v$P$AD_966_out0;
wire v$P$AD_967_out0;
wire v$P$AD_968_out0;
wire v$P$AD_969_out0;
wire v$P$AD_970_out0;
wire v$P$AD_971_out0;
wire v$P$AD_972_out0;
wire v$P$AD_973_out0;
wire v$P$AD_974_out0;
wire v$P$AD_975_out0;
wire v$P$AD_976_out0;
wire v$P$AD_977_out0;
wire v$P$AD_978_out0;
wire v$P$AD_979_out0;
wire v$P$AD_980_out0;
wire v$P$AD_981_out0;
wire v$P$AD_982_out0;
wire v$P$AD_983_out0;
wire v$P$AD_984_out0;
wire v$P$AD_985_out0;
wire v$P$AD_986_out0;
wire v$P$AD_987_out0;
wire v$P$AD_988_out0;
wire v$P$AD_989_out0;
wire v$P$AD_990_out0;
wire v$P$AD_991_out0;
wire v$P$AD_992_out0;
wire v$P$AD_993_out0;
wire v$P$AD_994_out0;
wire v$P$AD_995_out0;
wire v$P$CD_10906_out0;
wire v$P$CD_10907_out0;
wire v$P$CD_10908_out0;
wire v$P$CD_10909_out0;
wire v$P$CD_10910_out0;
wire v$P$CD_10911_out0;
wire v$P$CD_10912_out0;
wire v$P$CD_10913_out0;
wire v$P$CD_10914_out0;
wire v$P$CD_10915_out0;
wire v$P$CD_10916_out0;
wire v$P$CD_10917_out0;
wire v$P$CD_10918_out0;
wire v$P$CD_10919_out0;
wire v$P$CD_10920_out0;
wire v$P$CD_10921_out0;
wire v$P$CD_10922_out0;
wire v$P$CD_10923_out0;
wire v$P$CD_10924_out0;
wire v$P$CD_10925_out0;
wire v$P$CD_10926_out0;
wire v$P$CD_10927_out0;
wire v$P$CD_10928_out0;
wire v$P$CD_10929_out0;
wire v$P$CD_10930_out0;
wire v$P$CD_10931_out0;
wire v$P$CD_10932_out0;
wire v$P$CD_10933_out0;
wire v$P$CD_10934_out0;
wire v$P$CD_10935_out0;
wire v$P$CD_10936_out0;
wire v$P$CD_10937_out0;
wire v$P$CD_10938_out0;
wire v$P$CD_10939_out0;
wire v$P$CD_10940_out0;
wire v$P$CD_10941_out0;
wire v$P$CD_10942_out0;
wire v$P$CD_10943_out0;
wire v$P$CD_10944_out0;
wire v$P$CD_10945_out0;
wire v$P$CD_10946_out0;
wire v$P$CD_10947_out0;
wire v$P$CD_10948_out0;
wire v$P$CD_10949_out0;
wire v$P$CD_10950_out0;
wire v$P$CD_10951_out0;
wire v$P$CD_10952_out0;
wire v$P$CD_10953_out0;
wire v$P$CD_10954_out0;
wire v$P$CD_10955_out0;
wire v$P$CD_10956_out0;
wire v$P$CD_10957_out0;
wire v$P$CD_10958_out0;
wire v$P$CD_10959_out0;
wire v$P$CD_10960_out0;
wire v$P$CD_10961_out0;
wire v$P$CD_10962_out0;
wire v$P$CD_10963_out0;
wire v$P$CD_10964_out0;
wire v$P$CD_10965_out0;
wire v$P$CD_10966_out0;
wire v$P$CD_10967_out0;
wire v$P$CD_10968_out0;
wire v$P$CD_10969_out0;
wire v$P$CD_10970_out0;
wire v$P$CD_10971_out0;
wire v$P$CD_10972_out0;
wire v$P$CD_10973_out0;
wire v$P$CD_10974_out0;
wire v$P$CD_10975_out0;
wire v$P$CD_10976_out0;
wire v$P$CD_10977_out0;
wire v$P$CD_10978_out0;
wire v$P$CD_10979_out0;
wire v$P$CD_10980_out0;
wire v$P$CD_10981_out0;
wire v$P$CD_10982_out0;
wire v$P$CD_10983_out0;
wire v$P$CD_10984_out0;
wire v$P$CD_10985_out0;
wire v$P$CD_10986_out0;
wire v$P$CD_10987_out0;
wire v$P$CD_10988_out0;
wire v$P$CD_10989_out0;
wire v$P$CD_10990_out0;
wire v$P$CD_10991_out0;
wire v$P$CD_10992_out0;
wire v$P$CD_10993_out0;
wire v$P$CD_10994_out0;
wire v$P$CD_10995_out0;
wire v$P$CD_10996_out0;
wire v$P$CD_10997_out0;
wire v$P$CD_10998_out0;
wire v$P$CD_10999_out0;
wire v$P$CD_11000_out0;
wire v$P$CD_11001_out0;
wire v$P$CD_11002_out0;
wire v$P$CD_11003_out0;
wire v$P$CD_11004_out0;
wire v$P$CD_11005_out0;
wire v$P$CD_11006_out0;
wire v$P$CD_11007_out0;
wire v$P$CD_11008_out0;
wire v$P$CD_11009_out0;
wire v$P$CD_11010_out0;
wire v$P$CD_11011_out0;
wire v$P$CD_11012_out0;
wire v$P$CD_11013_out0;
wire v$P$CD_11014_out0;
wire v$P$CD_11015_out0;
wire v$P$CD_11016_out0;
wire v$P$CD_11017_out0;
wire v$P$CD_11018_out0;
wire v$P$CD_11019_out0;
wire v$P$CD_11020_out0;
wire v$P$CD_11021_out0;
wire v$P$CD_11022_out0;
wire v$P$CD_11023_out0;
wire v$P$CD_11024_out0;
wire v$P$CD_11025_out0;
wire v$P$CD_11026_out0;
wire v$P$CD_11027_out0;
wire v$P$CD_11028_out0;
wire v$P$CD_11029_out0;
wire v$P$CD_11030_out0;
wire v$P$CD_11031_out0;
wire v$P$CD_11032_out0;
wire v$P$CD_11033_out0;
wire v$P$CD_11034_out0;
wire v$P$CD_11035_out0;
wire v$P$CD_11036_out0;
wire v$P$CD_11037_out0;
wire v$P$CD_11038_out0;
wire v$P$CD_11039_out0;
wire v$P$CD_11040_out0;
wire v$P$CD_11041_out0;
wire v$P$CD_11042_out0;
wire v$P$CD_11043_out0;
wire v$P$CD_11044_out0;
wire v$P$CD_11045_out0;
wire v$P$CD_11046_out0;
wire v$P$CD_11047_out0;
wire v$P$CD_11048_out0;
wire v$P$CD_11049_out0;
wire v$P$CD_11050_out0;
wire v$P$CD_11051_out0;
wire v$P$CD_11052_out0;
wire v$P$CD_11053_out0;
wire v$P$CD_11054_out0;
wire v$P$CD_11055_out0;
wire v$P$CD_11056_out0;
wire v$P$CD_11057_out0;
wire v$P$CD_11058_out0;
wire v$P$CD_11059_out0;
wire v$P$CD_11060_out0;
wire v$P$CD_11061_out0;
wire v$P$CD_11062_out0;
wire v$P$CD_11063_out0;
wire v$P$CD_11064_out0;
wire v$P$CD_11065_out0;
wire v$P$CD_11066_out0;
wire v$P$CD_11067_out0;
wire v$P$CD_11068_out0;
wire v$P$CD_11069_out0;
wire v$P$CD_11070_out0;
wire v$P$CD_11071_out0;
wire v$P$CD_11072_out0;
wire v$P$CD_11073_out0;
wire v$P$CD_11074_out0;
wire v$P$CD_11075_out0;
wire v$P$CD_11076_out0;
wire v$P$CD_11077_out0;
wire v$P$CD_11078_out0;
wire v$P$CD_11079_out0;
wire v$P$CD_11080_out0;
wire v$P$CD_11081_out0;
wire v$P$CD_11082_out0;
wire v$P$CD_11083_out0;
wire v$P$CD_11084_out0;
wire v$P$CD_11085_out0;
wire v$P$CD_11086_out0;
wire v$P$CD_11087_out0;
wire v$P$CD_11088_out0;
wire v$P$CD_11089_out0;
wire v$P$CD_11090_out0;
wire v$P$CD_11091_out0;
wire v$P$CD_11092_out0;
wire v$P$CD_11093_out0;
wire v$P$CD_11094_out0;
wire v$P$CD_11095_out0;
wire v$P$CD_11096_out0;
wire v$P$CD_11097_out0;
wire v$P$CD_11098_out0;
wire v$P$CD_11099_out0;
wire v$P$CD_11100_out0;
wire v$P$CD_11101_out0;
wire v$P$CD_11102_out0;
wire v$P$CD_11103_out0;
wire v$P$CD_11104_out0;
wire v$P$CD_11105_out0;
wire v$P$CD_11106_out0;
wire v$P$CD_11107_out0;
wire v$P$CD_11108_out0;
wire v$P$CD_11109_out0;
wire v$P$CD_11110_out0;
wire v$P$CD_11111_out0;
wire v$P$CD_11112_out0;
wire v$P$CD_11113_out0;
wire v$P$CD_11114_out0;
wire v$P$CD_11115_out0;
wire v$P$CD_11116_out0;
wire v$P$CD_11117_out0;
wire v$P$CD_11118_out0;
wire v$P$CD_11119_out0;
wire v$P$CD_11120_out0;
wire v$P$CD_11121_out0;
wire v$P$CD_11122_out0;
wire v$P$CD_11123_out0;
wire v$P$CD_11124_out0;
wire v$P$CD_11125_out0;
wire v$P$CD_11126_out0;
wire v$P$CD_11127_out0;
wire v$P$CD_11128_out0;
wire v$P$CD_11129_out0;
wire v$P$CD_11130_out0;
wire v$P$CD_11131_out0;
wire v$P$CD_11132_out0;
wire v$P$CD_11133_out0;
wire v$P$CD_11134_out0;
wire v$P$CD_11135_out0;
wire v$P$CD_11136_out0;
wire v$P$CD_11137_out0;
wire v$P$CD_11138_out0;
wire v$P$CD_11139_out0;
wire v$P$CD_11140_out0;
wire v$P$CD_11141_out0;
wire v$P$CD_11142_out0;
wire v$P$CD_11143_out0;
wire v$P$CD_11144_out0;
wire v$P$CD_11145_out0;
wire v$P$CD_11146_out0;
wire v$P$CD_11147_out0;
wire v$P$CD_11148_out0;
wire v$P$CD_11149_out0;
wire v$P$CD_11150_out0;
wire v$P$CD_11151_out0;
wire v$P0_5023_out0;
wire v$P0_5024_out0;
wire v$P0_5025_out0;
wire v$P0_5026_out0;
wire v$P0_5027_out0;
wire v$P0_5028_out0;
wire v$P10_360_out0;
wire v$P10_361_out0;
wire v$P10_362_out0;
wire v$P10_363_out0;
wire v$P10_364_out0;
wire v$P10_365_out0;
wire v$P11_9992_out0;
wire v$P11_9993_out0;
wire v$P11_9994_out0;
wire v$P11_9995_out0;
wire v$P11_9996_out0;
wire v$P11_9997_out0;
wire v$P12_243_out0;
wire v$P12_244_out0;
wire v$P12_245_out0;
wire v$P12_246_out0;
wire v$P12_247_out0;
wire v$P12_248_out0;
wire v$P13_3245_out0;
wire v$P13_3246_out0;
wire v$P13_3247_out0;
wire v$P13_3248_out0;
wire v$P13_3249_out0;
wire v$P13_3250_out0;
wire v$P14_3369_out0;
wire v$P14_3370_out0;
wire v$P14_3371_out0;
wire v$P14_3372_out0;
wire v$P14_3373_out0;
wire v$P14_3374_out0;
wire v$P15_7183_out0;
wire v$P15_7184_out0;
wire v$P15_7185_out0;
wire v$P15_7186_out0;
wire v$P15_7187_out0;
wire v$P15_7188_out0;
wire v$P16_7243_out0;
wire v$P16_7244_out0;
wire v$P16_7245_out0;
wire v$P16_7246_out0;
wire v$P16_7247_out0;
wire v$P16_7248_out0;
wire v$P17_12328_out0;
wire v$P17_12329_out0;
wire v$P17_12330_out0;
wire v$P17_12331_out0;
wire v$P17_12332_out0;
wire v$P17_12333_out0;
wire v$P18_12290_out0;
wire v$P18_12291_out0;
wire v$P18_12292_out0;
wire v$P18_12293_out0;
wire v$P18_12294_out0;
wire v$P18_12295_out0;
wire v$P19_16932_out0;
wire v$P19_16933_out0;
wire v$P19_16934_out0;
wire v$P19_16935_out0;
wire v$P19_16936_out0;
wire v$P19_16937_out0;
wire v$P1_3168_out0;
wire v$P1_3169_out0;
wire v$P1_3170_out0;
wire v$P1_3171_out0;
wire v$P1_3172_out0;
wire v$P1_3173_out0;
wire v$P20_11152_out0;
wire v$P20_11153_out0;
wire v$P20_11154_out0;
wire v$P20_11155_out0;
wire v$P20_11156_out0;
wire v$P20_11157_out0;
wire v$P21_4981_out0;
wire v$P21_4982_out0;
wire v$P21_4983_out0;
wire v$P21_4984_out0;
wire v$P21_4985_out0;
wire v$P21_4986_out0;
wire v$P22_4945_out0;
wire v$P22_4946_out0;
wire v$P22_4947_out0;
wire v$P22_4948_out0;
wire v$P22_4949_out0;
wire v$P22_4950_out0;
wire v$P23_6626_out0;
wire v$P23_6627_out0;
wire v$P23_6628_out0;
wire v$P23_6629_out0;
wire v$P23_6630_out0;
wire v$P23_6631_out0;
wire v$P2_2424_out0;
wire v$P2_2425_out0;
wire v$P2_2426_out0;
wire v$P2_2427_out0;
wire v$P2_2428_out0;
wire v$P2_2429_out0;
wire v$P3_15921_out0;
wire v$P3_15922_out0;
wire v$P3_15923_out0;
wire v$P3_15924_out0;
wire v$P3_15925_out0;
wire v$P3_15926_out0;
wire v$P4_14214_out0;
wire v$P4_14215_out0;
wire v$P4_14216_out0;
wire v$P4_14217_out0;
wire v$P4_14218_out0;
wire v$P4_14219_out0;
wire v$P5_228_out0;
wire v$P5_229_out0;
wire v$P5_230_out0;
wire v$P5_231_out0;
wire v$P5_232_out0;
wire v$P5_233_out0;
wire v$P6_8418_out0;
wire v$P6_8419_out0;
wire v$P6_8420_out0;
wire v$P6_8421_out0;
wire v$P6_8422_out0;
wire v$P6_8423_out0;
wire v$P7_12338_out0;
wire v$P7_12339_out0;
wire v$P7_12340_out0;
wire v$P7_12341_out0;
wire v$P7_12342_out0;
wire v$P7_12343_out0;
wire v$P8_1861_out0;
wire v$P8_1862_out0;
wire v$P8_1863_out0;
wire v$P8_1864_out0;
wire v$P8_1865_out0;
wire v$P8_1866_out0;
wire v$P9_19053_out0;
wire v$P9_19054_out0;
wire v$P9_19055_out0;
wire v$P9_19056_out0;
wire v$P9_19057_out0;
wire v$P9_19058_out0;
wire v$PARITY_12637_out0;
wire v$PARITY_12638_out0;
wire v$PCHALTVIEWER_1929_out0;
wire v$PCHALT_13316_out0;
wire v$PCHALT_17182_out0;
wire v$PHALT0$PREV_7940_out0;
wire v$PHALT0_12199_out0;
wire v$PHALT1$PREV_7682_out0;
wire v$PHALT1_9264_out0;
wire v$PHALTVIEWER_2846_out0;
wire v$PHALT_15747_out0;
wire v$PHALT_1794_out0;
wire v$PHALT_18124_out0;
wire v$PIPELINE$RESTART_19235_out0;
wire v$PIPELINE$RESTART_19236_out0;
wire v$PIPELINE$RESTART_6348_out0;
wire v$PIPELINE$RESTART_6349_out0;
wire v$PIPELINEHALT_15423_out0;
wire v$PIPELINEHALT_15424_out0;
wire v$PIPELINERESTART_2611_out0;
wire v$PIPELINERESTART_2612_out0;
wire v$P_14453_out0;
wire v$P_14454_out0;
wire v$P_14455_out0;
wire v$P_14456_out0;
wire v$P_14457_out0;
wire v$P_14458_out0;
wire v$P_14459_out0;
wire v$P_14460_out0;
wire v$P_14461_out0;
wire v$P_14462_out0;
wire v$P_14463_out0;
wire v$P_14464_out0;
wire v$P_14465_out0;
wire v$P_14466_out0;
wire v$P_14467_out0;
wire v$P_14468_out0;
wire v$P_14469_out0;
wire v$P_14470_out0;
wire v$P_14471_out0;
wire v$P_14472_out0;
wire v$P_14473_out0;
wire v$P_14474_out0;
wire v$P_14475_out0;
wire v$P_14476_out0;
wire v$P_14477_out0;
wire v$P_14478_out0;
wire v$P_14479_out0;
wire v$P_14480_out0;
wire v$P_14481_out0;
wire v$P_14482_out0;
wire v$P_14483_out0;
wire v$P_14484_out0;
wire v$P_14485_out0;
wire v$P_14486_out0;
wire v$P_14487_out0;
wire v$P_14488_out0;
wire v$P_14489_out0;
wire v$P_14490_out0;
wire v$P_14491_out0;
wire v$P_14492_out0;
wire v$P_14493_out0;
wire v$P_14494_out0;
wire v$P_14495_out0;
wire v$P_14496_out0;
wire v$P_14497_out0;
wire v$P_14498_out0;
wire v$P_14499_out0;
wire v$P_14500_out0;
wire v$P_14501_out0;
wire v$P_14502_out0;
wire v$P_14503_out0;
wire v$P_14504_out0;
wire v$P_14505_out0;
wire v$P_14506_out0;
wire v$P_14507_out0;
wire v$P_14508_out0;
wire v$P_14509_out0;
wire v$P_14510_out0;
wire v$P_14511_out0;
wire v$P_14512_out0;
wire v$P_14513_out0;
wire v$P_14514_out0;
wire v$P_14515_out0;
wire v$P_14516_out0;
wire v$P_14517_out0;
wire v$P_14518_out0;
wire v$P_14519_out0;
wire v$P_14520_out0;
wire v$P_14521_out0;
wire v$P_14522_out0;
wire v$P_14523_out0;
wire v$P_14524_out0;
wire v$P_14525_out0;
wire v$P_14526_out0;
wire v$P_14527_out0;
wire v$P_14528_out0;
wire v$P_14529_out0;
wire v$P_14530_out0;
wire v$P_14531_out0;
wire v$P_14532_out0;
wire v$P_14533_out0;
wire v$P_14534_out0;
wire v$P_14535_out0;
wire v$P_14536_out0;
wire v$P_14537_out0;
wire v$P_14538_out0;
wire v$P_14539_out0;
wire v$P_14540_out0;
wire v$P_14541_out0;
wire v$P_14542_out0;
wire v$P_14543_out0;
wire v$P_14544_out0;
wire v$P_14545_out0;
wire v$P_14546_out0;
wire v$P_14547_out0;
wire v$P_14548_out0;
wire v$P_14549_out0;
wire v$P_14550_out0;
wire v$P_14551_out0;
wire v$P_14552_out0;
wire v$P_14553_out0;
wire v$P_14554_out0;
wire v$P_14555_out0;
wire v$P_14556_out0;
wire v$P_14557_out0;
wire v$P_14558_out0;
wire v$P_14559_out0;
wire v$P_14560_out0;
wire v$P_14561_out0;
wire v$P_14562_out0;
wire v$P_14563_out0;
wire v$P_14564_out0;
wire v$P_14565_out0;
wire v$P_14566_out0;
wire v$P_14567_out0;
wire v$P_14568_out0;
wire v$P_14569_out0;
wire v$P_14570_out0;
wire v$P_14571_out0;
wire v$P_14572_out0;
wire v$P_14573_out0;
wire v$P_14574_out0;
wire v$P_14575_out0;
wire v$P_14576_out0;
wire v$P_14577_out0;
wire v$P_14578_out0;
wire v$P_14579_out0;
wire v$P_14580_out0;
wire v$P_14581_out0;
wire v$P_14582_out0;
wire v$P_14583_out0;
wire v$P_14584_out0;
wire v$P_14585_out0;
wire v$P_14586_out0;
wire v$P_14587_out0;
wire v$P_14588_out0;
wire v$P_14589_out0;
wire v$P_14590_out0;
wire v$P_14591_out0;
wire v$P_14592_out0;
wire v$P_14593_out0;
wire v$P_14594_out0;
wire v$P_14595_out0;
wire v$P_14596_out0;
wire v$P_8621_out0;
wire v$P_8622_out0;
wire v$ParityCheck_16733_out0;
wire v$ParityCheck_16734_out0;
wire v$ParityEN_16385_out0;
wire v$ParityEN_16386_out0;
wire v$Q0P_12736_out0;
wire v$Q0P_12737_out0;
wire v$Q0P_17393_out0;
wire v$Q0P_17394_out0;
wire v$Q0_14284_out0;
wire v$Q0_14285_out0;
wire v$Q0_18924_out0;
wire v$Q0_18925_out0;
wire v$Q0_74_out0;
wire v$Q0_75_out0;
wire v$Q1P_11515_out0;
wire v$Q1P_11516_out0;
wire v$Q1P_6027_out0;
wire v$Q1P_6028_out0;
wire v$Q1_11427_out0;
wire v$Q1_11428_out0;
wire v$Q1_14930_out0;
wire v$Q1_14931_out0;
wire v$Q1_4619_out0;
wire v$Q1_4620_out0;
wire v$Q2P_4318_out0;
wire v$Q2P_4319_out0;
wire v$Q2P_6320_out0;
wire v$Q2P_6321_out0;
wire v$Q2_18125_out0;
wire v$Q2_18126_out0;
wire v$Q2_3367_out0;
wire v$Q2_3368_out0;
wire v$Q2_5696_out0;
wire v$Q2_5697_out0;
wire v$Q3P_12238_out0;
wire v$Q3P_12239_out0;
wire v$Q3P_14397_out0;
wire v$Q3P_14398_out0;
wire v$Q3_18893_out0;
wire v$Q3_18894_out0;
wire v$Q3_19033_out0;
wire v$Q3_19034_out0;
wire v$Q_14753_out0;
wire v$Q_14754_out0;
wire v$Q_14755_out0;
wire v$Q_14756_out0;
wire v$Q_14757_out0;
wire v$Q_14758_out0;
wire v$Q_14759_out0;
wire v$Q_14760_out0;
wire v$Q_14761_out0;
wire v$Q_14762_out0;
wire v$Q_14763_out0;
wire v$Q_14764_out0;
wire v$Q_14765_out0;
wire v$Q_14766_out0;
wire v$Q_14767_out0;
wire v$Q_14768_out0;
wire v$Q_14769_out0;
wire v$Q_14770_out0;
wire v$Q_14771_out0;
wire v$Q_14772_out0;
wire v$Q_14773_out0;
wire v$Q_14774_out0;
wire v$R0_15792_out0;
wire v$R0_15793_out0;
wire v$R0_2163_out0;
wire v$R0_6913_out0;
wire v$R1_12459_out0;
wire v$R1_15628_out0;
wire v$R1_15629_out0;
wire v$R1_18512_out0;
wire v$R2_4026_out0;
wire v$R2_4027_out0;
wire v$R3_15899_out0;
wire v$R3_15900_out0;
wire v$RAMWEN0_17189_out0;
wire v$RAMWEN1_11257_out0;
wire v$RAMWENVIEWER_17930_out0;
wire v$RAMWEN_16256_out0;
wire v$RAMWEN_16257_out0;
wire v$RAMWEN_18576_out0;
wire v$RAMWEN_8084_out0;
wire v$RAMWEN_8085_out0;
wire v$READ$REQUEST0_11924_out0;
wire v$READ$REQUEST0_19088_out0;
wire v$READ$REQUEST1_17439_out0;
wire v$READ$REQUEST1_6717_out0;
wire v$READ$REQUEST_15062_out0;
wire v$READ$REQUEST_15063_out0;
wire v$READ$REQUEST_17172_out0;
wire v$READ$REQUEST_17173_out0;
wire v$READ$REQUEST_8130_out0;
wire v$READ$REQUEST_8131_out0;
wire v$RECIEVEDPARITY_6488_out0;
wire v$RECIEVEDPARITY_6489_out0;
wire v$RR0VIEWER_15261_out0;
wire v$RR0_8403_out0;
wire v$RR1REGoutVIEWER_7695_out0;
wire v$RR1VIEWER_15650_out0;
wire v$RR1_2111_out0;
wire v$RXBIT_9243_out0;
wire v$RXBIT_9244_out0;
wire v$RXCLK_1393_out0;
wire v$RXCLK_1394_out0;
wire v$RXCLK_16448_out0;
wire v$RXCLK_16449_out0;
wire v$RXDISABLE_8214_out0;
wire v$RXDISABLE_8215_out0;
wire v$RXENABLE_3897_out0;
wire v$RXENABLE_3898_out0;
wire v$RXErrorSet_3679_out0;
wire v$RXErrorSet_3680_out0;
wire v$RXFLAG_12700_out0;
wire v$RXFLAG_12701_out0;
wire v$RXFLAG_15620_out0;
wire v$RXFLAG_15621_out0;
wire v$RXFlagSet_9435_out0;
wire v$RXFlagSet_9436_out0;
wire v$RXINTERRUPT_15456_out0;
wire v$RXINTERRUPT_15457_out0;
wire v$RXINTERRUPT_15935_out0;
wire v$RXINTERRUPT_15936_out0;
wire v$RXINT_13139_out0;
wire v$RXINT_13140_out0;
wire v$RXREAD_15931_out0;
wire v$RXREAD_15932_out0;
wire v$RXREAD_16458_out0;
wire v$RXREAD_16459_out0;
wire v$RXRead_16983_out0;
wire v$RXRead_16984_out0;
wire v$RXRegAdd_13546_out0;
wire v$RXRegAdd_13547_out0;
wire v$RXReset_17150_out0;
wire v$RXReset_17151_out0;
wire v$RXSET_15291_out0;
wire v$RXSET_15292_out0;
wire v$RXSHIFT_736_out0;
wire v$RXSHIFT_737_out0;
wire v$RX_3176_out0;
wire v$RX_3177_out0;
wire v$RX_44_out0;
wire v$RX_45_out0;
wire v$RX_5021_out0;
wire v$RX_5022_out0;
wire v$RX_6447_out0;
wire v$RX_6448_out0;
wire v$RX_6887_out0;
wire v$RX_6888_out0;
wire v$RXflag_16445_out0;
wire v$RXflag_16446_out0;
wire v$RXlast_13391_out0;
wire v$RXlast_13392_out0;
wire v$RXoverflow_9918_out0;
wire v$RXoverflow_9919_out0;
wire v$RXreset_6240_out0;
wire v$RXreset_6241_out0;
wire v$RXset_1859_out0;
wire v$RXset_1860_out0;
wire v$RXset_5317_out0;
wire v$RXset_5318_out0;
wire v$R_1639_out0;
wire v$R_1640_out0;
wire v$R_1641_out0;
wire v$R_1642_out0;
wire v$R_1643_out0;
wire v$R_1644_out0;
wire v$R_17367_out0;
wire v$R_1743_out0;
wire v$R_1744_out0;
wire v$R_1745_out0;
wire v$R_1746_out0;
wire v$R_1747_out0;
wire v$R_1748_out0;
wire v$R_1749_out0;
wire v$R_18936_out0;
wire v$R_18937_out0;
wire v$R_18938_out0;
wire v$R_18939_out0;
wire v$R_18940_out0;
wire v$R_18941_out0;
wire v$R_18942_out0;
wire v$R_18943_out0;
wire v$R_18944_out0;
wire v$R_18945_out0;
wire v$R_18946_out0;
wire v$R_18947_out0;
wire v$R_18948_out0;
wire v$R_18949_out0;
wire v$R_18950_out0;
wire v$R_18951_out0;
wire v$R_18952_out0;
wire v$R_18953_out0;
wire v$R_18954_out0;
wire v$R_18955_out0;
wire v$R_18956_out0;
wire v$R_18957_out0;
wire v$R_9127_out0;
wire v$R_9128_out0;
wire v$RceivedParity_19151_out0;
wire v$RceivedParity_19152_out0;
wire v$RecievedParity_9916_out0;
wire v$RecievedParity_9917_out0;
wire v$SAME$H_1301_out0;
wire v$SAME$H_1302_out0;
wire v$SAME$H_9245_out0;
wire v$SAME$H_9246_out0;
wire v$SAME$L_17063_out0;
wire v$SAME$L_17064_out0;
wire v$SAME$L_9837_out0;
wire v$SAME$L_9838_out0;
wire v$SAME_18968_out0;
wire v$SAME_18969_out0;
wire v$SAME_18970_out0;
wire v$SAME_18971_out0;
wire v$SAME_18972_out0;
wire v$SAME_18973_out0;
wire v$SAME_18974_out0;
wire v$SAME_18975_out0;
wire v$SAME_19333_out0;
wire v$SAME_19334_out0;
wire v$SAME_19335_out0;
wire v$SAME_19336_out0;
wire v$SAME_19337_out0;
wire v$SAME_19338_out0;
wire v$SAME_19339_out0;
wire v$SAME_19340_out0;
wire v$SAME_19341_out0;
wire v$SAME_19342_out0;
wire v$SAME_19343_out0;
wire v$SAME_19344_out0;
wire v$SAME_19345_out0;
wire v$SAME_19346_out0;
wire v$SAME_19347_out0;
wire v$SAME_19348_out0;
wire v$SAME_19349_out0;
wire v$SAME_19350_out0;
wire v$SAME_19351_out0;
wire v$SAME_19352_out0;
wire v$SAME_19353_out0;
wire v$SAME_19354_out0;
wire v$SAME_19355_out0;
wire v$SAME_19356_out0;
wire v$SAME_19357_out0;
wire v$SAME_19358_out0;
wire v$SAME_19359_out0;
wire v$SAME_19360_out0;
wire v$SAME_19361_out0;
wire v$SAME_19362_out0;
wire v$SAME_19363_out0;
wire v$SAME_19364_out0;
wire v$SAME_6530_out0;
wire v$SAME_6531_out0;
wire v$SAME_9249_out0;
wire v$SAME_9250_out0;
wire v$SAME_9251_out0;
wire v$SAME_9252_out0;
wire v$SEL10_13189_out0;
wire v$SEL10_13190_out0;
wire v$SEL10_13191_out0;
wire v$SEL10_13192_out0;
wire v$SEL10_13193_out0;
wire v$SEL10_13194_out0;
wire v$SEL10_13195_out0;
wire v$SEL10_13196_out0;
wire v$SEL10_13197_out0;
wire v$SEL10_13198_out0;
wire v$SEL10_13199_out0;
wire v$SEL10_13200_out0;
wire v$SEL10_13201_out0;
wire v$SEL10_13202_out0;
wire v$SEL10_13203_out0;
wire v$SEL10_13204_out0;
wire v$SEL10_13205_out0;
wire v$SEL10_13206_out0;
wire v$SEL10_13207_out0;
wire v$SEL10_13208_out0;
wire v$SEL10_13209_out0;
wire v$SEL10_13210_out0;
wire v$SEL10_13211_out0;
wire v$SEL10_13212_out0;
wire v$SEL10_4311_out0;
wire v$SEL10_4312_out0;
wire v$SEL10_7597_out0;
wire v$SEL10_7598_out0;
wire v$SEL10_9883_out0;
wire v$SEL10_9884_out0;
wire v$SEL10_9885_out0;
wire v$SEL10_9886_out0;
wire v$SEL11_12766_out0;
wire v$SEL11_12767_out0;
wire v$SEL11_16147_out0;
wire v$SEL11_16148_out0;
wire v$SEL11_16493_out0;
wire v$SEL11_16494_out0;
wire v$SEL11_7539_out0;
wire v$SEL11_7540_out0;
wire v$SEL11_7541_out0;
wire v$SEL11_7542_out0;
wire v$SEL11_8654_out0;
wire v$SEL11_8655_out0;
wire v$SEL12_14433_out0;
wire v$SEL12_14434_out0;
wire v$SEL12_14435_out0;
wire v$SEL12_14436_out0;
wire v$SEL12_1513_out0;
wire v$SEL12_1514_out0;
wire v$SEL13_13831_out0;
wire v$SEL13_13832_out0;
wire v$SEL13_18204_out0;
wire v$SEL13_18205_out0;
wire v$SEL13_7205_out0;
wire v$SEL13_7206_out0;
wire v$SEL13_7207_out0;
wire v$SEL13_7208_out0;
wire v$SEL14_16964_out0;
wire v$SEL14_16965_out0;
wire v$SEL14_16966_out0;
wire v$SEL14_16967_out0;
wire v$SEL15_14189_out0;
wire v$SEL15_14190_out0;
wire v$SEL15_5102_out0;
wire v$SEL15_5103_out0;
wire v$SEL15_5104_out0;
wire v$SEL15_5105_out0;
wire v$SEL16_17505_out0;
wire v$SEL16_17506_out0;
wire v$SEL16_17507_out0;
wire v$SEL16_17508_out0;
wire v$SEL17_16683_out0;
wire v$SEL17_16684_out0;
wire v$SEL17_16685_out0;
wire v$SEL17_16686_out0;
wire v$SEL18_11908_out0;
wire v$SEL18_11909_out0;
wire v$SEL18_11910_out0;
wire v$SEL18_11911_out0;
wire v$SEL19_13385_out0;
wire v$SEL19_13386_out0;
wire v$SEL19_13387_out0;
wire v$SEL19_13388_out0;
wire v$SEL1_13940_out0;
wire v$SEL1_13941_out0;
wire v$SEL1_13942_out0;
wire v$SEL1_13943_out0;
wire v$SEL1_14044_out0;
wire v$SEL1_14045_out0;
wire v$SEL1_14046_out0;
wire v$SEL1_14047_out0;
wire v$SEL1_14048_out0;
wire v$SEL1_14049_out0;
wire v$SEL1_14050_out0;
wire v$SEL1_14051_out0;
wire v$SEL1_14052_out0;
wire v$SEL1_14053_out0;
wire v$SEL1_14054_out0;
wire v$SEL1_14055_out0;
wire v$SEL1_14056_out0;
wire v$SEL1_14057_out0;
wire v$SEL1_14058_out0;
wire v$SEL1_14059_out0;
wire v$SEL1_14060_out0;
wire v$SEL1_14061_out0;
wire v$SEL1_14062_out0;
wire v$SEL1_14063_out0;
wire v$SEL1_14064_out0;
wire v$SEL1_14065_out0;
wire v$SEL1_14066_out0;
wire v$SEL1_14067_out0;
wire v$SEL1_14068_out0;
wire v$SEL1_14069_out0;
wire v$SEL1_14070_out0;
wire v$SEL1_14071_out0;
wire v$SEL1_14072_out0;
wire v$SEL1_14073_out0;
wire v$SEL1_14074_out0;
wire v$SEL1_14075_out0;
wire v$SEL1_14076_out0;
wire v$SEL1_14077_out0;
wire v$SEL1_14078_out0;
wire v$SEL1_14079_out0;
wire v$SEL1_1437_out0;
wire v$SEL1_1438_out0;
wire v$SEL1_18649_out0;
wire v$SEL1_18650_out0;
wire v$SEL1_18651_out0;
wire v$SEL1_18652_out0;
wire v$SEL1_2475_out0;
wire v$SEL1_2476_out0;
wire v$SEL1_2477_out0;
wire v$SEL1_2478_out0;
wire v$SEL1_2479_out0;
wire v$SEL1_2480_out0;
wire v$SEL1_2481_out0;
wire v$SEL1_2482_out0;
wire v$SEL1_3901_out0;
wire v$SEL1_3902_out0;
wire v$SEL1_7288_out0;
wire v$SEL1_7378_out0;
wire v$SEL1_7379_out0;
wire v$SEL1_7380_out0;
wire v$SEL1_7381_out0;
wire v$SEL20_8483_out0;
wire v$SEL20_8484_out0;
wire v$SEL20_8485_out0;
wire v$SEL20_8486_out0;
wire v$SEL21_11560_out0;
wire v$SEL21_11561_out0;
wire v$SEL21_11562_out0;
wire v$SEL21_11563_out0;
wire v$SEL22_7712_out0;
wire v$SEL22_7713_out0;
wire v$SEL22_7714_out0;
wire v$SEL22_7715_out0;
wire v$SEL23_7945_out0;
wire v$SEL23_7946_out0;
wire v$SEL23_7947_out0;
wire v$SEL23_7948_out0;
wire v$SEL24_17529_out0;
wire v$SEL24_17530_out0;
wire v$SEL24_17531_out0;
wire v$SEL24_17532_out0;
wire v$SEL27_16918_out0;
wire v$SEL27_16919_out0;
wire v$SEL27_16920_out0;
wire v$SEL27_16921_out0;
wire v$SEL28_7645_out0;
wire v$SEL28_7646_out0;
wire v$SEL28_7647_out0;
wire v$SEL28_7648_out0;
wire v$SEL29_17214_out0;
wire v$SEL29_17215_out0;
wire v$SEL29_17216_out0;
wire v$SEL29_17217_out0;
wire v$SEL2_13906_out0;
wire v$SEL2_13907_out0;
wire v$SEL2_13908_out0;
wire v$SEL2_13909_out0;
wire v$SEL2_14017_out0;
wire v$SEL2_14018_out0;
wire v$SEL2_16440_out0;
wire v$SEL2_17220_out0;
wire v$SEL2_17221_out0;
wire v$SEL2_17222_out0;
wire v$SEL2_17223_out0;
wire v$SEL2_17224_out0;
wire v$SEL2_17225_out0;
wire v$SEL2_17226_out0;
wire v$SEL2_17227_out0;
wire v$SEL2_17228_out0;
wire v$SEL2_17229_out0;
wire v$SEL2_17230_out0;
wire v$SEL2_17231_out0;
wire v$SEL2_17232_out0;
wire v$SEL2_17233_out0;
wire v$SEL2_17234_out0;
wire v$SEL2_17235_out0;
wire v$SEL2_17236_out0;
wire v$SEL2_17237_out0;
wire v$SEL2_17238_out0;
wire v$SEL2_17239_out0;
wire v$SEL2_17240_out0;
wire v$SEL2_17241_out0;
wire v$SEL2_17242_out0;
wire v$SEL2_17243_out0;
wire v$SEL2_18960_out0;
wire v$SEL2_18961_out0;
wire v$SEL2_18962_out0;
wire v$SEL2_18963_out0;
wire v$SEL2_18964_out0;
wire v$SEL2_18965_out0;
wire v$SEL2_18966_out0;
wire v$SEL2_18967_out0;
wire v$SEL2_19113_out0;
wire v$SEL2_19114_out0;
wire v$SEL2_19115_out0;
wire v$SEL2_19116_out0;
wire v$SEL2_3895_out0;
wire v$SEL2_3896_out0;
wire v$SEL2_7999_out0;
wire v$SEL2_8000_out0;
wire v$SEL2_8001_out0;
wire v$SEL2_8002_out0;
wire v$SEL2_8003_out0;
wire v$SEL2_8004_out0;
wire v$SEL2_8005_out0;
wire v$SEL2_8006_out0;
wire v$SEL2_8007_out0;
wire v$SEL2_8008_out0;
wire v$SEL2_8009_out0;
wire v$SEL2_8010_out0;
wire v$SEL2_8011_out0;
wire v$SEL2_8012_out0;
wire v$SEL2_8013_out0;
wire v$SEL2_8014_out0;
wire v$SEL2_8015_out0;
wire v$SEL2_8016_out0;
wire v$SEL2_8017_out0;
wire v$SEL2_8018_out0;
wire v$SEL2_8019_out0;
wire v$SEL2_8020_out0;
wire v$SEL2_8021_out0;
wire v$SEL2_8022_out0;
wire v$SEL2_8023_out0;
wire v$SEL2_8024_out0;
wire v$SEL2_8025_out0;
wire v$SEL2_8026_out0;
wire v$SEL2_8027_out0;
wire v$SEL2_8028_out0;
wire v$SEL2_8029_out0;
wire v$SEL2_8030_out0;
wire v$SEL2_8031_out0;
wire v$SEL2_8032_out0;
wire v$SEL2_8033_out0;
wire v$SEL2_8034_out0;
wire v$SEL2_9803_out0;
wire v$SEL2_9804_out0;
wire v$SEL3_12298_out0;
wire v$SEL3_12299_out0;
wire v$SEL3_12300_out0;
wire v$SEL3_12301_out0;
wire v$SEL3_1281_out0;
wire v$SEL3_1282_out0;
wire v$SEL3_1283_out0;
wire v$SEL3_1284_out0;
wire v$SEL3_1285_out0;
wire v$SEL3_1286_out0;
wire v$SEL3_1287_out0;
wire v$SEL3_1288_out0;
wire v$SEL3_14614_out0;
wire v$SEL3_14615_out0;
wire v$SEL3_14616_out0;
wire v$SEL3_14617_out0;
wire v$SEL3_18044_out0;
wire v$SEL3_18045_out0;
wire v$SEL3_19268_out0;
wire v$SEL3_19269_out0;
wire v$SEL3_2499_out0;
wire v$SEL3_2500_out0;
wire v$SEL3_2501_out0;
wire v$SEL3_2502_out0;
wire v$SEL3_2503_out0;
wire v$SEL3_2504_out0;
wire v$SEL3_2505_out0;
wire v$SEL3_2506_out0;
wire v$SEL3_2507_out0;
wire v$SEL3_2508_out0;
wire v$SEL3_2509_out0;
wire v$SEL3_2510_out0;
wire v$SEL3_2511_out0;
wire v$SEL3_2512_out0;
wire v$SEL3_2513_out0;
wire v$SEL3_2514_out0;
wire v$SEL3_2515_out0;
wire v$SEL3_2516_out0;
wire v$SEL3_2517_out0;
wire v$SEL3_2518_out0;
wire v$SEL3_2519_out0;
wire v$SEL3_2520_out0;
wire v$SEL3_2521_out0;
wire v$SEL3_2522_out0;
wire v$SEL3_2523_out0;
wire v$SEL3_2524_out0;
wire v$SEL3_2525_out0;
wire v$SEL3_2526_out0;
wire v$SEL3_2527_out0;
wire v$SEL3_2528_out0;
wire v$SEL3_2529_out0;
wire v$SEL3_2530_out0;
wire v$SEL3_2531_out0;
wire v$SEL3_2532_out0;
wire v$SEL3_2533_out0;
wire v$SEL3_2534_out0;
wire v$SEL3_3340_out0;
wire v$SEL3_8730_out0;
wire v$SEL3_8731_out0;
wire v$SEL3_8732_out0;
wire v$SEL3_8733_out0;
wire v$SEL3_8734_out0;
wire v$SEL3_8735_out0;
wire v$SEL3_8736_out0;
wire v$SEL3_8737_out0;
wire v$SEL3_8738_out0;
wire v$SEL3_8739_out0;
wire v$SEL3_8740_out0;
wire v$SEL3_8741_out0;
wire v$SEL3_8742_out0;
wire v$SEL3_8743_out0;
wire v$SEL3_8744_out0;
wire v$SEL3_8745_out0;
wire v$SEL3_8746_out0;
wire v$SEL3_8747_out0;
wire v$SEL3_8748_out0;
wire v$SEL3_8749_out0;
wire v$SEL3_8750_out0;
wire v$SEL3_8751_out0;
wire v$SEL3_8752_out0;
wire v$SEL3_8753_out0;
wire v$SEL4_17042_out0;
wire v$SEL4_2005_out0;
wire v$SEL4_2006_out0;
wire v$SEL4_2007_out0;
wire v$SEL4_2008_out0;
wire v$SEL4_5152_out0;
wire v$SEL4_5153_out0;
wire v$SEL4_5154_out0;
wire v$SEL4_5155_out0;
wire v$SEL4_5156_out0;
wire v$SEL4_5157_out0;
wire v$SEL4_5158_out0;
wire v$SEL4_5159_out0;
wire v$SEL4_6356_out0;
wire v$SEL4_6357_out0;
wire v$SEL4_6358_out0;
wire v$SEL4_6359_out0;
wire v$SEL4_6360_out0;
wire v$SEL4_6361_out0;
wire v$SEL4_6362_out0;
wire v$SEL4_6363_out0;
wire v$SEL4_6364_out0;
wire v$SEL4_6365_out0;
wire v$SEL4_6366_out0;
wire v$SEL4_6367_out0;
wire v$SEL4_6368_out0;
wire v$SEL4_6369_out0;
wire v$SEL4_6370_out0;
wire v$SEL4_6371_out0;
wire v$SEL4_6372_out0;
wire v$SEL4_6373_out0;
wire v$SEL4_6374_out0;
wire v$SEL4_6375_out0;
wire v$SEL4_6376_out0;
wire v$SEL4_6377_out0;
wire v$SEL4_6378_out0;
wire v$SEL4_6379_out0;
wire v$SEL4_6380_out0;
wire v$SEL4_6381_out0;
wire v$SEL4_6382_out0;
wire v$SEL4_6383_out0;
wire v$SEL4_6384_out0;
wire v$SEL4_6385_out0;
wire v$SEL4_6386_out0;
wire v$SEL4_6387_out0;
wire v$SEL4_6388_out0;
wire v$SEL4_6389_out0;
wire v$SEL4_6390_out0;
wire v$SEL4_6391_out0;
wire v$SEL4_7339_out0;
wire v$SEL4_7340_out0;
wire v$SEL4_7639_out0;
wire v$SEL4_7640_out0;
wire v$SEL4_7641_out0;
wire v$SEL4_7642_out0;
wire v$SEL4_7652_out0;
wire v$SEL4_7653_out0;
wire v$SEL4_7654_out0;
wire v$SEL4_7655_out0;
wire v$SEL4_7656_out0;
wire v$SEL4_7657_out0;
wire v$SEL4_7658_out0;
wire v$SEL4_7659_out0;
wire v$SEL4_7660_out0;
wire v$SEL4_7661_out0;
wire v$SEL4_7662_out0;
wire v$SEL4_7663_out0;
wire v$SEL4_7664_out0;
wire v$SEL4_7665_out0;
wire v$SEL4_7666_out0;
wire v$SEL4_7667_out0;
wire v$SEL4_7668_out0;
wire v$SEL4_7669_out0;
wire v$SEL4_7670_out0;
wire v$SEL4_7671_out0;
wire v$SEL4_7672_out0;
wire v$SEL4_7673_out0;
wire v$SEL4_7674_out0;
wire v$SEL4_7675_out0;
wire v$SEL5_12186_out0;
wire v$SEL5_12232_out0;
wire v$SEL5_12233_out0;
wire v$SEL5_12234_out0;
wire v$SEL5_12235_out0;
wire v$SEL5_12781_out0;
wire v$SEL5_12782_out0;
wire v$SEL5_12783_out0;
wire v$SEL5_12784_out0;
wire v$SEL5_12785_out0;
wire v$SEL5_12786_out0;
wire v$SEL5_12787_out0;
wire v$SEL5_12788_out0;
wire v$SEL5_13345_out0;
wire v$SEL5_13346_out0;
wire v$SEL5_13347_out0;
wire v$SEL5_13348_out0;
wire v$SEL5_13349_out0;
wire v$SEL5_13350_out0;
wire v$SEL5_13351_out0;
wire v$SEL5_13352_out0;
wire v$SEL5_13353_out0;
wire v$SEL5_13354_out0;
wire v$SEL5_13355_out0;
wire v$SEL5_13356_out0;
wire v$SEL5_13357_out0;
wire v$SEL5_13358_out0;
wire v$SEL5_13359_out0;
wire v$SEL5_13360_out0;
wire v$SEL5_13361_out0;
wire v$SEL5_13362_out0;
wire v$SEL5_13363_out0;
wire v$SEL5_13364_out0;
wire v$SEL5_13365_out0;
wire v$SEL5_13366_out0;
wire v$SEL5_13367_out0;
wire v$SEL5_13368_out0;
wire v$SEL5_16038_out0;
wire v$SEL5_16039_out0;
wire v$SEL5_16040_out0;
wire v$SEL5_16041_out0;
wire v$SEL5_326_out0;
wire v$SEL5_327_out0;
wire v$SEL6_13066_out0;
wire v$SEL6_13067_out0;
wire v$SEL6_13068_out0;
wire v$SEL6_13069_out0;
wire v$SEL6_14365_out0;
wire v$SEL6_14366_out0;
wire v$SEL6_14367_out0;
wire v$SEL6_14368_out0;
wire v$SEL6_14369_out0;
wire v$SEL6_14370_out0;
wire v$SEL6_14371_out0;
wire v$SEL6_14372_out0;
wire v$SEL6_14846_out0;
wire v$SEL6_15060_out0;
wire v$SEL6_15061_out0;
wire v$SEL6_6092_out0;
wire v$SEL6_6093_out0;
wire v$SEL6_6094_out0;
wire v$SEL6_6095_out0;
wire v$SEL7_14936_out0;
wire v$SEL7_14937_out0;
wire v$SEL7_14938_out0;
wire v$SEL7_14939_out0;
wire v$SEL7_16208_out0;
wire v$SEL7_16209_out0;
wire v$SEL7_17604_out0;
wire v$SEL7_4324_out0;
wire v$SEL7_4325_out0;
wire v$SEL7_4326_out0;
wire v$SEL7_4327_out0;
wire v$SEL7_4328_out0;
wire v$SEL7_4329_out0;
wire v$SEL7_4330_out0;
wire v$SEL7_4331_out0;
wire v$SEL7_4332_out0;
wire v$SEL7_4333_out0;
wire v$SEL7_4334_out0;
wire v$SEL7_4335_out0;
wire v$SEL7_4336_out0;
wire v$SEL7_4337_out0;
wire v$SEL7_4338_out0;
wire v$SEL7_4339_out0;
wire v$SEL7_4340_out0;
wire v$SEL7_4341_out0;
wire v$SEL7_4342_out0;
wire v$SEL7_4343_out0;
wire v$SEL7_4344_out0;
wire v$SEL7_4345_out0;
wire v$SEL7_4346_out0;
wire v$SEL7_4347_out0;
wire v$SEL7_6596_out0;
wire v$SEL7_6597_out0;
wire v$SEL7_6598_out0;
wire v$SEL7_6599_out0;
wire v$SEL7_6600_out0;
wire v$SEL7_6601_out0;
wire v$SEL7_6602_out0;
wire v$SEL7_6603_out0;
wire v$SEL8_13484_out0;
wire v$SEL8_13485_out0;
wire v$SEL8_13486_out0;
wire v$SEL8_13487_out0;
wire v$SEL8_13488_out0;
wire v$SEL8_13489_out0;
wire v$SEL8_13490_out0;
wire v$SEL8_13491_out0;
wire v$SEL8_13492_out0;
wire v$SEL8_13493_out0;
wire v$SEL8_13494_out0;
wire v$SEL8_13495_out0;
wire v$SEL8_13496_out0;
wire v$SEL8_13497_out0;
wire v$SEL8_13498_out0;
wire v$SEL8_13499_out0;
wire v$SEL8_13500_out0;
wire v$SEL8_13501_out0;
wire v$SEL8_13502_out0;
wire v$SEL8_13503_out0;
wire v$SEL8_13504_out0;
wire v$SEL8_13505_out0;
wire v$SEL8_13506_out0;
wire v$SEL8_13507_out0;
wire v$SEL8_17190_out0;
wire v$SEL8_17191_out0;
wire v$SEL8_17192_out0;
wire v$SEL8_17193_out0;
wire v$SEL8_17194_out0;
wire v$SEL8_17195_out0;
wire v$SEL8_17196_out0;
wire v$SEL8_17197_out0;
wire v$SEL8_18285_out0;
wire v$SEL8_18286_out0;
wire v$SEL8_18287_out0;
wire v$SEL8_18288_out0;
wire v$SEL8_2132_out0;
wire v$SEL9_10717_out0;
wire v$SEL9_10718_out0;
wire v$SEL9_10719_out0;
wire v$SEL9_10720_out0;
wire v$SEL9_11336_out0;
wire v$SEL9_11337_out0;
wire v$SEL9_11338_out0;
wire v$SEL9_11339_out0;
wire v$SEL9_11340_out0;
wire v$SEL9_11341_out0;
wire v$SEL9_11342_out0;
wire v$SEL9_11343_out0;
wire v$SEL9_11344_out0;
wire v$SEL9_11345_out0;
wire v$SEL9_11346_out0;
wire v$SEL9_11347_out0;
wire v$SEL9_11348_out0;
wire v$SEL9_11349_out0;
wire v$SEL9_11350_out0;
wire v$SEL9_11351_out0;
wire v$SEL9_11352_out0;
wire v$SEL9_11353_out0;
wire v$SEL9_11354_out0;
wire v$SEL9_11355_out0;
wire v$SEL9_11356_out0;
wire v$SEL9_11357_out0;
wire v$SEL9_11358_out0;
wire v$SEL9_11359_out0;
wire v$SELIN$VIEWER_11583_out0;
wire v$SELIN_18816_out0;
wire v$SELOUTVIEWER_7596_out0;
wire v$SELOUT_1880_out0;
wire v$SERIALIN_6011_out0;
wire v$SERIALIN_6012_out0;
wire v$SHIFTEN_10737_out0;
wire v$SHIFTEN_10738_out0;
wire v$SHIFTEN_13335_out0;
wire v$SHIFTEN_13336_out0;
wire v$SHIFTEN_7382_out0;
wire v$SHIFTEN_7383_out0;
wire v$SHIFTEN_9781_out0;
wire v$SHIFTEN_9782_out0;
wire v$SHIFTEN_9783_out0;
wire v$SHIFTEN_9784_out0;
wire v$SHIFTEN_9785_out0;
wire v$SHIFTEN_9786_out0;
wire v$SHIFTEN_9787_out0;
wire v$SHIFTEN_9788_out0;
wire v$SHIFTEN_9789_out0;
wire v$SHIFTEN_9790_out0;
wire v$SHIFTEN_9791_out0;
wire v$SHIFTEN_9792_out0;
wire v$SHOULD$STORE_13280_out0;
wire v$SHOULD$STORE_13281_out0;
wire v$SIGN_13329_out0;
wire v$SIGN_13330_out0;
wire v$SIGN_1529_out0;
wire v$SIGN_1530_out0;
wire v$SIGN_1531_out0;
wire v$SIGN_1532_out0;
wire v$SIN_100_out0;
wire v$SIN_101_out0;
wire v$SIN_102_out0;
wire v$SIN_103_out0;
wire v$SIN_92_out0;
wire v$SIN_93_out0;
wire v$SIN_94_out0;
wire v$SIN_95_out0;
wire v$SIN_96_out0;
wire v$SIN_97_out0;
wire v$SIN_98_out0;
wire v$SIN_99_out0;
wire v$SOUT1_2080_out0;
wire v$SOUT1_2081_out0;
wire v$SOUT1_2082_out0;
wire v$SOUT1_2083_out0;
wire v$SOUT1_2084_out0;
wire v$SOUT1_2085_out0;
wire v$SOUT1_2086_out0;
wire v$SOUT1_2087_out0;
wire v$SOUT1_2088_out0;
wire v$SOUT1_2089_out0;
wire v$SOUT1_2090_out0;
wire v$SOUT1_2091_out0;
wire v$SOUT_18793_out0;
wire v$SOUT_18794_out0;
wire v$STALL$FETCH$OCCURRED_2844_out0;
wire v$STALL$FETCH$OCCURRED_2845_out0;
wire v$STALL$IN$PREV_13795_out0;
wire v$STALL$IN$PREV_13796_out0;
wire v$STALL$PREV$CYCLE_6059_out0;
wire v$STALL$PREV$CYCLE_6060_out0;
wire v$STALL$PREV$PREV_6096_out0;
wire v$STALL$PREV$PREV_6097_out0;
wire v$STALL$VIEWER_18671_out0;
wire v$STALL$VIEWER_18672_out0;
wire v$STALL_12797_out0;
wire v$STALL_12798_out0;
wire v$STALL_13723_out0;
wire v$STALL_13724_out0;
wire v$STALL_16085_out0;
wire v$STALL_16086_out0;
wire v$STALL_18502_out0;
wire v$STALL_18503_out0;
wire v$START$PIPELINED$VIEWER_6640_out0;
wire v$START$PIPELINED$VIEWER_6641_out0;
wire v$START_14620_out0;
wire v$START_14621_out0;
wire v$START_16968_out0;
wire v$START_16969_out0;
wire v$START_19327_out0;
wire v$START_19328_out0;
wire v$START_3879_out0;
wire v$START_3880_out0;
wire v$START_4398_out0;
wire v$START_4399_out0;
wire v$START_5733_out0;
wire v$START_5734_out0;
wire v$STATE_16624_out0;
wire v$STATE_16625_out0;
wire v$STATE_16626_out0;
wire v$STATE_16627_out0;
wire v$STATE_16628_out0;
wire v$STATE_16629_out0;
wire v$STATE_16630_out0;
wire v$STATUSCLR_6234_out0;
wire v$STATUSCLR_6235_out0;
wire v$STATUSREAD_1795_out0;
wire v$STATUSREAD_1796_out0;
wire v$STClr_10669_out0;
wire v$STClr_10670_out0;
wire v$STOP$1_8134_out0;
wire v$STOP$1_8135_out0;
wire v$STOP$2_8543_out0;
wire v$STOP$2_8544_out0;
wire v$STOPBITERROR_12296_out0;
wire v$STOPBITERROR_12297_out0;
wire v$STOPERROR_306_out0;
wire v$STOPERROR_307_out0;
wire v$STP$DECODED_17154_out0;
wire v$STP$DECODED_17155_out0;
wire v$STP$SAVED_7884_out0;
wire v$STP$SAVED_7885_out0;
wire v$STPHALT_13514_out0;
wire v$STPHALT_13515_out0;
wire v$STPHALT_18735_out0;
wire v$STPHALT_18736_out0;
wire v$STPHALT_4478_out0;
wire v$STPHALT_4479_out0;
wire v$STP_11314_out0;
wire v$STP_11315_out0;
wire v$STP_12282_out0;
wire v$STP_12283_out0;
wire v$STP_18374_out0;
wire v$STP_18375_out0;
wire v$STP_6467_out0;
wire v$STP_6468_out0;
wire v$STRead_10348_out0;
wire v$STRead_10349_out0;
wire v$SUBEN_13429_out0;
wire v$SUBEN_13430_out0;
wire v$SUBTRACTION$SIGN_12445_out0;
wire v$SUBTRACTION$SIGN_12446_out0;
wire v$SUB_14377_out0;
wire v$SUB_14378_out0;
wire v$S_1004_out0;
wire v$S_1005_out0;
wire v$S_10809_out0;
wire v$S_10810_out0;
wire v$S_10894_out0;
wire v$S_10895_out0;
wire v$S_11196_out0;
wire v$S_11197_out0;
wire v$S_13233_out0;
wire v$S_13234_out0;
wire v$S_13389_out0;
wire v$S_13390_out0;
wire v$S_1377_out0;
wire v$S_16062_out0;
wire v$S_16063_out0;
wire v$S_16064_out0;
wire v$S_16065_out0;
wire v$S_16066_out0;
wire v$S_16067_out0;
wire v$S_17002_out0;
wire v$S_17003_out0;
wire v$S_17537_out0;
wire v$S_17538_out0;
wire v$S_17539_out0;
wire v$S_17540_out0;
wire v$S_17541_out0;
wire v$S_17542_out0;
wire v$S_17543_out0;
wire v$S_17544_out0;
wire v$S_17545_out0;
wire v$S_17546_out0;
wire v$S_17547_out0;
wire v$S_17548_out0;
wire v$S_17549_out0;
wire v$S_17550_out0;
wire v$S_17551_out0;
wire v$S_17552_out0;
wire v$S_17553_out0;
wire v$S_17554_out0;
wire v$S_17555_out0;
wire v$S_17556_out0;
wire v$S_17557_out0;
wire v$S_17558_out0;
wire v$S_18561_out0;
wire v$S_18562_out0;
wire v$S_2636_out0;
wire v$S_2637_out0;
wire v$S_4182_out0;
wire v$S_4183_out0;
wire v$S_4400_out0;
wire v$S_4401_out0;
wire v$S_6017_out0;
wire v$S_6018_out0;
wire v$S_8335_out0;
wire v$S_8336_out0;
wire v$S_8337_out0;
wire v$S_8338_out0;
wire v$S_8339_out0;
wire v$S_8340_out0;
wire v$S_8341_out0;
wire v$S_8475_out0;
wire v$S_8476_out0;
wire v$S_9799_out0;
wire v$S_9800_out0;
wire v$SetError_18196_out0;
wire v$SetError_18197_out0;
wire v$ShiftEN_6115_out0;
wire v$ShiftEN_6116_out0;
wire v$ShiftEN_8039_out0;
wire v$ShiftEN_8040_out0;
wire v$ShiftOut_16960_out0;
wire v$ShiftOut_16961_out0;
wire v$Shift_9986_out0;
wire v$Shift_9987_out0;
wire v$StatRegAdd1_15154_out0;
wire v$StatRegAdd1_15155_out0;
wire v$StatRegAdd_8059_out0;
wire v$StatRegAdd_8060_out0;
wire v$TAKEJUMP_11294_out0;
wire v$TAKEJUMP_11295_out0;
wire v$THRESHOLD$WRITE_7550_out0;
wire v$THRESHOLD$WRITE_7551_out0;
wire v$TWOS$COMPLEMENT$ADDER$COUT_3639_out0;
wire v$TWOS$COMPLEMENT$ADDER$COUT_3640_out0;
wire v$TXFLAG_15295_out0;
wire v$TXFLAG_15296_out0;
wire v$TXFLAG_4060_out0;
wire v$TXFLAG_4061_out0;
wire v$TXFlag_15829_out0;
wire v$TXFlag_15830_out0;
wire v$TXFlag_8035_out0;
wire v$TXFlag_8036_out0;
wire v$TXINTERRUPT_3824_out0;
wire v$TXINTERRUPT_3825_out0;
wire v$TXINT_5126_out0;
wire v$TXINT_5127_out0;
wire v$TXLast_11914_out0;
wire v$TXLast_11915_out0;
wire v$TXRST_16998_out0;
wire v$TXRST_16999_out0;
wire v$TXRST_8358_out0;
wire v$TXRST_8359_out0;
wire v$TXRegAdd_16193_out0;
wire v$TXRegAdd_16194_out0;
wire v$TXReset_18441_out0;
wire v$TXReset_18442_out0;
wire v$TXSet_13235_out0;
wire v$TXSet_13236_out0;
wire v$TXSet_14941_out0;
wire v$TXSet_14942_out0;
wire v$TXWRITE_11608_out0;
wire v$TXWRITE_11609_out0;
wire v$TXWRITE_16703_out0;
wire v$TXWRITE_16704_out0;
wire v$TXWrite_18136_out0;
wire v$TXWrite_18137_out0;
wire v$TX_12248_out0;
wire v$TX_12249_out0;
wire v$TX_1458_out0;
wire v$TX_1459_out0;
wire v$TX_18860_out0;
wire v$TX_18861_out0;
wire v$TX_439_out0;
wire v$TX_440_out0;
wire v$TXoverflow_4265_out0;
wire v$TXoverflow_4266_out0;
wire v$V0_7741_out0;
wire v$V0_9720_out0;
wire v$V1_17321_out0;
wire v$V1_18443_out0;
wire v$VALID$PREV_14013_out0;
wire v$VALID$PREV_14014_out0;
wire v$VALID0_13990_out0;
wire v$VALID1_9151_out0;
wire v$VALID_15094_out0;
wire v$VALID_15095_out0;
wire v$VALID_18531_out0;
wire v$VALID_18532_out0;
wire v$VALID_19282_out0;
wire v$VALID_19283_out0;
wire v$VALID_3893_out0;
wire v$VALID_3894_out0;
wire v$WB$HAZARD_9227_out0;
wire v$WB$HAZARD_9228_out0;
wire v$WEN$FPU_8623_out0;
wire v$WEN$FPU_8624_out0;
wire v$WEN3_2009_out0;
wire v$WEN3_2010_out0;
wire v$WEN3_3509_out0;
wire v$WEN3_3510_out0;
wire v$WENALU_16990_out0;
wire v$WENALU_16991_out0;
wire v$WENALU_19270_out0;
wire v$WENALU_19271_out0;
wire v$WENALU_4228_out0;
wire v$WENALU_4229_out0;
wire v$WENFPU_14322_out0;
wire v$WENFPU_14323_out0;
wire v$WENFPU_3698_out0;
wire v$WENFPU_3699_out0;
wire v$WENLDST_13078_out0;
wire v$WENLDST_13079_out0;
wire v$WENLDST_19239_out0;
wire v$WENLDST_19240_out0;
wire v$WENLDST_6924_out0;
wire v$WENLDST_6925_out0;
wire v$WENRAM0_10341_out0;
wire v$WENRAM1_1879_out0;
wire v$WENRAM_17680_out0;
wire v$WENRAM_17681_out0;
wire v$WENRAM_2535_out0;
wire v$WENRAM_2536_out0;
wire v$WENRAM_5184_out0;
wire v$WENRAM_5185_out0;
wire v$WEN_12738_out0;
wire v$WEN_12739_out0;
wire v$WEN_12900_out0;
wire v$WEN_12901_out0;
wire v$WEN_14820_out0;
wire v$WEN_14821_out0;
wire v$WEN_18998_out0;
wire v$WEN_18999_out0;
wire v$WEN_3862_out0;
wire v$WEN_3863_out0;
wire v$WEN_3983_out0;
wire v$WEN_3984_out0;
wire v$WR0VIEWER_16495_out0;
wire v$WR0_1478_out0;
wire v$WR0_14871_out0;
wire v$WR1VIEWER_16508_out0;
wire v$WR1_14940_out0;
wire v$WR1_315_out0;
wire v$WREN_11505_out0;
wire v$WREN_11506_out0;
wire v$WREN_2730_out0;
wire v$WREN_2731_out0;
wire v$Wordlength_5358_out0;
wire v$Wordlength_5359_out0;
wire v$Write_3479_out0;
wire v$Write_3480_out0;
wire v$Write_3481_out0;
wire v$Write_3482_out0;
wire v$Write_3483_out0;
wire v$Write_3484_out0;
wire v$Write_3485_out0;
wire v$Write_3486_out0;
wire v$Write_3487_out0;
wire v$Write_3488_out0;
wire v$Write_3489_out0;
wire v$Write_3490_out0;
wire v$Z1_17592_out0;
wire v$Z1_17593_out0;
wire v$Z1_17594_out0;
wire v$Z1_17595_out0;
wire v$Z1_17596_out0;
wire v$Z1_17597_out0;
wire v$Z1_17598_out0;
wire v$Z1_17599_out0;
wire v$Z1_18330_out0;
wire v$Z1_18331_out0;
wire v$Z1_6049_out0;
wire v$Z1_6050_out0;
wire v$Z1_6051_out0;
wire v$Z1_6052_out0;
wire v$Z1_6053_out0;
wire v$Z1_6054_out0;
wire v$Z1_6055_out0;
wire v$Z1_6056_out0;
wire v$Z1_6057_out0;
wire v$Z1_6058_out0;
wire v$Z2_180_out0;
wire v$Z2_181_out0;
wire v$Z2_182_out0;
wire v$Z2_183_out0;
wire v$Z2_184_out0;
wire v$Z2_185_out0;
wire v$Z2_186_out0;
wire v$Z2_187_out0;
wire v$Z2_188_out0;
wire v$Z2_189_out0;
wire v$Z2_2463_out0;
wire v$Z2_2464_out0;
wire v$Z2_6574_out0;
wire v$Z2_6575_out0;
wire v$Z2_6576_out0;
wire v$Z2_6577_out0;
wire v$Z2_6578_out0;
wire v$Z2_6579_out0;
wire v$Z2_6580_out0;
wire v$Z2_6581_out0;
wire v$Z3_12563_out0;
wire v$Z3_12564_out0;
wire v$Z3_18389_out0;
wire v$Z3_18390_out0;
wire v$Z3_18391_out0;
wire v$Z3_18392_out0;
wire v$Z4_8247_out0;
wire v$Z4_8248_out0;
wire v$Z4_8249_out0;
wire v$Z4_8250_out0;
wire v$Z_10787_out0;
wire v$Z_10788_out0;
wire v$Z_10789_out0;
wire v$Z_10790_out0;
wire v$Z_10791_out0;
wire v$Z_10792_out0;
wire v$Z_10793_out0;
wire v$Z_10794_out0;
wire v$Z_10795_out0;
wire v$Z_10796_out0;
wire v$Z_13147_out0;
wire v$Z_13148_out0;
wire v$Z_13149_out0;
wire v$Z_13150_out0;
wire v$Z_13151_out0;
wire v$Z_13152_out0;
wire v$Z_13153_out0;
wire v$Z_13154_out0;
wire v$Z_13155_out0;
wire v$Z_13156_out0;
wire v$Z_13157_out0;
wire v$Z_13158_out0;
wire v$Z_13159_out0;
wire v$Z_13160_out0;
wire v$Z_13161_out0;
wire v$Z_13162_out0;
wire v$Z_13163_out0;
wire v$Z_13164_out0;
wire v$Z_13165_out0;
wire v$Z_13166_out0;
wire v$Z_13167_out0;
wire v$Z_13168_out0;
wire v$Z_13169_out0;
wire v$Z_13170_out0;
wire v$Z_13171_out0;
wire v$Z_13172_out0;
wire v$Z_13173_out0;
wire v$Z_13174_out0;
wire v$Z_13175_out0;
wire v$Z_13176_out0;
wire v$Z_13177_out0;
wire v$Z_13178_out0;
wire v$Z_13179_out0;
wire v$Z_13180_out0;
wire v$Z_13181_out0;
wire v$Z_13182_out0;
wire v$Z_14128_out0;
wire v$Z_14129_out0;
wire v$Z_16411_out0;
wire v$Z_16412_out0;
wire v$Z_16413_out0;
wire v$Z_16414_out0;
wire v$Z_2747_out0;
wire v$Z_2748_out0;
wire v$Z_2749_out0;
wire v$Z_2750_out0;
wire v$Z_2751_out0;
wire v$Z_2752_out0;
wire v$Z_2753_out0;
wire v$Z_2754_out0;
wire v$_10697_out0;
wire v$_10697_out1;
wire v$_10698_out0;
wire v$_10698_out1;
wire v$_10733_out0;
wire v$_10734_out0;
wire v$_10739_out0;
wire v$_10739_out1;
wire v$_10740_out0;
wire v$_10740_out1;
wire v$_10741_out0;
wire v$_10741_out1;
wire v$_10742_out0;
wire v$_10742_out1;
wire v$_10743_out0;
wire v$_10743_out1;
wire v$_10744_out0;
wire v$_10744_out1;
wire v$_10868_out0;
wire v$_10869_out0;
wire v$_10898_out0;
wire v$_10899_out0;
wire v$_10900_out0;
wire v$_10901_out0;
wire v$_10902_out0;
wire v$_10903_out0;
wire v$_11264_out0;
wire v$_11265_out0;
wire v$_11266_out0;
wire v$_11267_out0;
wire v$_11268_out0;
wire v$_11269_out0;
wire v$_11282_out0;
wire v$_11283_out0;
wire v$_11413_out0;
wire v$_11414_out0;
wire v$_11415_out0;
wire v$_11416_out0;
wire v$_11417_out0;
wire v$_11418_out0;
wire v$_11531_out0;
wire v$_11531_out1;
wire v$_11532_out0;
wire v$_11532_out1;
wire v$_11533_out0;
wire v$_11533_out1;
wire v$_11534_out0;
wire v$_11534_out1;
wire v$_11535_out0;
wire v$_11535_out1;
wire v$_11536_out0;
wire v$_11536_out1;
wire v$_11568_out0;
wire v$_11568_out1;
wire v$_11569_out0;
wire v$_11569_out1;
wire v$_11596_out0;
wire v$_11597_out0;
wire v$_11598_out0;
wire v$_11599_out0;
wire v$_11600_out0;
wire v$_11601_out0;
wire v$_11920_out0;
wire v$_11921_out0;
wire v$_12178_out0;
wire v$_12178_out1;
wire v$_12179_out0;
wire v$_12179_out1;
wire v$_12180_out0;
wire v$_12180_out1;
wire v$_12181_out0;
wire v$_12181_out1;
wire v$_12182_out0;
wire v$_12182_out1;
wire v$_12183_out0;
wire v$_12183_out1;
wire v$_12334_out0;
wire v$_12335_out0;
wire v$_12431_out0;
wire v$_12431_out1;
wire v$_12432_out0;
wire v$_12432_out1;
wire v$_12433_out0;
wire v$_12433_out1;
wire v$_12434_out0;
wire v$_12434_out1;
wire v$_12435_out0;
wire v$_12435_out1;
wire v$_12436_out0;
wire v$_12436_out1;
wire v$_12437_out0;
wire v$_12437_out1;
wire v$_12438_out0;
wire v$_12438_out1;
wire v$_12439_out0;
wire v$_12439_out1;
wire v$_12440_out0;
wire v$_12440_out1;
wire v$_12441_out0;
wire v$_12441_out1;
wire v$_12442_out0;
wire v$_12442_out1;
wire v$_12641_out0;
wire v$_12641_out1;
wire v$_12642_out0;
wire v$_12642_out1;
wire v$_12643_out0;
wire v$_12643_out1;
wire v$_12644_out0;
wire v$_12644_out1;
wire v$_13333_out0;
wire v$_13334_out0;
wire v$_13341_out0;
wire v$_13342_out0;
wire v$_1345_out0;
wire v$_1346_out0;
wire v$_13758_out0;
wire v$_13758_out1;
wire v$_13759_out0;
wire v$_13759_out1;
wire v$_13760_out0;
wire v$_13760_out1;
wire v$_13761_out0;
wire v$_13761_out1;
wire v$_13762_out0;
wire v$_13762_out1;
wire v$_13763_out0;
wire v$_13763_out1;
wire v$_13853_out0;
wire v$_13856_out0;
wire v$_13873_out0;
wire v$_13874_out0;
wire v$_14119_out0;
wire v$_14120_out0;
wire v$_14272_out0;
wire v$_14273_out0;
wire v$_14431_out0;
wire v$_14431_out1;
wire v$_14432_out0;
wire v$_14432_out1;
wire v$_1462_out0;
wire v$_1463_out0;
wire v$_1464_out0;
wire v$_1465_out0;
wire v$_1466_out0;
wire v$_1467_out0;
wire v$_14689_out0;
wire v$_14689_out1;
wire v$_14690_out0;
wire v$_14690_out1;
wire v$_14849_out0;
wire v$_14849_out1;
wire v$_14850_out0;
wire v$_14850_out1;
wire v$_14928_out0;
wire v$_14929_out0;
wire v$_15108_out0;
wire v$_15108_out1;
wire v$_15109_out0;
wire v$_15109_out1;
wire v$_15110_out0;
wire v$_15110_out1;
wire v$_15111_out0;
wire v$_15111_out1;
wire v$_15112_out0;
wire v$_15112_out1;
wire v$_15113_out0;
wire v$_15113_out1;
wire v$_15114_out0;
wire v$_15114_out1;
wire v$_15115_out0;
wire v$_15115_out1;
wire v$_15116_out0;
wire v$_15116_out1;
wire v$_15117_out0;
wire v$_15117_out1;
wire v$_15118_out0;
wire v$_15118_out1;
wire v$_15119_out0;
wire v$_15119_out1;
wire v$_15120_out0;
wire v$_15120_out1;
wire v$_15121_out0;
wire v$_15121_out1;
wire v$_1515_out0;
wire v$_1516_out0;
wire v$_1517_out0;
wire v$_1518_out0;
wire v$_1519_out0;
wire v$_1520_out0;
wire v$_15249_out0;
wire v$_15249_out1;
wire v$_15250_out0;
wire v$_15250_out1;
wire v$_15748_out0;
wire v$_15749_out0;
wire v$_15758_out0;
wire v$_15759_out0;
wire v$_15760_out0;
wire v$_15761_out0;
wire v$_15762_out0;
wire v$_15763_out0;
wire v$_15786_out0;
wire v$_15786_out1;
wire v$_15787_out0;
wire v$_15787_out1;
wire v$_15788_out0;
wire v$_15788_out1;
wire v$_15789_out0;
wire v$_15789_out1;
wire v$_15905_out0;
wire v$_15905_out1;
wire v$_15906_out0;
wire v$_15906_out1;
wire v$_16339_out0;
wire v$_16339_out1;
wire v$_16340_out0;
wire v$_16340_out1;
wire v$_16341_out0;
wire v$_16341_out1;
wire v$_16342_out0;
wire v$_16342_out1;
wire v$_16343_out0;
wire v$_16343_out1;
wire v$_16344_out0;
wire v$_16344_out1;
wire v$_16443_out0;
wire v$_16443_out1;
wire v$_16444_out0;
wire v$_16444_out1;
wire v$_16742_out0;
wire v$_16743_out0;
wire v$_16744_out0;
wire v$_16745_out0;
wire v$_16746_out0;
wire v$_16747_out0;
wire v$_16750_out0;
wire v$_16750_out1;
wire v$_16751_out0;
wire v$_16751_out1;
wire v$_16791_out0;
wire v$_16791_out1;
wire v$_16792_out0;
wire v$_16792_out1;
wire v$_16793_out0;
wire v$_16793_out1;
wire v$_16794_out0;
wire v$_16794_out1;
wire v$_16795_out0;
wire v$_16795_out1;
wire v$_16796_out0;
wire v$_16796_out1;
wire v$_16876_out0;
wire v$_16877_out0;
wire v$_16878_out0;
wire v$_16879_out0;
wire v$_16880_out0;
wire v$_16881_out0;
wire v$_1709_out0;
wire v$_1710_out0;
wire v$_17170_out0;
wire v$_17170_out1;
wire v$_17171_out0;
wire v$_17171_out1;
wire v$_17208_out0;
wire v$_17208_out1;
wire v$_17209_out0;
wire v$_17209_out1;
wire v$_17210_out0;
wire v$_17210_out1;
wire v$_17211_out0;
wire v$_17211_out1;
wire v$_17212_out0;
wire v$_17212_out1;
wire v$_17213_out0;
wire v$_17213_out1;
wire v$_17322_out0;
wire v$_17322_out1;
wire v$_17323_out0;
wire v$_17323_out1;
wire v$_17324_out0;
wire v$_17324_out1;
wire v$_17325_out0;
wire v$_17325_out1;
wire v$_17326_out0;
wire v$_17326_out1;
wire v$_17327_out0;
wire v$_17327_out1;
wire v$_17361_out0;
wire v$_17362_out0;
wire v$_17363_out0;
wire v$_17364_out0;
wire v$_17365_out0;
wire v$_17366_out0;
wire v$_17577_out0;
wire v$_17577_out1;
wire v$_17578_out0;
wire v$_17578_out1;
wire v$_17965_out0;
wire v$_17965_out1;
wire v$_17966_out0;
wire v$_17966_out1;
wire v$_17967_out0;
wire v$_17967_out1;
wire v$_17968_out0;
wire v$_17968_out1;
wire v$_17969_out0;
wire v$_17969_out1;
wire v$_17970_out0;
wire v$_17970_out1;
wire v$_1797_out0;
wire v$_1797_out1;
wire v$_1798_out0;
wire v$_1798_out1;
wire v$_1799_out0;
wire v$_1799_out1;
wire v$_1800_out0;
wire v$_1800_out1;
wire v$_1801_out0;
wire v$_1801_out1;
wire v$_1802_out0;
wire v$_1802_out1;
wire v$_1803_out0;
wire v$_1803_out1;
wire v$_1804_out0;
wire v$_1804_out1;
wire v$_1805_out0;
wire v$_1805_out1;
wire v$_1806_out0;
wire v$_1806_out1;
wire v$_1807_out0;
wire v$_1807_out1;
wire v$_1808_out0;
wire v$_1808_out1;
wire v$_18366_out0;
wire v$_18366_out1;
wire v$_18367_out0;
wire v$_18367_out1;
wire v$_18368_out0;
wire v$_18368_out1;
wire v$_18369_out0;
wire v$_18369_out1;
wire v$_18370_out0;
wire v$_18370_out1;
wire v$_18371_out0;
wire v$_18371_out1;
wire v$_18599_out0;
wire v$_18599_out1;
wire v$_18600_out0;
wire v$_18600_out1;
wire v$_18623_out0;
wire v$_18624_out0;
wire v$_18787_out0;
wire v$_18788_out0;
wire v$_18789_out0;
wire v$_18790_out0;
wire v$_18791_out0;
wire v$_18792_out0;
wire v$_18901_out0;
wire v$_18902_out0;
wire v$_2014_out0;
wire v$_2015_out0;
wire v$_2016_out0;
wire v$_2017_out0;
wire v$_2018_out0;
wire v$_2019_out0;
wire v$_2130_out0;
wire v$_2131_out0;
wire v$_2640_out0;
wire v$_2641_out0;
wire v$_2849_out0;
wire v$_2850_out0;
wire v$_3129_out0;
wire v$_3130_out0;
wire v$_3131_out0;
wire v$_3132_out0;
wire v$_3133_out0;
wire v$_3134_out0;
wire v$_3193_out0;
wire v$_3194_out0;
wire v$_3322_out0;
wire v$_3322_out1;
wire v$_3323_out0;
wire v$_3323_out1;
wire v$_3332_out0;
wire v$_3332_out1;
wire v$_3333_out0;
wire v$_3333_out1;
wire v$_346_out0;
wire v$_346_out1;
wire v$_347_out0;
wire v$_347_out1;
wire v$_3685_out0;
wire v$_3685_out1;
wire v$_3686_out0;
wire v$_3686_out1;
wire v$_3864_out0;
wire v$_3864_out1;
wire v$_3865_out0;
wire v$_3865_out1;
wire v$_3969_out0;
wire v$_3969_out1;
wire v$_3970_out0;
wire v$_3970_out1;
wire v$_4148_out0;
wire v$_4148_out1;
wire v$_4149_out0;
wire v$_4149_out1;
wire v$_4172_out0;
wire v$_4172_out1;
wire v$_4173_out0;
wire v$_4173_out1;
wire v$_4176_out0;
wire v$_4176_out1;
wire v$_4177_out0;
wire v$_4177_out1;
wire v$_42_out0;
wire v$_43_out0;
wire v$_4987_out0;
wire v$_4987_out1;
wire v$_4988_out0;
wire v$_4988_out1;
wire v$_5108_out0;
wire v$_5108_out1;
wire v$_5109_out0;
wire v$_5109_out1;
wire v$_5112_out1;
wire v$_5113_out1;
wire v$_5255_out0;
wire v$_5255_out1;
wire v$_5256_out0;
wire v$_5256_out1;
wire v$_5293_out0;
wire v$_5293_out1;
wire v$_5294_out0;
wire v$_5294_out1;
wire v$_5646_out0;
wire v$_5646_out1;
wire v$_5647_out0;
wire v$_5647_out1;
wire v$_6074_out0;
wire v$_6074_out1;
wire v$_6075_out0;
wire v$_6075_out1;
wire v$_6228_out0;
wire v$_6228_out1;
wire v$_6229_out0;
wire v$_6229_out1;
wire v$_6230_out0;
wire v$_6230_out1;
wire v$_6231_out0;
wire v$_6231_out1;
wire v$_6232_out0;
wire v$_6232_out1;
wire v$_6233_out0;
wire v$_6233_out1;
wire v$_6352_out0;
wire v$_6353_out0;
wire v$_7176_out0;
wire v$_7176_out1;
wire v$_7177_out0;
wire v$_7177_out1;
wire v$_7178_out0;
wire v$_7178_out1;
wire v$_7179_out0;
wire v$_7179_out1;
wire v$_7180_out0;
wire v$_7180_out1;
wire v$_7181_out0;
wire v$_7181_out1;
wire v$_7258_out0;
wire v$_7258_out1;
wire v$_7259_out0;
wire v$_7259_out1;
wire v$_7260_out0;
wire v$_7260_out1;
wire v$_7261_out0;
wire v$_7261_out1;
wire v$_7262_out0;
wire v$_7262_out1;
wire v$_7263_out0;
wire v$_7263_out1;
wire v$_7264_out0;
wire v$_7264_out1;
wire v$_7265_out0;
wire v$_7265_out1;
wire v$_7355_out0;
wire v$_7356_out0;
wire v$_7357_out0;
wire v$_7358_out0;
wire v$_7359_out0;
wire v$_7360_out0;
wire v$_7560_out0;
wire v$_7560_out1;
wire v$_7561_out0;
wire v$_7561_out1;
wire v$_7605_out0;
wire v$_7605_out1;
wire v$_7606_out0;
wire v$_7606_out1;
wire v$_7607_out0;
wire v$_7608_out0;
wire v$_7676_out0;
wire v$_7676_out1;
wire v$_7677_out0;
wire v$_7677_out1;
wire v$_7678_out0;
wire v$_7678_out1;
wire v$_7679_out0;
wire v$_7679_out1;
wire v$_7680_out0;
wire v$_7680_out1;
wire v$_7681_out0;
wire v$_7681_out1;
wire v$_7710_out0;
wire v$_7710_out1;
wire v$_7711_out0;
wire v$_7711_out1;
wire v$_7794_out0;
wire v$_7795_out0;
wire v$_7985_out0;
wire v$_7985_out1;
wire v$_7986_out0;
wire v$_7986_out1;
wire v$_7987_out0;
wire v$_7987_out1;
wire v$_7988_out0;
wire v$_7988_out1;
wire v$_7989_out0;
wire v$_7989_out1;
wire v$_7990_out0;
wire v$_7990_out1;
wire v$_7991_out0;
wire v$_7991_out1;
wire v$_7992_out0;
wire v$_7992_out1;
wire v$_7993_out0;
wire v$_7993_out1;
wire v$_7994_out0;
wire v$_7994_out1;
wire v$_7995_out0;
wire v$_7995_out1;
wire v$_7996_out0;
wire v$_7996_out1;
wire v$_8088_out0;
wire v$_8089_out0;
wire v$_8090_out0;
wire v$_8091_out0;
wire v$_8092_out0;
wire v$_8093_out0;
wire v$_8297_out0;
wire v$_8297_out1;
wire v$_8298_out0;
wire v$_8298_out1;
wire v$_8404_out0;
wire v$_8404_out1;
wire v$_8405_out0;
wire v$_8405_out1;
wire v$_8541_out0;
wire v$_8542_out0;
wire v$_9123_out0;
wire v$_9124_out0;
wire v$_9125_out0;
wire v$_9125_out1;
wire v$_9126_out0;
wire v$_9126_out1;
wire v$_9157_out0;
wire v$_9157_out1;
wire v$_9158_out0;
wire v$_9158_out1;
wire v$_9389_out0;
wire v$_9390_out0;
wire v$_9391_out0;
wire v$_9392_out0;
wire v$_9393_out0;
wire v$_9394_out0;
wire v$_9398_out0;
wire v$_9398_out1;
wire v$_9399_out0;
wire v$_9399_out1;
wire v$_9437_out0;
wire v$_9437_out1;
wire v$_9438_out0;
wire v$_9438_out1;
wire v$_9743_out0;
wire v$_9743_out1;
wire v$_9744_out0;
wire v$_9744_out1;
wire v$_9753_out0;
wire v$_9753_out1;
wire v$_9754_out0;
wire v$_9754_out1;
wire v$_9755_out0;
wire v$_9755_out1;
wire v$_9756_out0;
wire v$_9756_out1;
wire v$_9757_out0;
wire v$_9757_out1;
wire v$_9758_out0;
wire v$_9758_out1;
wire v$_9857_out0;
wire v$_9857_out1;
wire v$_9858_out0;
wire v$_9858_out1;
wire v$_9873_out0;
wire v$_9873_out1;
wire v$_9874_out0;
wire v$_9874_out1;
wire v$_9875_out0;
wire v$_9875_out1;
wire v$_9876_out0;
wire v$_9876_out1;
wire v$_9877_out0;
wire v$_9877_out1;
wire v$_9878_out0;
wire v$_9878_out1;
wire v$_9960_out0;
wire v$_9961_out0;
wire v$_996_out0;
wire v$_997_out0;
wire v$increment_18454_out0;
wire v$increment_18455_out0;

always @(posedge clk) v$FF1_2_out0 <= v$NEWINTERRUPT_7309_out0;
always @(posedge clk) v$FF1_3_out0 <= v$NEWINTERRUPT_7310_out0;
always @(posedge clk) v$FF1_194_out0 <= v$G3_8354_out0;
always @(posedge clk) v$FF1_195_out0 <= v$G3_8355_out0;
always @(posedge clk) v$INT2_265_out0 <= v$I2EN_16345_out0 ? v$SEL1_12547_out0 : v$INT2_265_out0;
always @(posedge clk) v$INT2_266_out0 <= v$I2EN_16346_out0 ? v$SEL1_12548_out0 : v$INT2_266_out0;
always @(posedge clk) v$FF3_271_out0 <= v$ShiftEN_8039_out0 ? v$MUX3_18332_out0 : v$FF3_271_out0;
always @(posedge clk) v$FF3_272_out0 <= v$ShiftEN_8040_out0 ? v$MUX3_18333_out0 : v$FF3_272_out0;
always @(posedge clk) v$INT3_281_out0 <= v$I3EN_18387_out0 ? v$SEL1_12547_out0 : v$INT3_281_out0;
always @(posedge clk) v$INT3_282_out0 <= v$I3EN_18388_out0 ? v$SEL1_12548_out0 : v$INT3_282_out0;
always @(posedge clk) v$REG13_308_out0 <= v$HALT0_380_out0;
always @(posedge clk) v$FF0_716_out0 <= v$CLK4_12779_out0 ? v$G1_15877_out0 : v$FF0_716_out0;
always @(posedge clk) v$FF0_717_out0 <= v$CLK4_12780_out0 ? v$G1_15878_out0 : v$FF0_717_out0;
always @(posedge clk) v$REG2_718_out0 <= v$increment_18454_out0 ? v$A2_15432_out0 : v$REG2_718_out0;
always @(posedge clk) v$REG2_719_out0 <= v$increment_18455_out0 ? v$A2_15433_out0 : v$REG2_719_out0;
always @(posedge clk) v$REG1_1309_out0 <= v$G14_16418_out0 ? v$A_11554_out0 : v$REG1_1309_out0;
always @(posedge clk) v$REG1_1310_out0 <= v$G14_16419_out0 ? v$A_11555_out0 : v$REG1_1310_out0;
always @(posedge clk) v$FF1_1325_out0 <= v$CLK4_12779_out0 ? v$G21_18276_out0 : v$FF1_1325_out0;
always @(posedge clk) v$FF1_1326_out0 <= v$CLK4_12780_out0 ? v$G21_18277_out0 : v$FF1_1326_out0;
always @(posedge clk) v$FF2_1327_out0 <= v$LDMAIN_14395_out0;
always @(posedge clk) v$FF2_1328_out0 <= v$LDMAIN_14396_out0;
always @(posedge clk) v$FF3_1456_out0 <= v$Shift_9986_out0 ? v$FF1_16797_out0 : v$FF3_1456_out0;
always @(posedge clk) v$FF3_1457_out0 <= v$Shift_9987_out0 ? v$FF1_16798_out0 : v$FF3_1457_out0;
always @(posedge clk) v$FF1_1539_out0 <= v$NEWINTERRUPT_4598_out0;
always @(posedge clk) v$FF1_1540_out0 <= v$NEWINTERRUPT_4599_out0;
always @(posedge clk) v$FF2_1729_out0 <= v$Shift_9986_out0 ? v$FF7_15152_out0 : v$FF2_1729_out0;
always @(posedge clk) v$FF2_1730_out0 <= v$Shift_9987_out0 ? v$FF7_15153_out0 : v$FF2_1730_out0;
always @(posedge clk) v$FF5_1915_out0 <= v$SHIFTEN_9781_out0 ? v$MUX1_2776_out0 : v$FF5_1915_out0;
always @(posedge clk) v$FF5_1916_out0 <= v$SHIFTEN_9782_out0 ? v$MUX1_2777_out0 : v$FF5_1916_out0;
always @(posedge clk) v$FF5_1917_out0 <= v$SHIFTEN_9783_out0 ? v$MUX1_2778_out0 : v$FF5_1917_out0;
always @(posedge clk) v$FF5_1918_out0 <= v$SHIFTEN_9784_out0 ? v$MUX1_2779_out0 : v$FF5_1918_out0;
always @(posedge clk) v$FF5_1919_out0 <= v$SHIFTEN_9785_out0 ? v$MUX1_2780_out0 : v$FF5_1919_out0;
always @(posedge clk) v$FF5_1920_out0 <= v$SHIFTEN_9786_out0 ? v$MUX1_2781_out0 : v$FF5_1920_out0;
always @(posedge clk) v$FF5_1921_out0 <= v$SHIFTEN_9787_out0 ? v$MUX1_2782_out0 : v$FF5_1921_out0;
always @(posedge clk) v$FF5_1922_out0 <= v$SHIFTEN_9788_out0 ? v$MUX1_2783_out0 : v$FF5_1922_out0;
always @(posedge clk) v$FF5_1923_out0 <= v$SHIFTEN_9789_out0 ? v$MUX1_2784_out0 : v$FF5_1923_out0;
always @(posedge clk) v$FF5_1924_out0 <= v$SHIFTEN_9790_out0 ? v$MUX1_2785_out0 : v$FF5_1924_out0;
always @(posedge clk) v$FF5_1925_out0 <= v$SHIFTEN_9791_out0 ? v$MUX1_2786_out0 : v$FF5_1925_out0;
always @(posedge clk) v$FF5_1926_out0 <= v$SHIFTEN_9792_out0 ? v$MUX1_2787_out0 : v$FF5_1926_out0;
always @(posedge clk) v$FF4_2541_out0 <= v$ShiftEN_8039_out0 ? v$MUX4_16228_out0 : v$FF4_2541_out0;
always @(posedge clk) v$FF4_2542_out0 <= v$ShiftEN_8040_out0 ? v$MUX4_16229_out0 : v$FF4_2542_out0;
always @(posedge clk) v$FF11_2642_out0 <= v$G50_16979_out0;
always @(posedge clk) v$FF11_2643_out0 <= v$G50_16980_out0;
always @(posedge clk) v$FF1_2722_out0 <= v$G4_15287_out0;
always @(posedge clk) v$FF1_2723_out0 <= v$G4_15288_out0;
always @(posedge clk) v$FF6_2817_out0 <= v$SHIFTEN_9781_out0 ? v$MUX3_10374_out0 : v$FF6_2817_out0;
always @(posedge clk) v$FF6_2818_out0 <= v$SHIFTEN_9782_out0 ? v$MUX3_10375_out0 : v$FF6_2818_out0;
always @(posedge clk) v$FF6_2819_out0 <= v$SHIFTEN_9783_out0 ? v$MUX3_10376_out0 : v$FF6_2819_out0;
always @(posedge clk) v$FF6_2820_out0 <= v$SHIFTEN_9784_out0 ? v$MUX3_10377_out0 : v$FF6_2820_out0;
always @(posedge clk) v$FF6_2821_out0 <= v$SHIFTEN_9785_out0 ? v$MUX3_10378_out0 : v$FF6_2821_out0;
always @(posedge clk) v$FF6_2822_out0 <= v$SHIFTEN_9786_out0 ? v$MUX3_10379_out0 : v$FF6_2822_out0;
always @(posedge clk) v$FF6_2823_out0 <= v$SHIFTEN_9787_out0 ? v$MUX3_10380_out0 : v$FF6_2823_out0;
always @(posedge clk) v$FF6_2824_out0 <= v$SHIFTEN_9788_out0 ? v$MUX3_10381_out0 : v$FF6_2824_out0;
always @(posedge clk) v$FF6_2825_out0 <= v$SHIFTEN_9789_out0 ? v$MUX3_10382_out0 : v$FF6_2825_out0;
always @(posedge clk) v$FF6_2826_out0 <= v$SHIFTEN_9790_out0 ? v$MUX3_10383_out0 : v$FF6_2826_out0;
always @(posedge clk) v$FF6_2827_out0 <= v$SHIFTEN_9791_out0 ? v$MUX3_10384_out0 : v$FF6_2827_out0;
always @(posedge clk) v$FF6_2828_out0 <= v$SHIFTEN_9792_out0 ? v$MUX3_10385_out0 : v$FF6_2828_out0;
always @(posedge clk) v$REG3_3046_out0 <= v$G55_18799_out0 ? v$MUX5_12517_out0 : v$REG3_3046_out0;
always @(posedge clk) v$REG3_3047_out0 <= v$G55_18800_out0 ? v$MUX5_12518_out0 : v$REG3_3047_out0;
always @(posedge clk) v$FF2_3160_out0 <= v$ShiftEN_8039_out0 ? v$MUX2_13871_out0 : v$FF2_3160_out0;
always @(posedge clk) v$FF2_3161_out0 <= v$ShiftEN_8040_out0 ? v$MUX2_13872_out0 : v$FF2_3161_out0;
v$ROM1_3190 I3190 (v$ROM1_3190_out0, v$_2810_out0, clk);
always @(posedge clk) v$REG12_3553_out0 <= v$HALT1_4317_out0 ? v$RAMADDR1_13239_out0 : v$REG12_3553_out0;
always @(posedge clk) v$FF3_3598_out0 <= v$G53_18133_out0;
always @(posedge clk) v$FF4_3963_out0 <= v$CAPTURE_251_out0 ? v$G6_12692_out0 : v$FF4_3963_out0;
always @(posedge clk) v$FF4_3964_out0 <= v$CAPTURE_252_out0 ? v$G6_12693_out0 : v$FF4_3964_out0;
always @(posedge clk) v$REG1_4200_out0 <= v$EN_16500_out0 ? v$MODE_11296_out0 : v$REG1_4200_out0;
always @(posedge clk) v$REG1_4201_out0 <= v$EN_16501_out0 ? v$MODE_11297_out0 : v$REG1_4201_out0;
always @(posedge clk) v$REG2_4204_out0 <= v$START_5733_out0 ? v$_2012_out0 : v$REG2_4204_out0;
always @(posedge clk) v$REG2_4205_out0 <= v$START_5734_out0 ? v$_2013_out0 : v$REG2_4205_out0;
always @(posedge clk) v$REG8_4264_out0 <= v$SELIN_18816_out0;
always @(posedge clk) v$FF0_4488_out0 <= v$CLK4_18601_out0 ? v$MUX1_7971_out0 : v$FF0_4488_out0;
always @(posedge clk) v$FF0_4489_out0 <= v$CLK4_18602_out0 ? v$MUX1_7972_out0 : v$FF0_4489_out0;
always @(posedge clk) v$FF1_4502_out0 <= v$START_5733_out0 ? v$IS$32$BITS_14649_out0 : v$FF1_4502_out0;
always @(posedge clk) v$FF1_4503_out0 <= v$START_5734_out0 ? v$IS$32$BITS_14650_out0 : v$FF1_4503_out0;
always @(posedge clk) v$FF2_4510_out0 <= v$CLK4_18601_out0 ? v$MUX3_6396_out0 : v$FF2_4510_out0;
always @(posedge clk) v$FF2_4511_out0 <= v$CLK4_18602_out0 ? v$MUX3_6397_out0 : v$FF2_4511_out0;
always @(posedge clk) v$FF5_4957_out0 <= v$EQ2_12176_out0;
always @(posedge clk) v$FF5_4958_out0 <= v$EQ2_12177_out0;
always @(posedge clk) v$REG1_5110_out0 <= v$D1_14709_out1 ? v$DIN3_15022_out0 : v$REG1_5110_out0;
always @(posedge clk) v$REG1_5111_out0 <= v$D1_14710_out1 ? v$DIN3_15023_out0 : v$REG1_5111_out0;
always @(posedge clk) v$FF0_5223_out0 <= v$G1_13725_out0;
always @(posedge clk) v$FF0_5224_out0 <= v$G1_13726_out0;
always @(posedge clk) v$REG2_5345_out0 <= v$HALT_16989_out0 ? v$G8_16329_out0 : v$REG2_5345_out0;
always @(posedge clk) v$FF1_5439_out0 <= v$NEXTSTATE_14110_out0;
always @(posedge clk) v$FF1_5440_out0 <= v$NEXTSTATE_14111_out0;
always @(posedge clk) v$FF1_5441_out0 <= v$NEXTSTATE_14112_out0;
always @(posedge clk) v$FF1_5442_out0 <= v$NEXTSTATE_14113_out0;
always @(posedge clk) v$FF1_5443_out0 <= v$NEXTSTATE_14114_out0;
always @(posedge clk) v$FF1_5444_out0 <= v$NEXTSTATE_14115_out0;
always @(posedge clk) v$FF1_5688_out0 <= v$G45_15949_out0;
always @(posedge clk) v$REG14_5698_out0 <= v$HALT1_4317_out0;
always @(posedge clk) v$FF1_6306_out0 <= v$INTERRUPT0_12268_out0;
always @(posedge clk) v$FF1_6307_out0 <= v$INTERRUPT0_12269_out0;
always @(posedge clk) v$FF1_6414_out0 <= v$CAPTURE_251_out0 ? v$I3_5036_out0 : v$FF1_6414_out0;
always @(posedge clk) v$FF1_6415_out0 <= v$CAPTURE_252_out0 ? v$I3_5037_out0 : v$FF1_6415_out0;
always @(posedge clk) v$REG7_6442_out0 <= v$G84_1386_out0;
always @(posedge clk) v$REG4_6885_out0 <= v$G66_9020_out0 ? v$MUX1_15845_out0 : v$REG4_6885_out0;
always @(posedge clk) v$REG4_6886_out0 <= v$G66_9021_out0 ? v$MUX1_15846_out0 : v$REG4_6886_out0;
always @(posedge clk) v$FF4_7301_out0 <= v$EQ1_14926_out0;
always @(posedge clk) v$FF4_7302_out0 <= v$EQ1_14927_out0;
always @(posedge clk) v$REG1_7363_out0 <= v$HALTVALID_8061_out0 ? v$NEXTSTATE_14116_out0 : v$REG1_7363_out0;
v$ROM1_7586 I7586 (v$ROM1_7586_out0, v$_2613_out0, clk);
always @(posedge clk) v$FF3_7649_out0 <= v$RX_44_out0;
always @(posedge clk) v$FF3_7650_out0 <= v$RX_45_out0;
always @(posedge clk) v$FF3_7887_out0 <= v$CAPTURE_251_out0 ? v$G9_16121_out0 : v$FF3_7887_out0;
always @(posedge clk) v$FF3_7888_out0 <= v$CAPTURE_252_out0 ? v$G9_16122_out0 : v$FF3_7888_out0;
always @(posedge clk) v$REG1_8170_out0 <= v$START_5733_out0 ? v$_13118_out0 : v$REG1_8170_out0;
always @(posedge clk) v$REG1_8171_out0 <= v$START_5734_out0 ? v$_13119_out0 : v$REG1_8171_out0;
always @(posedge clk) v$FF10_8216_out0 <= v$HALT_13471_out0;
always @(posedge clk) v$FF10_8217_out0 <= v$HALT_13472_out0;
always @(posedge clk) v$FF8_8346_out0 <= v$ShiftEN_8039_out0 ? v$MUX8_1651_out0 : v$FF8_8346_out0;
always @(posedge clk) v$FF8_8347_out0 <= v$ShiftEN_8040_out0 ? v$MUX8_1652_out0 : v$FF8_8347_out0;
always @(posedge clk) v$FF4_8369_out0 <= v$G68_15784_out0;
always @(posedge clk) v$FF4_8370_out0 <= v$G68_15785_out0;
always @(posedge clk) v$FF7_8401_out0 <= v$G62_12324_out0 ? v$R_9127_out0 : v$FF7_8401_out0;
always @(posedge clk) v$FF7_8402_out0 <= v$G62_12325_out0 ? v$R_9128_out0 : v$FF7_8402_out0;
always @(posedge clk) v$FF1_8531_out0 <= v$EXEC2_8362_out0 ? v$S_18561_out0 : v$FF1_8531_out0;
always @(posedge clk) v$FF1_8532_out0 <= v$EXEC2_8363_out0 ? v$S_18562_out0 : v$FF1_8532_out0;
always @(posedge clk) v$FF4_8562_out0 <= v$Shift_9986_out0 ? v$RX_3176_out0 : v$FF4_8562_out0;
always @(posedge clk) v$FF4_8563_out0 <= v$Shift_9987_out0 ? v$RX_3177_out0 : v$FF4_8563_out0;
always @(posedge clk) v$FF7_8609_out0 <= v$SHIFTEN_9781_out0 ? v$MUX8_3792_out0 : v$FF7_8609_out0;
always @(posedge clk) v$FF7_8610_out0 <= v$SHIFTEN_9782_out0 ? v$MUX8_3793_out0 : v$FF7_8610_out0;
always @(posedge clk) v$FF7_8611_out0 <= v$SHIFTEN_9783_out0 ? v$MUX8_3794_out0 : v$FF7_8611_out0;
always @(posedge clk) v$FF7_8612_out0 <= v$SHIFTEN_9784_out0 ? v$MUX8_3795_out0 : v$FF7_8612_out0;
always @(posedge clk) v$FF7_8613_out0 <= v$SHIFTEN_9785_out0 ? v$MUX8_3796_out0 : v$FF7_8613_out0;
always @(posedge clk) v$FF7_8614_out0 <= v$SHIFTEN_9786_out0 ? v$MUX8_3797_out0 : v$FF7_8614_out0;
always @(posedge clk) v$FF7_8615_out0 <= v$SHIFTEN_9787_out0 ? v$MUX8_3798_out0 : v$FF7_8615_out0;
always @(posedge clk) v$FF7_8616_out0 <= v$SHIFTEN_9788_out0 ? v$MUX8_3799_out0 : v$FF7_8616_out0;
always @(posedge clk) v$FF7_8617_out0 <= v$SHIFTEN_9789_out0 ? v$MUX8_3800_out0 : v$FF7_8617_out0;
always @(posedge clk) v$FF7_8618_out0 <= v$SHIFTEN_9790_out0 ? v$MUX8_3801_out0 : v$FF7_8618_out0;
always @(posedge clk) v$FF7_8619_out0 <= v$SHIFTEN_9791_out0 ? v$MUX8_3802_out0 : v$FF7_8619_out0;
always @(posedge clk) v$FF7_8620_out0 <= v$SHIFTEN_9792_out0 ? v$MUX8_3803_out0 : v$FF7_8620_out0;
always @(posedge clk) v$REG1_9169_out0 <= v$G6_3703_out0;
always @(posedge clk) v$REG1_9225_out0 <= v$EXEC2_9813_out0 ? v$MUX5_15088_out0 : v$REG1_9225_out0;
always @(posedge clk) v$REG1_9226_out0 <= v$EXEC2_9814_out0 ? v$MUX5_15089_out0 : v$REG1_9226_out0;
always @(posedge clk) v$FF6_9289_out0 <= v$Shift_9986_out0 ? v$FF8_17348_out0 : v$FF6_9289_out0;
always @(posedge clk) v$FF6_9290_out0 <= v$Shift_9987_out0 ? v$FF8_17349_out0 : v$FF6_9290_out0;
always @(posedge clk) v$FF0_9775_out0 <= v$G12_2420_out0;
always @(posedge clk) v$FF0_9776_out0 <= v$G12_2421_out0;
always @(posedge clk) v$FF2_9793_out0 <= v$STATUSREAD_1795_out0;
always @(posedge clk) v$FF2_9794_out0 <= v$STATUSREAD_1796_out0;
always @(posedge clk) v$FF1_9797_out0 <= v$ShiftEN_8039_out0 ? v$MUX1_435_out0 : v$FF1_9797_out0;
always @(posedge clk) v$FF1_9798_out0 <= v$ShiftEN_8040_out0 ? v$MUX1_436_out0 : v$FF1_9798_out0;
always @(posedge clk) v$FF1_9988_out0 <= v$CLK4_18601_out0 ? v$MUX2_6922_out0 : v$FF1_9988_out0;
always @(posedge clk) v$FF1_9989_out0 <= v$CLK4_18602_out0 ? v$MUX2_6923_out0 : v$FF1_9989_out0;
always @(posedge clk) v$REG11_10004_out0 <= v$HALT1_4317_out0 ? v$DATAIN1_10016_out0 : v$REG11_10004_out0;
always @(posedge clk) v$FF1_10012_out0 <= v$G2_5471_out0;
always @(posedge clk) v$FF1_10013_out0 <= v$G2_5472_out0;
always @(posedge clk) v$FF3_10396_out0 <= v$SHIFTEN_9781_out0 ? v$MUX5_9902_out0 : v$FF3_10396_out0;
always @(posedge clk) v$FF3_10397_out0 <= v$SHIFTEN_9782_out0 ? v$MUX5_9903_out0 : v$FF3_10397_out0;
always @(posedge clk) v$FF3_10398_out0 <= v$SHIFTEN_9783_out0 ? v$MUX5_9904_out0 : v$FF3_10398_out0;
always @(posedge clk) v$FF3_10399_out0 <= v$SHIFTEN_9784_out0 ? v$MUX5_9905_out0 : v$FF3_10399_out0;
always @(posedge clk) v$FF3_10400_out0 <= v$SHIFTEN_9785_out0 ? v$MUX5_9906_out0 : v$FF3_10400_out0;
always @(posedge clk) v$FF3_10401_out0 <= v$SHIFTEN_9786_out0 ? v$MUX5_9907_out0 : v$FF3_10401_out0;
always @(posedge clk) v$FF3_10402_out0 <= v$SHIFTEN_9787_out0 ? v$MUX5_9908_out0 : v$FF3_10402_out0;
always @(posedge clk) v$FF3_10403_out0 <= v$SHIFTEN_9788_out0 ? v$MUX5_9909_out0 : v$FF3_10403_out0;
always @(posedge clk) v$FF3_10404_out0 <= v$SHIFTEN_9789_out0 ? v$MUX5_9910_out0 : v$FF3_10404_out0;
always @(posedge clk) v$FF3_10405_out0 <= v$SHIFTEN_9790_out0 ? v$MUX5_9911_out0 : v$FF3_10405_out0;
always @(posedge clk) v$FF3_10406_out0 <= v$SHIFTEN_9791_out0 ? v$MUX5_9912_out0 : v$FF3_10406_out0;
always @(posedge clk) v$FF3_10407_out0 <= v$SHIFTEN_9792_out0 ? v$MUX5_9913_out0 : v$FF3_10407_out0;
always @(posedge clk) v$REG1_10757_out0 <= v$EXEC2_8362_out0 ? v$MUX6_14288_out0 : v$REG1_10757_out0;
always @(posedge clk) v$REG1_10758_out0 <= v$EXEC2_8363_out0 ? v$MUX6_14289_out0 : v$REG1_10758_out0;
always @(posedge clk) v$FF1_10761_out0 <= v$G5_7910_out0 ? v$A1_9805_out1 : v$FF1_10761_out0;
always @(posedge clk) v$FF1_10762_out0 <= v$G5_7911_out0 ? v$A1_9806_out1 : v$FF1_10762_out0;
always @(posedge clk) v$FF8_10797_out0 <= v$EQ3_4362_out0;
always @(posedge clk) v$FF8_10798_out0 <= v$EQ3_4363_out0;
always @(posedge clk) v$FF9_11158_out0 <= v$STP$DECODED_17154_out0;
always @(posedge clk) v$FF9_11159_out0 <= v$STP$DECODED_17155_out0;
always @(posedge clk) v$REG4_11270_out0 <= v$START_3879_out0 ? v$RD_12364_out0 : v$REG4_11270_out0;
always @(posedge clk) v$REG4_11271_out0 <= v$START_3880_out0 ? v$RD_12365_out0 : v$REG4_11271_out0;
always @(posedge clk) v$S$FF_11312_out0 <= v$EXEC2_1313_out0 ? v$S_11196_out0 : v$S$FF_11312_out0;
always @(posedge clk) v$S$FF_11313_out0 <= v$EXEC2_1314_out0 ? v$S_11197_out0 : v$S$FF_11313_out0;
always @(posedge clk) v$REG1_11407_out0 <= v$EXEC2_1621_out0 ? v$MUX5_8281_out0 : v$REG1_11407_out0;
always @(posedge clk) v$REG1_11408_out0 <= v$EXEC2_1622_out0 ? v$MUX5_8282_out0 : v$REG1_11408_out0;
always @(posedge clk) v$FF14_11409_out0 <= v$VALID_3893_out0;
always @(posedge clk) v$FF14_11410_out0 <= v$VALID_3894_out0;
always @(posedge clk) v$FF3_11419_out0 <= v$CLK4_18601_out0 ? v$MUX4_17682_out0 : v$FF3_11419_out0;
always @(posedge clk) v$FF3_11420_out0 <= v$CLK4_18602_out0 ? v$MUX4_17683_out0 : v$FF3_11420_out0;
always @(posedge clk) v$REG4_11502_out0 <= v$G88_7716_out0;
always @(posedge clk) v$REG3_11509_out0 <= v$D1_14709_out3 ? v$DIN3_15022_out0 : v$REG3_11509_out0;
always @(posedge clk) v$REG3_11510_out0 <= v$D1_14710_out3 ? v$DIN3_15023_out0 : v$REG3_11510_out0;
always @(posedge clk) v$FF1_11566_out0 <= v$G1_4372_out0;
always @(posedge clk) v$FF1_11567_out0 <= v$G1_4373_out0;
always @(posedge clk) v$REG3_12336_out0 <= v$G33_338_out0 ? v$SEL4_9936_out0 : v$REG3_12336_out0;
always @(posedge clk) v$REG3_12337_out0 <= v$G33_339_out0 ? v$SEL4_9937_out0 : v$REG3_12337_out0;
always @(posedge clk) v$REG2_12370_out0 <= v$IR2$VALID_13833_out0 ? v$_9123_out0 : v$REG2_12370_out0;
always @(posedge clk) v$REG2_12371_out0 <= v$IR2$VALID_13834_out0 ? v$_9124_out0 : v$REG2_12371_out0;
always @(posedge clk) v$REG1_12653_out0 <= v$OUT_15545_out0;
always @(posedge clk) v$REG1_12654_out0 <= v$OUT_15576_out0;
always @(posedge clk) v$FF15_13286_out0 <= v$HALT$PREV$PREV_18681_out0;
always @(posedge clk) v$FF15_13287_out0 <= v$HALT$PREV$PREV_18682_out0;
always @(posedge clk) v$FF7_13325_out0 <= v$STALL_18502_out0;
always @(posedge clk) v$FF7_13326_out0 <= v$STALL_18503_out0;
always @(posedge clk) v$PCNORMAL_13337_out0 <= v$G33_11239_out0 ? v$SUM_14246_out0 : v$PCNORMAL_13337_out0;
always @(posedge clk) v$PCNORMAL_13338_out0 <= v$G33_11240_out0 ? v$SUM_14247_out0 : v$PCNORMAL_13338_out0;
v$RAM1_13483 I13483 (v$RAM1_13483_out0, v$RAMADDR_14184_out0, v$MUX2_16447_out0, v$RAMWEN_18576_out0, clk);
always @(posedge clk) v$FF2_13615_out0 <= v$G7_14734_out0;
always @(posedge clk) v$FF2_13616_out0 <= v$G7_14735_out0;
always @(posedge clk) v$FF2_13617_out0 <= v$G7_14736_out0;
always @(posedge clk) v$FF2_13618_out0 <= v$G7_14737_out0;
always @(posedge clk) v$FF2_13619_out0 <= v$G7_14738_out0;
always @(posedge clk) v$FF2_13620_out0 <= v$G7_14739_out0;
always @(posedge clk) v$FF2_13621_out0 <= v$G4_12405_out0;
always @(posedge clk) v$FF2_13622_out0 <= v$G4_12406_out0;
always @(posedge clk) v$FF2_13623_out0 <= v$G4_12407_out0;
always @(posedge clk) v$FF2_13624_out0 <= v$G4_12408_out0;
always @(posedge clk) v$FF2_13625_out0 <= v$G4_12409_out0;
always @(posedge clk) v$FF2_13626_out0 <= v$G7_14740_out0;
always @(posedge clk) v$FF2_13627_out0 <= v$G7_14741_out0;
always @(posedge clk) v$FF2_13628_out0 <= v$G7_14742_out0;
always @(posedge clk) v$FF2_13629_out0 <= v$G7_14743_out0;
always @(posedge clk) v$FF2_13630_out0 <= v$G7_14744_out0;
always @(posedge clk) v$FF2_13631_out0 <= v$G7_14745_out0;
always @(posedge clk) v$FF2_13632_out0 <= v$G4_12410_out0;
always @(posedge clk) v$FF2_13633_out0 <= v$G4_12411_out0;
always @(posedge clk) v$FF2_13634_out0 <= v$G4_12412_out0;
always @(posedge clk) v$FF2_13635_out0 <= v$G4_12413_out0;
always @(posedge clk) v$FF2_13636_out0 <= v$G4_12414_out0;
always @(posedge clk) v$FF1_13671_out0 <= v$G16_6632_out0 ? v$G7_1991_out0 : v$FF1_13671_out0;
always @(posedge clk) v$FF1_13672_out0 <= v$G16_6633_out0 ? v$G7_1992_out0 : v$FF1_13672_out0;
always @(posedge clk) v$FF2_14043_out0 <= v$G51_19373_out0;
always @(posedge clk) v$FF4_14125_out0 <= v$G54_13869_out0;
always @(posedge clk) v$REG1_14166_out0 <= v$MUX1_18934_out0;
always @(posedge clk) v$REG1_14167_out0 <= v$MUX1_18935_out0;
always @(posedge clk) v$FF1_14261_out0 <= v$EXEC2_9813_out0 ? v$S_10809_out0 : v$FF1_14261_out0;
always @(posedge clk) v$FF1_14262_out0 <= v$EXEC2_9814_out0 ? v$S_10810_out0 : v$FF1_14262_out0;
always @(posedge clk) v$REG1_14701_out0 <= v$G1_12789_out0 ? v$MUX1_5354_out0 : v$REG1_14701_out0;
always @(posedge clk) v$REG1_14702_out0 <= v$G1_12790_out0 ? v$MUX1_5355_out0 : v$REG1_14702_out0;
always @(posedge clk) v$REG1_14711_out0 <= v$IR1$VALID_62_out0 ? v$RM_18797_out0 : v$REG1_14711_out0;
always @(posedge clk) v$REG1_14712_out0 <= v$IR1$VALID_63_out0 ? v$RM_18798_out0 : v$REG1_14712_out0;
always @(posedge clk) v$FF10_14804_out0 <= v$WREN_11505_out0;
always @(posedge clk) v$FF10_14805_out0 <= v$WREN_11506_out0;
always @(posedge clk) v$FF8_15064_out0 <= v$SHIFTEN_9781_out0 ? v$MUX4_17458_out0 : v$FF8_15064_out0;
always @(posedge clk) v$FF8_15065_out0 <= v$SHIFTEN_9782_out0 ? v$MUX4_17459_out0 : v$FF8_15065_out0;
always @(posedge clk) v$FF8_15066_out0 <= v$SHIFTEN_9783_out0 ? v$MUX4_17460_out0 : v$FF8_15066_out0;
always @(posedge clk) v$FF8_15067_out0 <= v$SHIFTEN_9784_out0 ? v$MUX4_17461_out0 : v$FF8_15067_out0;
always @(posedge clk) v$FF8_15068_out0 <= v$SHIFTEN_9785_out0 ? v$MUX4_17462_out0 : v$FF8_15068_out0;
always @(posedge clk) v$FF8_15069_out0 <= v$SHIFTEN_9786_out0 ? v$MUX4_17463_out0 : v$FF8_15069_out0;
always @(posedge clk) v$FF8_15070_out0 <= v$SHIFTEN_9787_out0 ? v$MUX4_17464_out0 : v$FF8_15070_out0;
always @(posedge clk) v$FF8_15071_out0 <= v$SHIFTEN_9788_out0 ? v$MUX4_17465_out0 : v$FF8_15071_out0;
always @(posedge clk) v$FF8_15072_out0 <= v$SHIFTEN_9789_out0 ? v$MUX4_17466_out0 : v$FF8_15072_out0;
always @(posedge clk) v$FF8_15073_out0 <= v$SHIFTEN_9790_out0 ? v$MUX4_17467_out0 : v$FF8_15073_out0;
always @(posedge clk) v$FF8_15074_out0 <= v$SHIFTEN_9791_out0 ? v$MUX4_17468_out0 : v$FF8_15074_out0;
always @(posedge clk) v$FF8_15075_out0 <= v$SHIFTEN_9792_out0 ? v$MUX4_17469_out0 : v$FF8_15075_out0;
always @(posedge clk) v$FF7_15152_out0 <= v$Shift_9986_out0 ? v$FF6_9289_out0 : v$FF7_15152_out0;
always @(posedge clk) v$FF7_15153_out0 <= v$Shift_9987_out0 ? v$FF6_9290_out0 : v$FF7_15153_out0;
always @(posedge clk) v$FF2_15233_out0 <= v$CLK4_12779_out0 ? v$G24_10000_out0 : v$FF2_15233_out0;
always @(posedge clk) v$FF2_15234_out0 <= v$CLK4_12780_out0 ? v$G24_10001_out0 : v$FF2_15234_out0;
always @(posedge clk) v$FF2_15390_out0 <= v$SHIFTEN_9781_out0 ? v$MUX6_10839_out0 : v$FF2_15390_out0;
always @(posedge clk) v$FF2_15391_out0 <= v$SHIFTEN_9782_out0 ? v$MUX6_10840_out0 : v$FF2_15391_out0;
always @(posedge clk) v$FF2_15392_out0 <= v$SHIFTEN_9783_out0 ? v$MUX6_10841_out0 : v$FF2_15392_out0;
always @(posedge clk) v$FF2_15393_out0 <= v$SHIFTEN_9784_out0 ? v$MUX6_10842_out0 : v$FF2_15393_out0;
always @(posedge clk) v$FF2_15394_out0 <= v$SHIFTEN_9785_out0 ? v$MUX6_10843_out0 : v$FF2_15394_out0;
always @(posedge clk) v$FF2_15395_out0 <= v$SHIFTEN_9786_out0 ? v$MUX6_10844_out0 : v$FF2_15395_out0;
always @(posedge clk) v$FF2_15396_out0 <= v$SHIFTEN_9787_out0 ? v$MUX6_10845_out0 : v$FF2_15396_out0;
always @(posedge clk) v$FF2_15397_out0 <= v$SHIFTEN_9788_out0 ? v$MUX6_10846_out0 : v$FF2_15397_out0;
always @(posedge clk) v$FF2_15398_out0 <= v$SHIFTEN_9789_out0 ? v$MUX6_10847_out0 : v$FF2_15398_out0;
always @(posedge clk) v$FF2_15399_out0 <= v$SHIFTEN_9790_out0 ? v$MUX6_10848_out0 : v$FF2_15399_out0;
always @(posedge clk) v$FF2_15400_out0 <= v$SHIFTEN_9791_out0 ? v$MUX6_10849_out0 : v$FF2_15400_out0;
always @(posedge clk) v$FF2_15401_out0 <= v$SHIFTEN_9792_out0 ? v$MUX6_10850_out0 : v$FF2_15401_out0;
always @(posedge clk) v$REG1_15444_out0 <= v$MUX1_10337_out0;
always @(posedge clk) v$REG1_15445_out0 <= v$MUX1_10338_out0;
always @(posedge clk) v$REG2_15622_out0 <= v$R_18958_out0;
always @(posedge clk) v$REG2_15623_out0 <= v$R_18959_out0;
always @(posedge clk) v$FF3_15648_out0 <= v$INTERRUPT2_1821_out0;
always @(posedge clk) v$FF3_15649_out0 <= v$INTERRUPT2_1822_out0;
always @(posedge clk) v$FF6_15909_out0 <= v$ShiftEN_8039_out0 ? v$MUX6_9458_out0 : v$FF6_15909_out0;
always @(posedge clk) v$FF6_15910_out0 <= v$ShiftEN_8040_out0 ? v$MUX6_9459_out0 : v$FF6_15910_out0;
always @(posedge clk) v$FF2_16070_out0 <= v$G1_5662_out0;
always @(posedge clk) v$FF2_16071_out0 <= v$G1_5663_out0;
always @(posedge clk) v$REG2_16210_out0 <= v$G13_8221_out0 ? v$B_3590_out0 : v$REG2_16210_out0;
always @(posedge clk) v$REG2_16211_out0 <= v$G13_8222_out0 ? v$B_3591_out0 : v$REG2_16211_out0;
always @(posedge clk) v$INT0_16488_out0 <= v$I0EN_8356_out0 ? v$SEL1_12547_out0 : v$INT0_16488_out0;
always @(posedge clk) v$INT0_16489_out0 <= v$I0EN_8357_out0 ? v$SEL1_12548_out0 : v$INT0_16489_out0;
always @(posedge clk) v$FF3_16564_out0 <= v$CLK4_12779_out0 ? v$G32_16952_out0 : v$FF3_16564_out0;
always @(posedge clk) v$FF3_16565_out0 <= v$CLK4_12780_out0 ? v$G32_16953_out0 : v$FF3_16565_out0;
always @(posedge clk) v$FF4_16584_out0 <= v$SHIFTEN_9781_out0 ? v$MUX2_14407_out0 : v$FF4_16584_out0;
always @(posedge clk) v$FF4_16585_out0 <= v$SHIFTEN_9782_out0 ? v$MUX2_14408_out0 : v$FF4_16585_out0;
always @(posedge clk) v$FF4_16586_out0 <= v$SHIFTEN_9783_out0 ? v$MUX2_14409_out0 : v$FF4_16586_out0;
always @(posedge clk) v$FF4_16587_out0 <= v$SHIFTEN_9784_out0 ? v$MUX2_14410_out0 : v$FF4_16587_out0;
always @(posedge clk) v$FF4_16588_out0 <= v$SHIFTEN_9785_out0 ? v$MUX2_14411_out0 : v$FF4_16588_out0;
always @(posedge clk) v$FF4_16589_out0 <= v$SHIFTEN_9786_out0 ? v$MUX2_14412_out0 : v$FF4_16589_out0;
always @(posedge clk) v$FF4_16590_out0 <= v$SHIFTEN_9787_out0 ? v$MUX2_14413_out0 : v$FF4_16590_out0;
always @(posedge clk) v$FF4_16591_out0 <= v$SHIFTEN_9788_out0 ? v$MUX2_14414_out0 : v$FF4_16591_out0;
always @(posedge clk) v$FF4_16592_out0 <= v$SHIFTEN_9789_out0 ? v$MUX2_14415_out0 : v$FF4_16592_out0;
always @(posedge clk) v$FF4_16593_out0 <= v$SHIFTEN_9790_out0 ? v$MUX2_14416_out0 : v$FF4_16593_out0;
always @(posedge clk) v$FF4_16594_out0 <= v$SHIFTEN_9791_out0 ? v$MUX2_14417_out0 : v$FF4_16594_out0;
always @(posedge clk) v$FF4_16595_out0 <= v$SHIFTEN_9792_out0 ? v$MUX2_14418_out0 : v$FF4_16595_out0;
always @(posedge clk) v$FF9_16635_out0 <= v$FF10_14804_out0 ? v$G26_16633_out0 : v$FF9_16635_out0;
always @(posedge clk) v$FF9_16636_out0 <= v$FF10_14805_out0 ? v$G26_16634_out0 : v$FF9_16636_out0;
always @(posedge clk) v$FF1_16687_out0 <= v$SHIFTEN_9781_out0 ? v$MUX7_18517_out0 : v$FF1_16687_out0;
always @(posedge clk) v$FF1_16688_out0 <= v$SHIFTEN_9782_out0 ? v$MUX7_18518_out0 : v$FF1_16688_out0;
always @(posedge clk) v$FF1_16689_out0 <= v$SHIFTEN_9783_out0 ? v$MUX7_18519_out0 : v$FF1_16689_out0;
always @(posedge clk) v$FF1_16690_out0 <= v$SHIFTEN_9784_out0 ? v$MUX7_18520_out0 : v$FF1_16690_out0;
always @(posedge clk) v$FF1_16691_out0 <= v$SHIFTEN_9785_out0 ? v$MUX7_18521_out0 : v$FF1_16691_out0;
always @(posedge clk) v$FF1_16692_out0 <= v$SHIFTEN_9786_out0 ? v$MUX7_18522_out0 : v$FF1_16692_out0;
always @(posedge clk) v$FF1_16693_out0 <= v$SHIFTEN_9787_out0 ? v$MUX7_18523_out0 : v$FF1_16693_out0;
always @(posedge clk) v$FF1_16694_out0 <= v$SHIFTEN_9788_out0 ? v$MUX7_18524_out0 : v$FF1_16694_out0;
always @(posedge clk) v$FF1_16695_out0 <= v$SHIFTEN_9789_out0 ? v$MUX7_18525_out0 : v$FF1_16695_out0;
always @(posedge clk) v$FF1_16696_out0 <= v$SHIFTEN_9790_out0 ? v$MUX7_18526_out0 : v$FF1_16696_out0;
always @(posedge clk) v$FF1_16697_out0 <= v$SHIFTEN_9791_out0 ? v$MUX7_18527_out0 : v$FF1_16697_out0;
always @(posedge clk) v$FF1_16698_out0 <= v$SHIFTEN_9792_out0 ? v$MUX7_18528_out0 : v$FF1_16698_out0;
always @(posedge clk) v$REG9_16701_out0 <= v$HALT0_380_out0 ? v$RAMADDR0_17579_out0 : v$REG9_16701_out0;
always @(posedge clk) v$FF6_16780_out0 <= v$PHALT1_9264_out0;
always @(posedge clk) v$FF1_16797_out0 <= v$Shift_9986_out0 ? v$FF2_1729_out0 : v$FF1_16797_out0;
always @(posedge clk) v$FF1_16798_out0 <= v$Shift_9987_out0 ? v$FF2_1730_out0 : v$FF1_16798_out0;
always @(posedge clk) v$REG0_16864_out0 <= v$D1_14709_out0 ? v$DIN3_15022_out0 : v$REG0_16864_out0;
always @(posedge clk) v$REG0_16865_out0 <= v$D1_14710_out0 ? v$DIN3_15023_out0 : v$REG0_16865_out0;
always @(posedge clk) v$FF1_16930_out0 <= v$EXEC2_1621_out0 ? v$S_10894_out0 : v$FF1_16930_out0;
always @(posedge clk) v$FF1_16931_out0 <= v$EXEC2_1622_out0 ? v$S_10895_out0 : v$FF1_16931_out0;
always @(posedge clk) v$FF2_16954_out0 <= v$CAPTURE_251_out0 ? v$G1_14123_out0 : v$FF2_16954_out0;
always @(posedge clk) v$FF2_16955_out0 <= v$CAPTURE_252_out0 ? v$G1_14124_out0 : v$FF2_16955_out0;
always @(posedge clk) v$FF5_16956_out0 <= v$ShiftEN_8039_out0 ? v$MUX5_19171_out0 : v$FF5_16956_out0;
always @(posedge clk) v$FF5_16957_out0 <= v$ShiftEN_8040_out0 ? v$MUX5_19172_out0 : v$FF5_16957_out0;
always @(posedge clk) v$REG2_16962_out0 <= v$THRESHOLD$WRITE_7550_out0 ? v$THRESHOLD_16123_out0 : v$REG2_16962_out0;
always @(posedge clk) v$REG2_16963_out0 <= v$THRESHOLD$WRITE_7551_out0 ? v$THRESHOLD_16124_out0 : v$REG2_16963_out0;
always @(posedge clk) v$FF5_17047_out0 <= v$PHALT0_12199_out0;
always @(posedge clk) v$FF12_17048_out0 <= v$FF10_8216_out0;
always @(posedge clk) v$FF12_17049_out0 <= v$FF10_8217_out0;
always @(posedge clk) v$REG10_17089_out0 <= v$HALT0_380_out0 ? v$DATAIN0_11570_out0 : v$REG10_17089_out0;
always @(posedge clk) v$FF2_17272_out0 <= v$INTERRUPT1_18306_out0;
always @(posedge clk) v$FF2_17273_out0 <= v$INTERRUPT1_18307_out0;
always @(posedge clk) v$FF8_17348_out0 <= v$Shift_9986_out0 ? v$FF4_8562_out0 : v$FF8_17348_out0;
always @(posedge clk) v$FF8_17349_out0 <= v$Shift_9987_out0 ? v$FF4_8563_out0 : v$FF8_17349_out0;
always @(posedge clk) v$REG2_17420_out0 <= v$_7693_out0;
always @(posedge clk) v$REG2_17421_out0 <= v$_7694_out0;
always @(posedge clk) v$REG2_18120_out0 <= v$D1_14709_out2 ? v$DIN3_15022_out0 : v$REG2_18120_out0;
always @(posedge clk) v$REG2_18121_out0 <= v$D1_14710_out2 ? v$DIN3_15023_out0 : v$REG2_18121_out0;
always @(posedge clk) v$REG3_18364_out0 <= v$IR2$VALID_13833_out0 ? v$EQ1_16882_out0 : v$REG3_18364_out0;
always @(posedge clk) v$REG3_18365_out0 <= v$IR2$VALID_13834_out0 ? v$EQ1_16883_out0 : v$REG3_18365_out0;
always @(posedge clk) v$PCINTERRUPT_18413_out0 <= v$ININTERRUPT_1277_out0 ? v$SUM_14246_out0 : v$PCINTERRUPT_18413_out0;
always @(posedge clk) v$PCINTERRUPT_18414_out0 <= v$ININTERRUPT_1278_out0 ? v$SUM_14247_out0 : v$PCINTERRUPT_18414_out0;
always @(posedge clk) v$FF4_18456_out0 <= v$C1_5674_out0;
always @(posedge clk) v$FF4_18457_out0 <= v$C1_5675_out0;
always @(posedge clk) v$FF3_18727_out0 <= v$G29_8174_out0;
always @(posedge clk) v$FF3_18728_out0 <= v$G29_8175_out0;
always @(posedge clk) v$FF7_18731_out0 <= v$ShiftEN_8039_out0 ? v$MUX7_9855_out0 : v$FF7_18731_out0;
always @(posedge clk) v$FF7_18732_out0 <= v$ShiftEN_8040_out0 ? v$MUX7_9856_out0 : v$FF7_18732_out0;
always @(posedge clk) v$FF4_19047_out0 <= v$INTERRUPT3_3040_out0;
always @(posedge clk) v$FF4_19048_out0 <= v$INTERRUPT3_3041_out0;
always @(posedge clk) v$FF5_19083_out0 <= v$Shift_9986_out0 ? v$FF3_1456_out0 : v$FF5_19083_out0;
always @(posedge clk) v$FF5_19084_out0 <= v$Shift_9987_out0 ? v$FF3_1457_out0 : v$FF5_19084_out0;
always @(posedge clk) v$LSB$FF_19125_out0 <= v$EXEC2_1313_out0 ? v$MUX5_17662_out0 : v$LSB$FF_19125_out0;
always @(posedge clk) v$LSB$FF_19126_out0 <= v$EXEC2_1314_out0 ? v$MUX5_17663_out0 : v$LSB$FF_19126_out0;
always @(posedge clk) v$INT1_19145_out0 <= v$I1EN_19009_out0 ? v$SEL1_12547_out0 : v$INT1_19145_out0;
always @(posedge clk) v$INT1_19146_out0 <= v$I1EN_19010_out0 ? v$SEL1_12548_out0 : v$INT1_19146_out0;
always @(posedge clk) v$FF13_19153_out0 <= v$FF7_13325_out0;
always @(posedge clk) v$FF13_19154_out0 <= v$FF7_13326_out0;
always @(posedge clk) v$REG1_19272_out0 <= v$MODEWRITE_15321_out0 ? v$SEL1_18848_out0 : v$REG1_19272_out0;
always @(posedge clk) v$REG1_19273_out0 <= v$MODEWRITE_15322_out0 ? v$SEL1_18849_out0 : v$REG1_19273_out0;
assign v$C9_19372_out0 = 16'h0;
assign v$C9_19371_out0 = 16'h0;
assign v$C3_19164_out0 = 1'h0;
assign v$C3_19163_out0 = 1'h0;
assign v$C3_19046_out0 = 24'h0;
assign v$C3_19045_out0 = 24'h0;
assign v$C2_18927_out0 = 1'h0;
assign v$C2_18926_out0 = 1'h0;
assign v$CIN_18833_out0 = 1'h1;
assign v$CIN_18832_out0 = 1'h1;
assign v$CIN_18831_out0 = 1'h1;
assign v$CIN_18830_out0 = 1'h1;
assign v$CIN_18829_out0 = 1'h1;
assign v$CIN_18828_out0 = 1'h1;
assign v$CIN_18827_out0 = 1'h1;
assign v$CIN_18826_out0 = 1'h1;
assign v$C1_18810_out0 = 16'h0;
assign v$C1_18809_out0 = 16'h0;
assign v$C3_18740_out0 = 1'h0;
assign v$C3_18739_out0 = 1'h0;
assign v$C2_18618_out0 = 15'h0;
assign v$C2_18617_out0 = 15'h0;
assign v$C4_18590_out0 = 24'h0;
assign v$C4_18589_out0 = 24'h0;
assign v$C1_18275_out0 = 1'h0;
assign v$C1_18274_out0 = 1'h0;
assign v$C1_18273_out0 = 1'h0;
assign v$C1_18272_out0 = 1'h0;
assign v$C1_18271_out0 = 1'h0;
assign v$C1_18270_out0 = 1'h0;
assign v$C1_18269_out0 = 1'h0;
assign v$C1_18268_out0 = 1'h0;
assign v$C1_18267_out0 = 1'h0;
assign v$C1_18266_out0 = 1'h0;
assign v$C1_17982_out0 = 1'h1;
assign v$C1_17981_out0 = 1'h1;
assign v$C1_17980_out0 = 1'h1;
assign v$C1_17979_out0 = 1'h1;
assign v$C2_17615_out0 = 1'h0;
assign v$C2_17614_out0 = 1'h0;
assign v$C5_17526_out0 = 2'h2;
assign v$C5_17525_out0 = 1'h0;
assign v$C5_17524_out0 = 2'h2;
assign v$C5_17523_out0 = 1'h0;
assign v$C5_17522_out0 = 2'h2;
assign v$C5_17521_out0 = 1'h0;
assign v$C5_17520_out0 = 2'h2;
assign v$C5_17519_out0 = 1'h0;
assign v$C1_17455_out0 = 3'h0;
assign v$C1_17454_out0 = 3'h0;
assign v$C4_17137_out0 = 2'h1;
assign v$C4_17136_out0 = 2'h1;
assign v$C4_17135_out0 = 2'h1;
assign v$C4_17134_out0 = 2'h1;
assign v$CON4_17062_out0 = 1'h0;
assign v$CON4_17061_out0 = 1'h0;
assign v$CON4_17060_out0 = 1'h0;
assign v$CON4_17059_out0 = 1'h0;
assign v$CON4_17058_out0 = 1'h0;
assign v$CON4_17057_out0 = 1'h0;
assign v$C2_16949_out0 = 1'h1;
assign v$C2_16948_out0 = 1'h1;
assign v$C2_16947_out0 = 1'h1;
assign v$C2_16946_out0 = 1'h1;
assign v$C1_16939_out0 = 16'h0;
assign v$C1_16938_out0 = 16'h0;
assign v$C4_16917_out0 = 2'h0;
assign v$C4_16916_out0 = 2'h0;
assign v$C2_16897_out0 = 1'h0;
assign v$C2_16896_out0 = 1'h0;
assign v$C2_16895_out0 = 1'h0;
assign v$C2_16894_out0 = 1'h0;
assign v$C2_16852_out0 = 1'h1;
assign v$C2_16851_out0 = 1'h1;
assign v$C1_16844_out0 = 24'h0;
assign v$C1_16843_out0 = 24'h0;
assign v$C5_16706_out0 = 1'h0;
assign v$C5_16705_out0 = 1'h0;
assign v$C2_16597_out0 = 6'h1;
assign v$C2_16596_out0 = 6'h1;
assign v$C1_16547_out0 = 12'h0;
assign v$C1_16546_out0 = 12'h0;
assign v$C1_16527_out0 = 1'h1;
assign v$C1_16526_out0 = 1'h1;
assign v$C4_16510_out0 = 12'h0;
assign v$C4_16509_out0 = 12'h0;
assign v$C1_16408_out0 = 11'h0;
assign v$C1_16407_out0 = 11'h0;
assign v$C1_16333_out0 = 5'h1f;
assign v$C1_16332_out0 = 5'h1f;
assign v$C1_16320_out0 = 1'h0;
assign v$C1_16319_out0 = 1'h0;
assign v$C1_16318_out0 = 1'h0;
assign v$C1_16317_out0 = 1'h0;
assign v$C1_16273_out0 = 5'h0;
assign v$C1_16272_out0 = 5'h0;
assign v$C5_16213_out0 = 23'h0;
assign v$C5_16212_out0 = 23'h0;
assign v$C9_15848_out0 = 24'hffffff;
assign v$C9_15847_out0 = 24'hffffff;
assign v$C1_15810_out0 = 32'h0;
assign v$C1_15809_out0 = 32'h0;
assign v$C2_15781_out0 = 1'h0;
assign v$C2_15780_out0 = 1'h0;
assign v$C2_15779_out0 = 1'h0;
assign v$C2_15778_out0 = 1'h0;
assign v$C4_15443_out0 = 1'h1;
assign v$C4_15442_out0 = 1'h1;
assign v$C4_15441_out0 = 1'h1;
assign v$C4_15440_out0 = 1'h1;
assign v$C1_15420_out0 = 8'h0;
assign v$C1_15419_out0 = 8'h0;
assign v$C4_15260_out0 = 5'h0;
assign v$C4_15259_out0 = 5'h0;
assign v$C7_15248_out0 = 24'h0;
assign v$C7_15247_out0 = 24'h0;
assign v$CON2_14976_out0 = 1'h0;
assign v$CON2_14975_out0 = 1'h0;
assign v$CON2_14974_out0 = 1'h0;
assign v$CON2_14973_out0 = 1'h0;
assign v$CON2_14972_out0 = 1'h0;
assign v$CON2_14971_out0 = 1'h0;
assign v$C1_14856_out0 = 2'h3;
assign v$C1_14855_out0 = 2'h3;
assign v$C1_14640_out0 = 1'h0;
assign v$C1_14639_out0 = 1'h0;
assign v$C4_14637_out0 = 32'h0;
assign v$C4_14636_out0 = 32'h0;
assign v$C1_14600_out0 = 8'h0;
assign v$C1_14599_out0 = 8'h0;
assign v$C8_14200_out0 = 24'hffffff;
assign v$C8_14199_out0 = 24'hffffff;
assign v$C1_14155_out0 = 8'hff;
assign v$C1_14154_out0 = 5'h1f;
assign v$C1_14153_out0 = 8'hff;
assign v$C1_14152_out0 = 5'h1f;
assign v$C1_14151_out0 = 8'hff;
assign v$C1_14150_out0 = 5'h1f;
assign v$C1_14149_out0 = 8'hff;
assign v$C1_14148_out0 = 5'h1f;
assign v$C10_14118_out0 = 3'h0;
assign v$C10_14117_out0 = 3'h0;
assign v$C3_14093_out0 = 1'h1;
assign v$C3_14092_out0 = 1'h1;
assign v$C3_14091_out0 = 1'h1;
assign v$C3_14090_out0 = 1'h1;
assign v$C2_14083_out0 = 1'h0;
assign v$C2_14082_out0 = 1'h0;
assign v$C1_14034_out0 = 8'h0;
assign v$C1_14033_out0 = 8'h0;
assign v$C2_13972_out0 = 2'h1;
assign v$C2_13971_out0 = 2'h1;
assign v$C2_13911_out0 = 3'h0;
assign v$C2_13910_out0 = 3'h0;
assign v$C3_13742_out0 = 6'h0;
assign v$C3_13741_out0 = 6'h0;
assign v$CON6_13576_out0 = 1'h0;
assign v$CON6_13575_out0 = 1'h0;
assign v$CON6_13574_out0 = 1'h0;
assign v$CON6_13573_out0 = 1'h0;
assign v$CON6_13572_out0 = 1'h0;
assign v$CON6_13571_out0 = 1'h0;
assign v$C1_13424_out0 = 1'h0;
assign v$C1_13423_out0 = 1'h0;
assign v$C1_13396_out0 = 4'h0;
assign v$C1_13395_out0 = 4'h0;
assign v$C6_13146_out0 = 1'h1;
assign v$C6_13145_out0 = 1'h1;
assign v$C2_12773_out0 = 16'hffff;
assign v$C2_12772_out0 = 16'hffff;
assign v$C3_12771_out0 = 16'h0;
assign v$C3_12770_out0 = 16'h0;
assign v$C2_11199_out0 = 1'h1;
assign v$C2_11198_out0 = 1'h1;
assign v$CON5_11181_out0 = 1'h0;
assign v$CON5_11180_out0 = 1'h0;
assign v$CON5_11179_out0 = 1'h0;
assign v$CON5_11178_out0 = 1'h0;
assign v$CON5_11177_out0 = 1'h0;
assign v$CON5_11176_out0 = 1'h0;
assign v$C2_10435_out0 = 16'hffff;
assign v$C2_10434_out0 = 16'hffff;
assign v$C7_9872_out0 = 1'h1;
assign v$C7_9871_out0 = 1'h1;
assign v$C10_9280_out0 = 13'h0;
assign v$C10_9279_out0 = 13'h0;
assign v$C6_9183_out0 = 1'h0;
assign v$C6_9182_out0 = 1'h0;
assign v$C5_9115_out0 = 1'h1;
assign v$C5_9114_out0 = 1'h1;
assign v$C5_9113_out0 = 1'h1;
assign v$C5_9112_out0 = 1'h1;
assign v$C4_8569_out0 = 31'h0;
assign v$C4_8568_out0 = 15'h0;
assign v$C4_8567_out0 = 31'h0;
assign v$C4_8566_out0 = 15'h0;
assign v$C8_8516_out0 = 13'h0;
assign v$C8_8515_out0 = 13'h0;
assign v$C6_8361_out0 = 6'h1;
assign v$C6_8360_out0 = 6'h1;
assign v$C1_8294_out0 = 8'h0;
assign v$C1_8293_out0 = 4'h0;
assign v$C1_8292_out0 = 2'h0;
assign v$C1_8291_out0 = 1'h0;
assign v$C1_8290_out0 = 8'h0;
assign v$C1_8289_out0 = 4'h0;
assign v$C1_8288_out0 = 2'h0;
assign v$C1_8287_out0 = 1'h0;
assign v$CON3_8244_out0 = 1'h0;
assign v$CON3_8243_out0 = 1'h0;
assign v$CON3_8242_out0 = 1'h0;
assign v$CON3_8241_out0 = 1'h0;
assign v$CON3_8240_out0 = 1'h0;
assign v$CON3_8239_out0 = 1'h0;
assign v$C1_8042_out0 = 2'h2;
assign v$C1_8041_out0 = 2'h2;
assign v$C2_7960_out0 = 1'h1;
assign v$C2_7959_out0 = 1'h1;
assign v$C2_7958_out0 = 1'h1;
assign v$C2_7957_out0 = 1'h1;
assign v$C2_7956_out0 = 1'h1;
assign v$C2_7955_out0 = 1'h1;
assign v$C2_7954_out0 = 1'h1;
assign v$C2_7953_out0 = 1'h1;
assign v$C2_7952_out0 = 1'h1;
assign v$C2_7951_out0 = 1'h1;
assign v$C1_7743_out0 = 5'h0;
assign v$C1_7742_out0 = 5'h0;
assign v$C8_7600_out0 = 4'h0;
assign v$C8_7599_out0 = 4'h0;
assign v$C3_7298_out0 = 5'h17;
assign v$C3_7297_out0 = 5'h17;
assign v$C4_6860_out0 = 3'h0;
assign v$C4_6859_out0 = 3'h0;
assign v$C6_6778_out0 = 2'h3;
assign v$C6_6777_out0 = 2'h2;
assign v$C6_6776_out0 = 2'h3;
assign v$C6_6775_out0 = 2'h2;
assign v$C6_6774_out0 = 2'h3;
assign v$C6_6773_out0 = 2'h2;
assign v$C6_6772_out0 = 2'h3;
assign v$C6_6771_out0 = 2'h2;
assign v$C1_6704_out0 = 1'h0;
assign v$C1_6703_out0 = 1'h0;
assign v$C10_6625_out0 = 16'h0;
assign v$C10_6624_out0 = 16'h0;
assign v$C4_6607_out0 = 1'h0;
assign v$C4_6606_out0 = 1'h0;
assign v$C7_6319_out0 = 13'h0;
assign v$C7_6318_out0 = 13'h0;
assign v$C1_6303_out0 = 1'h0;
assign v$C1_6302_out0 = 2'h0;
assign v$C1_6301_out0 = 16'h0;
assign v$C1_6300_out0 = 4'h0;
assign v$C1_6299_out0 = 8'h0;
assign v$C1_6298_out0 = 1'h0;
assign v$C1_6297_out0 = 2'h0;
assign v$C1_6296_out0 = 4'h0;
assign v$C1_6295_out0 = 1'h0;
assign v$C1_6294_out0 = 8'h0;
assign v$C1_6293_out0 = 16'h0;
assign v$C1_6292_out0 = 2'h0;
assign v$C1_6291_out0 = 16'h0;
assign v$C1_6290_out0 = 4'h0;
assign v$C1_6289_out0 = 8'h0;
assign v$C1_6288_out0 = 1'h0;
assign v$C1_6287_out0 = 2'h0;
assign v$C1_6286_out0 = 4'h0;
assign v$C1_6285_out0 = 1'h0;
assign v$C1_6284_out0 = 8'h0;
assign v$C1_6283_out0 = 16'h0;
assign v$C1_6282_out0 = 2'h0;
assign v$C1_6281_out0 = 4'h0;
assign v$C1_6280_out0 = 1'h0;
assign v$C1_6279_out0 = 8'h0;
assign v$C1_6278_out0 = 16'h0;
assign v$C1_6277_out0 = 2'h0;
assign v$C1_6276_out0 = 4'h0;
assign v$C1_6275_out0 = 1'h0;
assign v$C1_6274_out0 = 8'h0;
assign v$C1_6273_out0 = 16'h0;
assign v$C1_6272_out0 = 1'h0;
assign v$C1_6271_out0 = 2'h0;
assign v$C1_6270_out0 = 16'h0;
assign v$C1_6269_out0 = 4'h0;
assign v$C1_6268_out0 = 8'h0;
assign v$C1_6267_out0 = 1'h0;
assign v$C1_6266_out0 = 2'h0;
assign v$C1_6265_out0 = 4'h0;
assign v$C1_6264_out0 = 1'h0;
assign v$C1_6263_out0 = 8'h0;
assign v$C1_6262_out0 = 16'h0;
assign v$C1_6261_out0 = 2'h0;
assign v$C1_6260_out0 = 16'h0;
assign v$C1_6259_out0 = 4'h0;
assign v$C1_6258_out0 = 8'h0;
assign v$C1_6257_out0 = 1'h0;
assign v$C1_6256_out0 = 2'h0;
assign v$C1_6255_out0 = 4'h0;
assign v$C1_6254_out0 = 1'h0;
assign v$C1_6253_out0 = 8'h0;
assign v$C1_6252_out0 = 16'h0;
assign v$C1_6251_out0 = 2'h0;
assign v$C1_6250_out0 = 4'h0;
assign v$C1_6249_out0 = 1'h0;
assign v$C1_6248_out0 = 8'h0;
assign v$C1_6247_out0 = 16'h0;
assign v$C1_6246_out0 = 2'h0;
assign v$C1_6245_out0 = 4'h0;
assign v$C1_6244_out0 = 1'h0;
assign v$C1_6243_out0 = 8'h0;
assign v$C1_6242_out0 = 16'h0;
assign v$C1_6239_out0 = 8'h81;
assign v$C1_6238_out0 = 5'h11;
assign v$C1_6237_out0 = 8'h81;
assign v$C1_6236_out0 = 5'h11;
assign v$C1_5675_out0 = 1'h1;
assign v$C1_5674_out0 = 1'h1;
assign v$C1_5655_out0 = 4'h0;
assign v$C1_5654_out0 = 4'h0;
assign v$C3_5629_out0 = 1'h1;
assign v$C3_5628_out0 = 1'h1;
assign v$C1_5456_out0 = 5'h0;
assign v$C1_5455_out0 = 5'h0;
assign v$C1_4638_out0 = 1'h0;
assign v$C1_4637_out0 = 1'h0;
assign v$C1_4636_out0 = 1'h0;
assign v$C1_4635_out0 = 1'h0;
assign v$C1_4634_out0 = 1'h0;
assign v$C1_4633_out0 = 1'h0;
assign v$C1_4630_out0 = 24'h0;
assign v$C1_4629_out0 = 24'h0;
assign v$C1_4628_out0 = 24'h0;
assign v$C1_4627_out0 = 24'h0;
assign v$C1_4626_out0 = 24'h0;
assign v$C1_4625_out0 = 24'h0;
assign v$C1_4624_out0 = 24'h0;
assign v$C1_4623_out0 = 24'h0;
assign v$C1_4521_out0 = 1'h1;
assign v$C1_4520_out0 = 1'h1;
assign v$C5_4270_out0 = 32'h0;
assign v$C5_4269_out0 = 32'h0;
assign v$CON1_4241_out0 = 1'h0;
assign v$CON1_4240_out0 = 1'h0;
assign v$CON1_4239_out0 = 1'h0;
assign v$CON1_4238_out0 = 1'h0;
assign v$CON1_4237_out0 = 1'h0;
assign v$CON1_4236_out0 = 1'h0;
assign v$C4_3936_out0 = 1'h1;
assign v$C4_3935_out0 = 1'h1;
assign v$C11_3823_out0 = 1'h0;
assign v$C11_3822_out0 = 1'h0;
assign v$C2_3819_out0 = 1'h1;
assign v$C2_3818_out0 = 1'h1;
assign v$C3_3530_out0 = 2'h0;
assign v$C3_3529_out0 = 2'h0;
assign v$C3_3528_out0 = 2'h0;
assign v$C3_3527_out0 = 2'h0;
assign v$C9_3526_out0 = 16'h0;
assign v$C9_3525_out0 = 16'h0;
assign v$C1_3230_out0 = 2'h0;
assign v$C1_3229_out0 = 2'h0;
assign v$C2_3186_out0 = 1'h1;
assign v$C2_3185_out0 = 1'h1;
assign v$C4_3128_out0 = 1'h1;
assign v$C4_3127_out0 = 1'h1;
assign v$C2_2864_out0 = 1'h0;
assign v$C2_2863_out0 = 1'h0;
assign v$C1_2841_out0 = 1'h1;
assign v$C1_2840_out0 = 1'h1;
assign v$C1_2839_out0 = 1'h1;
assign v$C1_2838_out0 = 1'h1;
assign v$C1_2837_out0 = 1'h1;
assign v$C1_2836_out0 = 1'h1;
assign v$C1_2835_out0 = 1'h1;
assign v$C1_2834_out0 = 1'h1;
assign v$C1_2833_out0 = 1'h1;
assign v$C1_2832_out0 = 1'h1;
assign v$C1_2831_out0 = 1'h1;
assign v$C1_2830_out0 = 1'h1;
assign v$C4_2645_out0 = 13'h0;
assign v$C4_2644_out0 = 13'h0;
assign v$CON7_2619_out0 = 1'h0;
assign v$CON7_2618_out0 = 1'h0;
assign v$CON7_2617_out0 = 1'h0;
assign v$CON7_2616_out0 = 1'h0;
assign v$CON7_2615_out0 = 1'h0;
assign v$CON7_2614_out0 = 1'h0;
assign v$C7_1868_out0 = 16'h0;
assign v$C7_1867_out0 = 16'h0;
assign v$C6_1726_out0 = 1'h1;
assign v$C6_1725_out0 = 1'h1;
assign v$C1_1712_out0 = 8'hff;
assign v$C1_1711_out0 = 8'hff;
assign v$C6_1690_out0 = 13'h0;
assign v$C6_1689_out0 = 13'h0;
assign v$C1_1670_out0 = 1'h0;
assign v$C1_1669_out0 = 1'h0;
assign v$C1_1624_out0 = 1'h0;
assign v$C1_1623_out0 = 1'h0;
assign v$C2_1608_out0 = 1'h1;
assign v$C2_1607_out0 = 1'h1;
assign v$C3_1526_out0 = 1'h1;
assign v$C3_1525_out0 = 1'h1;
assign v$C2_1318_out0 = 1'h1;
assign v$C2_1317_out0 = 1'h1;
assign v$C7_355_out0 = 1'h0;
assign v$C7_354_out0 = 1'h0;
assign v$C2_165_out0 = 1'h0;
assign v$C2_164_out0 = 2'h0;
assign v$C2_163_out0 = 16'h0;
assign v$C2_162_out0 = 4'h0;
assign v$C2_161_out0 = 8'h0;
assign v$C2_160_out0 = 1'h0;
assign v$C2_159_out0 = 2'h0;
assign v$C2_158_out0 = 4'h0;
assign v$C2_157_out0 = 1'h0;
assign v$C2_156_out0 = 8'h0;
assign v$C2_155_out0 = 16'h0;
assign v$C2_154_out0 = 2'h0;
assign v$C2_153_out0 = 16'h0;
assign v$C2_152_out0 = 4'h0;
assign v$C2_151_out0 = 8'h0;
assign v$C2_150_out0 = 1'h0;
assign v$C2_149_out0 = 2'h0;
assign v$C2_148_out0 = 4'h0;
assign v$C2_147_out0 = 1'h0;
assign v$C2_146_out0 = 8'h0;
assign v$C2_145_out0 = 16'h0;
assign v$C2_144_out0 = 2'h0;
assign v$C2_143_out0 = 4'h0;
assign v$C2_142_out0 = 1'h0;
assign v$C2_141_out0 = 8'h0;
assign v$C2_140_out0 = 16'h0;
assign v$C2_139_out0 = 2'h0;
assign v$C2_138_out0 = 4'h0;
assign v$C2_137_out0 = 1'h0;
assign v$C2_136_out0 = 8'h0;
assign v$C2_135_out0 = 16'h0;
assign v$C2_134_out0 = 1'h0;
assign v$C2_133_out0 = 2'h0;
assign v$C2_132_out0 = 16'h0;
assign v$C2_131_out0 = 4'h0;
assign v$C2_130_out0 = 8'h0;
assign v$C2_129_out0 = 1'h0;
assign v$C2_128_out0 = 2'h0;
assign v$C2_127_out0 = 4'h0;
assign v$C2_126_out0 = 1'h0;
assign v$C2_125_out0 = 8'h0;
assign v$C2_124_out0 = 16'h0;
assign v$C2_123_out0 = 2'h0;
assign v$C2_122_out0 = 16'h0;
assign v$C2_121_out0 = 4'h0;
assign v$C2_120_out0 = 8'h0;
assign v$C2_119_out0 = 1'h0;
assign v$C2_118_out0 = 2'h0;
assign v$C2_117_out0 = 4'h0;
assign v$C2_116_out0 = 1'h0;
assign v$C2_115_out0 = 8'h0;
assign v$C2_114_out0 = 16'h0;
assign v$C2_113_out0 = 2'h0;
assign v$C2_112_out0 = 4'h0;
assign v$C2_111_out0 = 1'h0;
assign v$C2_110_out0 = 8'h0;
assign v$C2_109_out0 = 16'h0;
assign v$C2_108_out0 = 2'h0;
assign v$C2_107_out0 = 4'h0;
assign v$C2_106_out0 = 1'h0;
assign v$C2_105_out0 = 8'h0;
assign v$C2_104_out0 = 16'h0;
assign v$G3_20_out0 = !(v$FF0_5223_out0 || v$FF1_10012_out0);
assign v$G3_21_out0 = !(v$FF0_5224_out0 || v$FF1_10013_out0);
assign v$G2_66_out0 = ! v$FF1_194_out0;
assign v$G2_67_out0 = ! v$FF1_195_out0;
assign v$Q0_74_out0 = v$FF0_9775_out0;
assign v$Q0_75_out0 = v$FF0_9776_out0;
assign v$SIN_95_out0 = v$C7_354_out0;
assign v$SIN_101_out0 = v$C7_355_out0;
assign v$G58_168_out0 = ! v$FF5_4957_out0;
assign v$G58_169_out0 = ! v$FF5_4958_out0;
assign v$_1429_out0 = { v$FF0_9775_out0,v$FF1_2722_out0 };
assign v$_1430_out0 = { v$FF0_9776_out0,v$FF1_2723_out0 };
assign v$G2_1447_out0 = ((v$FF5_19083_out0 && !v$FF3_1456_out0) || (!v$FF5_19083_out0) && v$FF3_1456_out0);
assign v$G2_1448_out0 = ((v$FF5_19084_out0 && !v$FF3_1457_out0) || (!v$FF5_19084_out0) && v$FF3_1457_out0);
assign v$INITIAL$FETCH$OCCURRED_1691_out0 = v$FF4_18456_out0;
assign v$INITIAL$FETCH$OCCURRED_1692_out0 = v$FF4_18457_out0;
assign v$PHALT_1794_out0 = v$REG2_5345_out0;
assign v$SELOUT_1880_out0 = v$REG8_4264_out0;
assign v$SOUT1_2080_out0 = v$FF4_16584_out0;
assign v$SOUT1_2081_out0 = v$FF4_16585_out0;
assign v$SOUT1_2082_out0 = v$FF4_16586_out0;
assign v$SOUT1_2083_out0 = v$FF4_16587_out0;
assign v$SOUT1_2084_out0 = v$FF4_16588_out0;
assign v$SOUT1_2085_out0 = v$FF4_16589_out0;
assign v$SOUT1_2086_out0 = v$FF4_16590_out0;
assign v$SOUT1_2087_out0 = v$FF4_16591_out0;
assign v$SOUT1_2088_out0 = v$FF4_16592_out0;
assign v$SOUT1_2089_out0 = v$FF4_16593_out0;
assign v$SOUT1_2090_out0 = v$FF4_16594_out0;
assign v$SOUT1_2091_out0 = v$FF4_16595_out0;
assign v$I2P_2465_out0 = v$FF2_16954_out0;
assign v$I2P_2466_out0 = v$FF2_16955_out0;
assign v$_2471_out0 = { v$FF7_18731_out0,v$FF8_8346_out0 };
assign v$_2472_out0 = { v$FF7_18732_out0,v$FF8_8347_out0 };
assign v$PIPELINERESTART_2611_out0 = v$FF1_2_out0;
assign v$PIPELINERESTART_2612_out0 = v$FF1_3_out0;
assign v$G4_3096_out0 = ((v$FF7_15152_out0 && !v$FF6_9289_out0) || (!v$FF7_15152_out0) && v$FF6_9289_out0);
assign v$G4_3097_out0 = ((v$FF7_15153_out0 && !v$FF6_9290_out0) || (!v$FF7_15153_out0) && v$FF6_9290_out0);
assign v$LEFT$SHIT_3270_out0 = v$C1_17979_out0;
assign v$LEFT$SHIT_3271_out0 = v$C4_15440_out0;
assign v$LEFT$SHIT_3272_out0 = v$C3_14090_out0;
assign v$LEFT$SHIT_3273_out0 = v$C5_9112_out0;
assign v$LEFT$SHIT_3274_out0 = v$C2_16946_out0;
assign v$LEFT$SHIT_3280_out0 = v$C1_17980_out0;
assign v$LEFT$SHIT_3281_out0 = v$C4_15441_out0;
assign v$LEFT$SHIT_3282_out0 = v$C3_14091_out0;
assign v$LEFT$SHIT_3283_out0 = v$C5_9113_out0;
assign v$LEFT$SHIT_3284_out0 = v$C2_16947_out0;
assign v$LEFT$SHIT_3285_out0 = v$C1_14639_out0;
assign v$LEFT$SHIT_3301_out0 = v$C1_17981_out0;
assign v$LEFT$SHIT_3302_out0 = v$C4_15442_out0;
assign v$LEFT$SHIT_3303_out0 = v$C3_14092_out0;
assign v$LEFT$SHIT_3304_out0 = v$C5_9114_out0;
assign v$LEFT$SHIT_3305_out0 = v$C2_16948_out0;
assign v$LEFT$SHIT_3311_out0 = v$C1_17982_out0;
assign v$LEFT$SHIT_3312_out0 = v$C4_15443_out0;
assign v$LEFT$SHIT_3313_out0 = v$C3_14093_out0;
assign v$LEFT$SHIT_3314_out0 = v$C5_9115_out0;
assign v$LEFT$SHIT_3315_out0 = v$C2_16949_out0;
assign v$LEFT$SHIT_3316_out0 = v$C1_14640_out0;
assign v$Q2_3367_out0 = v$FF2_16070_out0;
assign v$Q2_3368_out0 = v$FF2_16071_out0;
assign v$R0_3503_out0 = v$REG0_16864_out0;
assign v$R0_3504_out0 = v$REG0_16865_out0;
assign v$S$REG_3653_out0 = v$REG1_11407_out0;
assign v$S$REG_3654_out0 = v$REG1_11408_out0;
assign v$A$SAVED_3877_out0 = v$REG1_1309_out0;
assign v$A$SAVED_3878_out0 = v$REG1_1310_out0;
assign v$_3967_out0 = { v$FF7_15152_out0,v$FF6_9289_out0 };
assign v$_3968_out0 = { v$FF7_15153_out0,v$FF6_9290_out0 };
assign v$EN_4056_out0 = v$C7_9871_out0;
assign v$EN_4059_out0 = v$C7_9872_out0;
assign {v$A1_4168_out1,v$A1_4168_out0 } = v$REG1_15444_out0 + v$C2_16596_out0 + v$C1_1669_out0;
assign {v$A1_4169_out1,v$A1_4169_out0 } = v$REG1_15445_out0 + v$C2_16597_out0 + v$C1_1670_out0;
assign v$Q1_4619_out0 = v$FF1_9988_out0;
assign v$Q1_4620_out0 = v$FF1_9989_out0;
assign v$B$SAVED_4961_out0 = v$REG2_16210_out0;
assign v$B$SAVED_4962_out0 = v$REG2_16211_out0;
assign v$_5112_out0 = v$REG1_19272_out0[2:0];
assign v$_5112_out1 = v$REG1_19272_out0[3:1];
assign v$_5113_out0 = v$REG1_19273_out0[2:0];
assign v$_5113_out1 = v$REG1_19273_out0[3:1];
assign v$RESULT_5279_out0 = v$REG2_17420_out0;
assign v$RESULT_5280_out0 = v$REG2_17421_out0;
assign v$Wordlength_5358_out0 = v$REG1_15444_out0 == 6'h27;
assign v$Wordlength_5359_out0 = v$REG1_15445_out0 == 6'h27;
assign v$G2_5471_out0 = ((v$FF0_5223_out0 && !v$FF1_10012_out0) || (!v$FF0_5223_out0) && v$FF1_10012_out0);
assign v$G2_5472_out0 = ((v$FF0_5224_out0 && !v$FF1_10013_out0) || (!v$FF0_5224_out0) && v$FF1_10013_out0);
assign v$OUT_5477_out0 = v$ROM1_7586_out0;
assign v$Q2_5696_out0 = v$FF2_15233_out0;
assign v$Q2_5697_out0 = v$FF2_15234_out0;
assign v$G17_5717_out0 = ! v$FF2_17272_out0;
assign v$G17_5718_out0 = ! v$FF2_17273_out0;
assign v$D_6009_out0 = v$REG1_14701_out0;
assign v$D_6010_out0 = v$REG1_14702_out0;
assign v$STALL$PREV$CYCLE_6059_out0 = v$FF7_13325_out0;
assign v$STALL$PREV$CYCLE_6060_out0 = v$FF7_13326_out0;
assign v$STALL$PREV$PREV_6096_out0 = v$FF13_19153_out0;
assign v$STALL$PREV$PREV_6097_out0 = v$FF13_19154_out0;
assign v$IR$READ$IN$PREV$CYCLE_6449_out0 = v$REG2_15622_out0;
assign v$IR$READ$IN$PREV$CYCLE_6450_out0 = v$REG2_15623_out0;
assign v$I1P_6684_out0 = v$FF3_7887_out0;
assign v$I1P_6685_out0 = v$FF3_7888_out0;
assign v$EQ1_7213_out0 = v$REG2_16962_out0 == 16'h0;
assign v$EQ1_7214_out0 = v$REG2_16963_out0 == 16'h0;
assign v$PHALT1$PREV_7682_out0 = v$FF6_16780_out0;
assign v$G20_7717_out0 = ((v$FF7_18731_out0 && !v$FF8_8346_out0) || (!v$FF7_18731_out0) && v$FF8_8346_out0);
assign v$G20_7718_out0 = ((v$FF7_18732_out0 && !v$FF8_8347_out0) || (!v$FF7_18732_out0) && v$FF8_8347_out0);
assign v$PHALT0$PREV_7940_out0 = v$FF5_17047_out0;
assign v$HALT$PREV$PREV$PREV_8049_out0 = v$FF15_13286_out0;
assign v$HALT$PREV$PREV$PREV_8050_out0 = v$FF15_13287_out0;
assign v$_8051_out0 = { v$FF3_271_out0,v$FF4_2541_out0 };
assign v$_8052_out0 = { v$FF3_272_out0,v$FF4_2542_out0 };
assign v$LSB_8138_out0 = v$LSB$FF_19125_out0;
assign v$LSB_8139_out0 = v$LSB$FF_19126_out0;
assign v$LSBS_8263_out0 = v$REG1_10757_out0;
assign v$LSBS_8264_out0 = v$REG1_10758_out0;
assign v$R2_8285_out0 = v$REG2_18120_out0;
assign v$R2_8286_out0 = v$REG2_18121_out0;
assign v$OUT_8651_out0 = v$ROM1_3190_out0;
assign v$B2_8720_out0 = v$C7_15247_out0;
assign v$B2_8723_out0 = v$C7_15248_out0;
assign v$CINA_8777_out0 = v$CON6_13571_out0;
assign v$CINA_8778_out0 = v$CON7_2614_out0;
assign v$CINA_8790_out0 = v$CON4_17057_out0;
assign v$CINA_8792_out0 = v$CON5_11176_out0;
assign v$CINA_8795_out0 = v$CON2_14971_out0;
assign v$CINA_8801_out0 = v$CON1_4236_out0;
assign v$CINA_8806_out0 = v$CON3_8239_out0;
assign v$CINA_8818_out0 = v$CON6_13572_out0;
assign v$CINA_8819_out0 = v$CON7_2615_out0;
assign v$CINA_8831_out0 = v$CON4_17058_out0;
assign v$CINA_8833_out0 = v$CON5_11177_out0;
assign v$CINA_8836_out0 = v$CON2_14972_out0;
assign v$CINA_8842_out0 = v$CON1_4237_out0;
assign v$CINA_8847_out0 = v$CON3_8240_out0;
assign v$CINA_8859_out0 = v$CON6_13573_out0;
assign v$CINA_8860_out0 = v$CON7_2616_out0;
assign v$CINA_8872_out0 = v$CON4_17059_out0;
assign v$CINA_8874_out0 = v$CON5_11178_out0;
assign v$CINA_8877_out0 = v$CON2_14973_out0;
assign v$CINA_8883_out0 = v$CON1_4238_out0;
assign v$CINA_8888_out0 = v$CON3_8241_out0;
assign v$CINA_8900_out0 = v$CON6_13574_out0;
assign v$CINA_8901_out0 = v$CON7_2617_out0;
assign v$CINA_8913_out0 = v$CON4_17060_out0;
assign v$CINA_8915_out0 = v$CON5_11179_out0;
assign v$CINA_8918_out0 = v$CON2_14974_out0;
assign v$CINA_8924_out0 = v$CON1_4239_out0;
assign v$CINA_8929_out0 = v$CON3_8242_out0;
assign v$CINA_8941_out0 = v$CON6_13575_out0;
assign v$CINA_8942_out0 = v$CON7_2618_out0;
assign v$CINA_8954_out0 = v$CON4_17061_out0;
assign v$CINA_8956_out0 = v$CON5_11180_out0;
assign v$CINA_8959_out0 = v$CON2_14975_out0;
assign v$CINA_8965_out0 = v$CON1_4240_out0;
assign v$CINA_8970_out0 = v$CON3_8243_out0;
assign v$CINA_8982_out0 = v$CON6_13576_out0;
assign v$CINA_8983_out0 = v$CON7_2619_out0;
assign v$CINA_8995_out0 = v$CON4_17062_out0;
assign v$CINA_8997_out0 = v$CON5_11181_out0;
assign v$CINA_9000_out0 = v$CON2_14976_out0;
assign v$CINA_9006_out0 = v$CON1_4241_out0;
assign v$CINA_9011_out0 = v$CON3_8244_out0;
assign v$PHALT1_9264_out0 = v$REG14_5698_out0;
assign v$I3P_9295_out0 = v$FF1_6414_out0;
assign v$I3P_9296_out0 = v$FF1_6415_out0;
assign v$G23_9729_out0 = ((v$FF1_9797_out0 && !v$FF2_3160_out0) || (!v$FF1_9797_out0) && v$FF2_3160_out0);
assign v$G23_9730_out0 = ((v$FF1_9798_out0 && !v$FF2_3161_out0) || (!v$FF1_9798_out0) && v$FF2_3161_out0);
assign v$SHIFTEN_9781_out0 = v$C1_2830_out0;
assign v$SHIFTEN_9782_out0 = v$C1_2831_out0;
assign v$SHIFTEN_9783_out0 = v$C1_2832_out0;
assign v$SHIFTEN_9784_out0 = v$C1_2833_out0;
assign v$SHIFTEN_9785_out0 = v$C1_2834_out0;
assign v$SHIFTEN_9786_out0 = v$C1_2835_out0;
assign v$SHIFTEN_9787_out0 = v$C1_2836_out0;
assign v$SHIFTEN_9788_out0 = v$C1_2837_out0;
assign v$SHIFTEN_9789_out0 = v$C1_2838_out0;
assign v$SHIFTEN_9790_out0 = v$C1_2839_out0;
assign v$SHIFTEN_9791_out0 = v$C1_2840_out0;
assign v$SHIFTEN_9792_out0 = v$C1_2841_out0;
assign v$_9811_out0 = { v$FF8_17348_out0,v$FF4_8562_out0 };
assign v$_9812_out0 = { v$FF8_17349_out0,v$FF4_8563_out0 };
assign v$RecievedParity_9916_out0 = v$FF7_8401_out0;
assign v$RecievedParity_9917_out0 = v$FF7_8402_out0;
assign v$G31_10014_out0 = ! v$FF4_19047_out0;
assign v$G31_10015_out0 = ! v$FF4_19048_out0;
assign v$G63_10444_out0 = ! v$FF8_10797_out0;
assign v$G63_10445_out0 = ! v$FF8_10798_out0;
assign v$I0P_10763_out0 = v$FF4_3963_out0;
assign v$I0P_10764_out0 = v$FF4_3964_out0;
assign v$OUTPUT_10799_out0 = v$FF1_5439_out0;
assign v$OUTPUT_10800_out0 = v$FF1_5440_out0;
assign v$OUTPUT_10801_out0 = v$FF1_5441_out0;
assign v$OUTPUT_10802_out0 = v$FF1_5442_out0;
assign v$OUTPUT_10803_out0 = v$FF1_5443_out0;
assign v$OUTPUT_10804_out0 = v$FF1_5444_out0;
assign v$HALT$PREV_10837_out0 = v$FF10_8216_out0;
assign v$HALT$PREV_10838_out0 = v$FF10_8217_out0;
assign v$R3_11234_out0 = v$REG3_11509_out0;
assign v$R3_11235_out0 = v$REG3_11510_out0;
assign v$Q1_11427_out0 = v$FF1_1325_out0;
assign v$Q1_11428_out0 = v$FF1_1326_out0;
assign v$PHALT0_12199_out0 = v$REG13_308_out0;
assign v$ISINTERRUPTED_12429_out0 = v$FF1_13671_out0;
assign v$ISINTERRUPTED_12430_out0 = v$FF1_13672_out0;
assign v$G21_12447_out0 = ((v$FF5_16956_out0 && !v$FF6_15909_out0) || (!v$FF5_16956_out0) && v$FF6_15909_out0);
assign v$G21_12448_out0 = ((v$FF5_16957_out0 && !v$FF6_15910_out0) || (!v$FF5_16957_out0) && v$FF6_15910_out0);
assign v$G24_12651_out0 = ! v$FF3_15648_out0;
assign v$G24_12652_out0 = ! v$FF3_15649_out0;
assign v$LASTQ_12664_out0 = v$FF2_13615_out0;
assign v$LASTQ_12665_out0 = v$FF2_13616_out0;
assign v$LASTQ_12666_out0 = v$FF2_13617_out0;
assign v$LASTQ_12667_out0 = v$FF2_13618_out0;
assign v$LASTQ_12668_out0 = v$FF2_13619_out0;
assign v$LASTQ_12669_out0 = v$FF2_13620_out0;
assign v$LASTQ_12670_out0 = v$FF2_13621_out0;
assign v$LASTQ_12671_out0 = v$FF2_13622_out0;
assign v$LASTQ_12672_out0 = v$FF2_13623_out0;
assign v$LASTQ_12673_out0 = v$FF2_13624_out0;
assign v$LASTQ_12674_out0 = v$FF2_13625_out0;
assign v$LASTQ_12675_out0 = v$FF2_13626_out0;
assign v$LASTQ_12676_out0 = v$FF2_13627_out0;
assign v$LASTQ_12677_out0 = v$FF2_13628_out0;
assign v$LASTQ_12678_out0 = v$FF2_13629_out0;
assign v$LASTQ_12679_out0 = v$FF2_13630_out0;
assign v$LASTQ_12680_out0 = v$FF2_13631_out0;
assign v$LASTQ_12681_out0 = v$FF2_13632_out0;
assign v$LASTQ_12682_out0 = v$FF2_13633_out0;
assign v$LASTQ_12683_out0 = v$FF2_13634_out0;
assign v$LASTQ_12684_out0 = v$FF2_13635_out0;
assign v$LASTQ_12685_out0 = v$FF2_13636_out0;
assign v$PCHALT_13316_out0 = v$REG1_9169_out0;
assign v$LEFT$SHIFT_13403_out0 = v$C11_3822_out0;
assign v$LEFT$SHIFT_13404_out0 = v$C2_17614_out0;
assign v$LEFT$SHIFT_13405_out0 = v$C3_1525_out0;
assign v$LEFT$SHIFT_13406_out0 = v$C3_18739_out0;
assign v$LEFT$SHIFT_13407_out0 = v$C11_3823_out0;
assign v$LEFT$SHIFT_13408_out0 = v$C2_17615_out0;
assign v$LEFT$SHIFT_13409_out0 = v$C3_1526_out0;
assign v$LEFT$SHIFT_13410_out0 = v$C3_18740_out0;
assign v$RMORIGINAL_13550_out0 = v$REG1_14711_out0;
assign v$RMORIGINAL_13551_out0 = v$REG1_14712_out0;
assign v$G1_13725_out0 = ! v$FF0_5223_out0;
assign v$G1_13726_out0 = ! v$FF0_5224_out0;
assign v$VALID$PREV_14013_out0 = v$FF14_11409_out0;
assign v$VALID$PREV_14014_out0 = v$FF14_11410_out0;
assign v$CARRY_14027_out0 = v$FF1_10761_out0;
assign v$CARRY_14028_out0 = v$FF1_10762_out0;
assign v$Q0_14284_out0 = v$FF0_716_out0;
assign v$Q0_14285_out0 = v$FF0_717_out0;
assign v$R1_14351_out0 = v$REG1_5110_out0;
assign v$R1_14352_out0 = v$REG1_5111_out0;
assign v$B$SHIFTED_14379_out0 = v$REG1_12653_out0;
assign v$B$SHIFTED_14380_out0 = v$REG1_12654_out0;
assign v$Q1_14930_out0 = v$FF1_2722_out0;
assign v$Q1_14931_out0 = v$FF1_2723_out0;
assign v$G1_15078_out0 = ! v$FF1_6306_out0;
assign v$G1_15079_out0 = ! v$FF1_6307_out0;
assign v$ADDRESS_15181_out0 = v$REG2_718_out0;
assign v$ADDRESS_15182_out0 = v$REG2_719_out0;
assign v$G5_15257_out0 = ((v$FF8_17348_out0 && !v$FF4_8562_out0) || (!v$FF8_17348_out0) && v$FF4_8562_out0);
assign v$G5_15258_out0 = ((v$FF8_17349_out0 && !v$FF4_8563_out0) || (!v$FF8_17349_out0) && v$FF4_8563_out0);
assign v$_15382_out0 = { v$FF1_9797_out0,v$FF2_3160_out0 };
assign v$_15383_out0 = { v$FF1_9798_out0,v$FF2_3161_out0 };
assign {v$A2_15432_out1,v$A2_15432_out0 } = v$REG2_718_out0 + v$C6_8360_out0 + v$C4_6606_out0;
assign {v$A2_15433_out1,v$A2_15433_out0 } = v$REG2_719_out0 + v$C6_8361_out0 + v$C4_6607_out0;
assign v$_15509_out0 = { v$FF1_16797_out0,v$FF2_1729_out0 };
assign v$_15510_out0 = { v$FF1_16798_out0,v$FF2_1730_out0 };
assign v$CIN_15669_out0 = v$C6_13145_out0;
assign v$CIN_15671_out0 = v$C5_16705_out0;
assign v$CIN_15672_out0 = v$C6_13146_out0;
assign v$CIN_15674_out0 = v$C5_16706_out0;
assign v$G71_15857_out0 = ! v$FF4_8369_out0;
assign v$G71_15858_out0 = ! v$FF4_8370_out0;
assign v$LSBS_15901_out0 = v$REG1_9225_out0;
assign v$LSBS_15902_out0 = v$REG1_9226_out0;
assign v$EQ1_15907_out0 = v$REG1_15444_out0 == 6'h1e;
assign v$EQ1_15908_out0 = v$REG1_15445_out0 == 6'h1e;
assign v$G3_16441_out0 = ((v$FF1_16797_out0 && !v$FF2_1729_out0) || (!v$FF1_16797_out0) && v$FF2_1729_out0);
assign v$G3_16442_out0 = ((v$FF1_16798_out0 && !v$FF2_1730_out0) || (!v$FF1_16798_out0) && v$FF2_1730_out0);
assign v$G52_16544_out0 = ! v$FF4_7301_out0;
assign v$G52_16545_out0 = ! v$FF4_7302_out0;
assign v$_16562_out0 = { v$FF5_16956_out0,v$FF6_15909_out0 };
assign v$_16563_out0 = { v$FF5_16957_out0,v$FF6_15910_out0 };
assign v$STATE_16624_out0 = v$FF1_5439_out0;
assign v$STATE_16625_out0 = v$FF1_5440_out0;
assign v$STATE_16626_out0 = v$FF1_5441_out0;
assign v$STATE_16627_out0 = v$FF1_5442_out0;
assign v$STATE_16628_out0 = v$FF1_5443_out0;
assign v$STATE_16629_out0 = v$FF1_5444_out0;
assign v$STATE_16630_out0 = v$REG1_7363_out0;
assign v$IR2_17178_out0 = v$REG4_6885_out0;
assign v$IR2_17179_out0 = v$REG4_6886_out0;
assign v$G24_17612_out0 = ((v$FF3_271_out0 && !v$FF4_2541_out0) || (!v$FF3_271_out0) && v$FF4_2541_out0);
assign v$G24_17613_out0 = ((v$FF3_272_out0 && !v$FF4_2542_out0) || (!v$FF3_272_out0) && v$FF4_2542_out0);
assign v$A_17640_out0 = v$REG1_14166_out0;
assign v$A_17641_out0 = v$REG1_14167_out0;
assign v$Q2_18125_out0 = v$FF2_4510_out0;
assign v$Q2_18126_out0 = v$FF2_4511_out0;
assign v$RD$OUT_18500_out0 = v$REG4_11270_out0;
assign v$RD$OUT_18501_out0 = v$REG4_11271_out0;
assign v$B_18591_out0 = v$REG2_16962_out0;
assign v$B_18592_out0 = v$REG2_16963_out0;
assign v$HALT$PREV$PREV_18681_out0 = v$FF12_17048_out0;
assign v$HALT$PREV$PREV_18682_out0 = v$FF12_17049_out0;
assign v$INT3_18737_out0 = v$C2_18926_out0;
assign v$INT3_18738_out0 = v$C2_18927_out0;
assign v$SOUT_18793_out0 = v$FF1_9797_out0;
assign v$SOUT_18794_out0 = v$FF1_9798_out0;
assign v$AUTODISABLE_18814_out0 = v$FF3_18727_out0;
assign v$AUTODISABLE_18815_out0 = v$FF3_18728_out0;
assign v$Q3_18893_out0 = v$FF3_16564_out0;
assign v$Q3_18894_out0 = v$FF3_16565_out0;
assign v$EPARITY_18914_out0 = v$FF9_16635_out0;
assign v$EPARITY_18915_out0 = v$FF9_16636_out0;
assign v$Q0_18924_out0 = v$FF0_4488_out0;
assign v$Q0_18925_out0 = v$FF0_4489_out0;
assign v$_19017_out0 = { v$FF5_19083_out0,v$FF3_1456_out0 };
assign v$_19018_out0 = { v$FF5_19084_out0,v$FF3_1457_out0 };
assign v$Q3_19033_out0 = v$FF3_11419_out0;
assign v$Q3_19034_out0 = v$FF3_11420_out0;
assign v$_19069_out0 = v$REG1_4200_out0[3:0];
assign v$_19069_out1 = v$REG1_4200_out0[7:4];
assign v$_19070_out0 = v$REG1_4201_out0[3:0];
assign v$_19070_out1 = v$REG1_4201_out0[7:4];
assign v$OUTPUT_19087_out0 = v$REG1_7363_out0;
assign v$G1_34_out0 = v$Wordlength_5358_out0 || v$G2_66_out0;
assign v$G1_35_out0 = v$Wordlength_5359_out0 || v$G2_67_out0;
assign v$SIN_92_out0 = v$SOUT1_2081_out0;
assign v$SIN_93_out0 = v$SOUT1_2084_out0;
assign v$SIN_94_out0 = v$SOUT1_2085_out0;
assign v$SIN_96_out0 = v$SOUT1_2083_out0;
assign v$SIN_97_out0 = v$SOUT1_2080_out0;
assign v$SIN_98_out0 = v$SOUT1_2087_out0;
assign v$SIN_99_out0 = v$SOUT1_2090_out0;
assign v$SIN_100_out0 = v$SOUT1_2091_out0;
assign v$SIN_102_out0 = v$SOUT1_2089_out0;
assign v$SIN_103_out0 = v$SOUT1_2086_out0;
assign v$CALCULATING_1647_out0 = v$OUTPUT_10799_out0;
assign v$CALCULATING_1648_out0 = v$OUTPUT_10802_out0;
assign v$_1683_out0 = v$A_17640_out0[7:0];
assign v$_1683_out1 = v$A_17640_out0[15:8];
assign v$_1684_out0 = v$A_17641_out0[7:0];
assign v$_1684_out1 = v$A_17641_out0[15:8];
assign v$G1_1750_out0 = ! v$Q0_18924_out0;
assign v$G1_1751_out0 = ! v$Q0_18925_out0;
assign v$IR2_1911_out0 = v$IR2_17178_out0;
assign v$IR2_1912_out0 = v$IR2_17179_out0;
assign v$_1989_out0 = { v$Q0_18924_out0,v$Q1_4619_out0 };
assign v$_1990_out0 = { v$Q0_18925_out0,v$Q1_4620_out0 };
assign v$G8_2473_out0 = ! v$Q1_14930_out0;
assign v$G8_2474_out0 = ! v$Q1_14931_out0;
assign v$I1P_2710_out0 = v$I1P_6684_out0;
assign v$I1P_2711_out0 = v$I1P_6685_out0;
assign v$IR2_3141_out0 = v$IR2_17178_out0;
assign v$IR2_3142_out0 = v$IR2_17179_out0;
assign {v$A1_3146_out1,v$A1_3146_out0 } = v$D_6009_out0 + v$C1_5455_out0 + v$C2_11198_out0;
assign {v$A1_3147_out1,v$A1_3147_out0 } = v$D_6010_out0 + v$C1_5456_out0 + v$C2_11199_out0;
assign v$G18_3199_out0 = ! v$ISINTERRUPTED_12429_out0;
assign v$G18_3200_out0 = ! v$ISINTERRUPTED_12430_out0;
assign v$END4_3491_out0 = v$LASTQ_12674_out0;
assign v$END4_3492_out0 = v$LASTQ_12685_out0;
assign v$G6_3580_out0 = ((v$Q0_74_out0 && !v$Q1_14930_out0) || (!v$Q0_74_out0) && v$Q1_14930_out0);
assign v$G6_3581_out0 = ((v$Q0_75_out0 && !v$Q1_14931_out0) || (!v$Q0_75_out0) && v$Q1_14931_out0);
assign v$INTERRUPT3_3708_out0 = v$INT3_18737_out0;
assign v$INTERRUPT3_3709_out0 = v$INT3_18738_out0;
assign v$B$SAVED_4066_out0 = v$B$SAVED_4961_out0;
assign v$B$SAVED_4067_out0 = v$B$SAVED_4962_out0;
assign v$_4140_out0 = v$B2_8720_out0[11:0];
assign v$_4140_out1 = v$B2_8720_out0[23:12];
assign v$_4143_out0 = v$B2_8723_out0[11:0];
assign v$_4143_out1 = v$B2_8723_out0[23:12];
assign v$OFF_4196_out0 = v$EQ1_7213_out0;
assign v$OFF_4197_out0 = v$EQ1_7214_out0;
assign v$G22_4474_out0 = ((v$Q1_11427_out0 && !v$Q0_14284_out0) || (!v$Q1_11427_out0) && v$Q0_14284_out0);
assign v$G22_4475_out0 = ((v$Q1_11428_out0 && !v$Q0_14285_out0) || (!v$Q1_11428_out0) && v$Q0_14285_out0);
assign v$G35_4476_out0 = v$Q1_4619_out0 && v$Q0_18924_out0;
assign v$G35_4477_out0 = v$Q1_4620_out0 && v$Q0_18925_out0;
assign v$I0P_4512_out0 = v$I0P_10763_out0;
assign v$I0P_4513_out0 = v$I0P_10764_out0;
assign v$B$SAVED_4522_out0 = v$B$SAVED_4961_out0;
assign v$B$SAVED_4523_out0 = v$B$SAVED_4962_out0;
assign v$G48_5092_out0 = ! v$STALL$PREV$CYCLE_6059_out0;
assign v$G48_5093_out0 = ! v$STALL$PREV$CYCLE_6060_out0;
assign v$G87_5362_out0 = ! v$PHALT0_12199_out0;
assign v$_5715_out0 = { v$_15382_out0,v$_8051_out0 };
assign v$_5716_out0 = { v$_15383_out0,v$_8052_out0 };
assign v$_5759_out0 = { v$_19017_out0,v$_15509_out0 };
assign v$_5760_out0 = { v$_19018_out0,v$_15510_out0 };
assign v$SERIALIN_6011_out0 = v$SOUT_18793_out0;
assign v$SERIALIN_6012_out0 = v$SOUT_18794_out0;
assign v$PIPELINE$RESTART_6348_out0 = v$PIPELINERESTART_2611_out0;
assign v$PIPELINE$RESTART_6349_out0 = v$PIPELINERESTART_2612_out0;
assign v$RECIEVEDPARITY_6488_out0 = v$RecievedParity_9916_out0;
assign v$RECIEVEDPARITY_6489_out0 = v$RecievedParity_9917_out0;
assign v$G64_6638_out0 = v$HALT$PREV_10837_out0 && v$STALL$PREV$PREV_6096_out0;
assign v$G64_6639_out0 = v$HALT$PREV_10838_out0 && v$STALL$PREV$PREV_6097_out0;
assign v$END1_7241_out0 = v$LASTQ_12673_out0;
assign v$END1_7242_out0 = v$LASTQ_12684_out0;
assign v$END1_7268_out0 = v$A2_15432_out1;
assign v$END1_7269_out0 = v$A2_15433_out1;
assign v$_7307_out0 = { v$_16562_out0,v$_2471_out0 };
assign v$_7308_out0 = { v$_16563_out0,v$_2472_out0 };
assign v$G22_7584_out0 = ((v$G21_12447_out0 && !v$G20_7717_out0) || (!v$G21_12447_out0) && v$G20_7717_out0);
assign v$G22_7585_out0 = ((v$G21_12448_out0 && !v$G20_7718_out0) || (!v$G21_12448_out0) && v$G20_7718_out0);
assign v$I2P_7810_out0 = v$I2P_2465_out0;
assign v$I2P_7811_out0 = v$I2P_2466_out0;
assign v$R3TEST_7858_out0 = v$R3_11234_out0;
assign v$R3TEST_7859_out0 = v$R3_11235_out0;
assign v$END6_7866_out0 = v$LASTQ_12668_out0;
assign v$END6_7867_out0 = v$LASTQ_12679_out0;
assign v$G2_7886_out0 = ! v$OUTPUT_19087_out0;
assign v$CALCULATING_8122_out0 = v$OUTPUT_10800_out0;
assign v$CALCULATING_8123_out0 = v$OUTPUT_10803_out0;
assign v$G7_8168_out0 = ! v$Q3_18893_out0;
assign v$G7_8169_out0 = ! v$Q3_18894_out0;
assign v$DM1_8182_out0 = v$SELOUT_1880_out0 ? 16'h0 : v$RAM1_13483_out0;
assign v$DM1_8182_out1 = v$SELOUT_1880_out0 ? v$RAM1_13483_out0 : 16'h0;
assign v$RXDISABLE_8214_out0 = v$_5112_out1;
assign v$RXDISABLE_8215_out0 = v$_5113_out1;
assign v$G3_8354_out0 = v$FF1_194_out0 || v$G2_66_out0;
assign v$G3_8355_out0 = v$FF1_195_out0 || v$G2_67_out0;
assign v$END_8410_out0 = v$A1_4168_out1;
assign v$END_8411_out0 = v$A1_4169_out1;
assign v$_8414_out0 = { v$_1429_out0,v$Q2_3367_out0 };
assign v$_8415_out0 = { v$_1430_out0,v$Q2_3368_out0 };
assign v$END4_8432_out0 = v$LASTQ_12665_out0;
assign v$END4_8433_out0 = v$LASTQ_12676_out0;
assign v$R0TEST_8545_out0 = v$R0_3503_out0;
assign v$R0TEST_8546_out0 = v$R0_3504_out0;
assign v$LEFT$SHIFT_9143_out0 = v$LEFT$SHIFT_13403_out0;
assign v$LEFT$SHIFT_9144_out0 = v$LEFT$SHIFT_13404_out0;
assign v$LEFT$SHIFT_9145_out0 = v$LEFT$SHIFT_13405_out0;
assign v$LEFT$SHIFT_9146_out0 = v$LEFT$SHIFT_13406_out0;
assign v$LEFT$SHIFT_9147_out0 = v$LEFT$SHIFT_13407_out0;
assign v$LEFT$SHIFT_9148_out0 = v$LEFT$SHIFT_13408_out0;
assign v$LEFT$SHIFT_9149_out0 = v$LEFT$SHIFT_13409_out0;
assign v$LEFT$SHIFT_9150_out0 = v$LEFT$SHIFT_13410_out0;
assign v$_9303_out0 = v$B_18591_out0[7:0];
assign v$_9303_out1 = v$B_18591_out0[15:8];
assign v$_9304_out0 = v$B_18592_out0[7:0];
assign v$_9304_out1 = v$B_18592_out0[15:8];
assign v$G6_9404_out0 = ! v$Q2_5696_out0;
assign v$G6_9405_out0 = ! v$Q2_5697_out0;
assign v$MODE_9454_out0 = v$_5112_out0;
assign v$MODE_9455_out0 = v$_5113_out0;
assign v$A$SAVED_10392_out0 = v$A$SAVED_3877_out0;
assign v$A$SAVED_10393_out0 = v$A$SAVED_3878_out0;
assign v$G38_10705_out0 = v$Q0_18924_out0 || v$Q1_4619_out0;
assign v$G38_10706_out0 = v$Q0_18925_out0 || v$Q1_4620_out0;
assign v$INIT_11241_out0 = v$G2_66_out0;
assign v$INIT_11242_out0 = v$G2_67_out0;
assign v$_11306_out0 = v$_19069_out0[1:0];
assign v$_11306_out1 = v$_19069_out0[3:2];
assign v$_11307_out0 = v$_19070_out0[1:0];
assign v$_11307_out1 = v$_19070_out0[3:2];
assign v$I3P_11324_out0 = v$I3P_9295_out0;
assign v$I3P_11325_out0 = v$I3P_9296_out0;
assign v$CARRY_11411_out0 = v$CARRY_14027_out0;
assign v$CARRY_11412_out0 = v$CARRY_14028_out0;
assign v$TXLast_11914_out0 = v$LASTQ_12670_out0;
assign v$TXLast_11915_out0 = v$LASTQ_12681_out0;
assign v$G57_12214_out0 = ! v$HALT$PREV_10837_out0;
assign v$G57_12215_out0 = ! v$HALT$PREV_10838_out0;
assign v$G27_12274_out0 = v$Q0_14284_out0 && v$Q1_11427_out0;
assign v$G27_12275_out0 = v$Q0_14285_out0 && v$Q1_11428_out0;
assign v$_12388_out0 = v$_19069_out1[1:0];
assign v$_12388_out1 = v$_19069_out1[3:2];
assign v$_12389_out0 = v$_19070_out1[1:0];
assign v$_12389_out1 = v$_19070_out1[3:2];
assign v$HALTED_12399_out0 = v$OUTPUT_10801_out0;
assign v$HALTED_12400_out0 = v$OUTPUT_10804_out0;
assign v$INSTR$READ1_12546_out0 = v$OUT_8651_out0;
assign v$RXlast_13391_out0 = v$LASTQ_12671_out0;
assign v$RXlast_13392_out0 = v$LASTQ_12682_out0;
assign v$RD$FPU_13518_out0 = v$RD$OUT_18500_out0;
assign v$RD$FPU_13519_out0 = v$RD$OUT_18501_out0;
assign v$G6_13585_out0 = ((v$G2_1447_out0 && !v$G3_16441_out0) || (!v$G2_1447_out0) && v$G3_16441_out0);
assign v$G6_13586_out0 = ((v$G2_1448_out0 && !v$G3_16442_out0) || (!v$G2_1448_out0) && v$G3_16442_out0);
assign v$_13995_out0 = { v$Q2_18125_out0,v$Q3_19033_out0 };
assign v$_13996_out0 = { v$Q2_18126_out0,v$Q3_19034_out0 };
assign v$G7_14015_out0 = ((v$G4_3096_out0 && !v$G5_15257_out0) || (!v$G4_3096_out0) && v$G5_15257_out0);
assign v$G7_14016_out0 = ((v$G4_3097_out0 && !v$G5_15258_out0) || (!v$G4_3097_out0) && v$G5_15258_out0);
assign v$G86_14102_out0 = ! v$PHALT1_9264_out0;
assign v$EVENPARITY_14162_out0 = v$EPARITY_18914_out0;
assign v$EVENPARITY_14163_out0 = v$EPARITY_18915_out0;
assign v$G4_14607_out0 = ! v$Q0_14284_out0;
assign v$G4_14608_out0 = ! v$Q0_14285_out0;
assign v$G51_14624_out0 = ! v$HALT$PREV_10837_out0;
assign v$G51_14625_out0 = ! v$HALT$PREV_10838_out0;
assign v$G25_14641_out0 = ((v$Q0_18924_out0 && !v$Q1_4619_out0) || (!v$Q0_18924_out0) && v$Q1_4619_out0);
assign v$G25_14642_out0 = ((v$Q0_18925_out0 && !v$Q1_4620_out0) || (!v$Q0_18925_out0) && v$Q1_4620_out0);
assign v$INSTR$READ0_14785_out0 = v$OUT_5477_out0;
assign v$G7_14914_out0 = ! v$Q2_3367_out0;
assign v$G7_14915_out0 = ! v$Q2_3368_out0;
assign v$A$SAVED_15235_out0 = v$A$SAVED_3877_out0;
assign v$A$SAVED_15236_out0 = v$A$SAVED_3878_out0;
assign v$PHALT_15747_out0 = v$PHALT_1794_out0;
assign v$R1TEST_15756_out0 = v$R1_14351_out0;
assign v$R1TEST_15757_out0 = v$R1_14352_out0;
assign v$R2TEST_16315_out0 = v$R2_8285_out0;
assign v$R2TEST_16316_out0 = v$R2_8286_out0;
assign v$G2_16361_out0 = ! v$Q1_4619_out0;
assign v$G2_16362_out0 = ! v$Q1_4620_out0;
assign v$G25_16715_out0 = ((v$G23_9729_out0 && !v$G24_17612_out0) || (!v$G23_9729_out0) && v$G24_17612_out0);
assign v$G25_16716_out0 = ((v$G23_9730_out0 && !v$G24_17613_out0) || (!v$G23_9730_out0) && v$G24_17613_out0);
assign v$_16740_out0 = { v$_3967_out0,v$_9811_out0 };
assign v$_16741_out0 = { v$_3968_out0,v$_9812_out0 };
assign v$G5_16764_out0 = ! v$Q1_11427_out0;
assign v$G5_16765_out0 = ! v$Q1_11428_out0;
v$AROM1_16768 I16768 (v$AROM1_16768_out0, v$ADDRESS_15181_out0);
v$AROM1_16769 I16769 (v$AROM1_16769_out0, v$ADDRESS_15182_out0);
assign v$G61_17069_out0 = ! v$HALT$PREV_10837_out0;
assign v$G61_17070_out0 = ! v$HALT$PREV_10838_out0;
assign v$G9_17120_out0 = ! v$Q0_74_out0;
assign v$G9_17121_out0 = ! v$Q0_75_out0;
assign v$PCHALT_17182_out0 = v$PCHALT_13316_out0;
assign v$CLK4_17354_out0 = v$G3_20_out0;
assign v$CLK4_17355_out0 = v$G3_21_out0;
assign v$END_17644_out0 = v$LASTQ_12672_out0;
assign v$END_17645_out0 = v$LASTQ_12683_out0;
assign v$CIN_17983_out0 = v$CIN_15669_out0;
assign v$CIN_17985_out0 = v$CIN_15671_out0;
assign v$CIN_17986_out0 = v$CIN_15672_out0;
assign v$CIN_17988_out0 = v$CIN_15674_out0;
assign v$G4_18209_out0 = ! v$Q3_19033_out0;
assign v$G4_18210_out0 = ! v$Q3_19034_out0;
assign v$increment_18454_out0 = v$EQ1_15907_out0;
assign v$increment_18455_out0 = v$EQ1_15908_out0;
assign v$G55_18799_out0 = ! v$HALT$PREV_10837_out0;
assign v$G55_18800_out0 = ! v$HALT$PREV_10838_out0;
assign v$_18932_out0 = { v$Q2_5696_out0,v$Q3_18893_out0 };
assign v$_18933_out0 = { v$Q2_5697_out0,v$Q3_18894_out0 };
assign v$G3_19021_out0 = ! v$Q2_18125_out0;
assign v$G3_19022_out0 = ! v$Q2_18126_out0;
assign v$G41_19089_out0 = v$Q0_18924_out0 && v$Q1_4619_out0;
assign v$G41_19090_out0 = v$Q0_18925_out0 && v$Q1_4620_out0;
assign v$_19129_out0 = { v$Q0_14284_out0,v$Q1_11427_out0 };
assign v$_19130_out0 = { v$Q0_14285_out0,v$Q1_11428_out0 };
assign v$NQ1_263_out0 = v$G5_16764_out0;
assign v$NQ1_264_out0 = v$G5_16765_out0;
assign v$SEL5_704_out0 = v$IR2_1911_out0[11:10];
assign v$SEL5_705_out0 = v$IR2_1912_out0[11:10];
assign v$G1_1343_out0 = ! v$OFF_4196_out0;
assign v$G1_1344_out0 = ! v$OFF_4197_out0;
assign v$_1369_out0 = v$_4140_out1[5:0];
assign v$_1369_out1 = v$_4140_out1[11:6];
assign v$_1372_out0 = v$_4143_out1[5:0];
assign v$_1372_out1 = v$_4143_out1[11:6];
assign v$NQ3_1645_out0 = v$G7_8168_out0;
assign v$NQ3_1646_out0 = v$G7_8169_out0;
assign v$_1677_out0 = v$_4140_out0[5:0];
assign v$_1677_out1 = v$_4140_out0[11:6];
assign v$_1680_out0 = v$_4143_out0[5:0];
assign v$_1680_out1 = v$_4143_out0[11:6];
assign v$MODE_1773_out0 = v$MODE_9454_out0;
assign v$MODE_1774_out0 = v$MODE_9455_out0;
assign v$IR2_2422_out0 = v$IR2_3141_out0;
assign v$IR2_2423_out0 = v$IR2_3142_out0;
assign v$_2539_out0 = v$_9303_out0[3:0];
assign v$_2539_out1 = v$_9303_out0[7:4];
assign v$_2540_out0 = v$_9304_out0[3:0];
assign v$_2540_out1 = v$_9304_out0[7:4];
assign v$G58_2714_out0 = v$FF11_2642_out0 && v$G57_12214_out0;
assign v$G58_2715_out0 = v$FF11_2643_out0 && v$G57_12215_out0;
assign v$_3104_out0 = v$_9303_out1[3:0];
assign v$_3104_out1 = v$_9303_out1[7:4];
assign v$_3105_out0 = v$_9304_out1[3:0];
assign v$_3105_out1 = v$_9304_out1[7:4];
assign v$NQ2_3191_out0 = v$G6_9404_out0;
assign v$NQ2_3192_out0 = v$G6_9405_out0;
assign v$NQ3_3209_out0 = v$G4_18209_out0;
assign v$NQ3_3210_out0 = v$G4_18210_out0;
assign v$LEFT$SHIT_3255_out0 = v$LEFT$SHIFT_9143_out0;
assign v$LEFT$SHIT_3256_out0 = v$LEFT$SHIFT_9143_out0;
assign v$LEFT$SHIT_3257_out0 = v$LEFT$SHIFT_9143_out0;
assign v$LEFT$SHIT_3258_out0 = v$LEFT$SHIFT_9143_out0;
assign v$LEFT$SHIT_3259_out0 = v$LEFT$SHIFT_9143_out0;
assign v$LEFT$SHIT_3260_out0 = v$LEFT$SHIFT_9144_out0;
assign v$LEFT$SHIT_3261_out0 = v$LEFT$SHIFT_9144_out0;
assign v$LEFT$SHIT_3262_out0 = v$LEFT$SHIFT_9144_out0;
assign v$LEFT$SHIT_3263_out0 = v$LEFT$SHIFT_9144_out0;
assign v$LEFT$SHIT_3264_out0 = v$LEFT$SHIFT_9144_out0;
assign v$LEFT$SHIT_3265_out0 = v$LEFT$SHIFT_9145_out0;
assign v$LEFT$SHIT_3266_out0 = v$LEFT$SHIFT_9145_out0;
assign v$LEFT$SHIT_3267_out0 = v$LEFT$SHIFT_9145_out0;
assign v$LEFT$SHIT_3268_out0 = v$LEFT$SHIFT_9145_out0;
assign v$LEFT$SHIT_3269_out0 = v$LEFT$SHIFT_9145_out0;
assign v$LEFT$SHIT_3275_out0 = v$LEFT$SHIFT_9146_out0;
assign v$LEFT$SHIT_3276_out0 = v$LEFT$SHIFT_9146_out0;
assign v$LEFT$SHIT_3277_out0 = v$LEFT$SHIFT_9146_out0;
assign v$LEFT$SHIT_3278_out0 = v$LEFT$SHIFT_9146_out0;
assign v$LEFT$SHIT_3279_out0 = v$LEFT$SHIFT_9146_out0;
assign v$LEFT$SHIT_3286_out0 = v$LEFT$SHIFT_9147_out0;
assign v$LEFT$SHIT_3287_out0 = v$LEFT$SHIFT_9147_out0;
assign v$LEFT$SHIT_3288_out0 = v$LEFT$SHIFT_9147_out0;
assign v$LEFT$SHIT_3289_out0 = v$LEFT$SHIFT_9147_out0;
assign v$LEFT$SHIT_3290_out0 = v$LEFT$SHIFT_9147_out0;
assign v$LEFT$SHIT_3291_out0 = v$LEFT$SHIFT_9148_out0;
assign v$LEFT$SHIT_3292_out0 = v$LEFT$SHIFT_9148_out0;
assign v$LEFT$SHIT_3293_out0 = v$LEFT$SHIFT_9148_out0;
assign v$LEFT$SHIT_3294_out0 = v$LEFT$SHIFT_9148_out0;
assign v$LEFT$SHIT_3295_out0 = v$LEFT$SHIFT_9148_out0;
assign v$LEFT$SHIT_3296_out0 = v$LEFT$SHIFT_9149_out0;
assign v$LEFT$SHIT_3297_out0 = v$LEFT$SHIFT_9149_out0;
assign v$LEFT$SHIT_3298_out0 = v$LEFT$SHIFT_9149_out0;
assign v$LEFT$SHIT_3299_out0 = v$LEFT$SHIFT_9149_out0;
assign v$LEFT$SHIT_3300_out0 = v$LEFT$SHIFT_9149_out0;
assign v$LEFT$SHIT_3306_out0 = v$LEFT$SHIFT_9150_out0;
assign v$LEFT$SHIT_3307_out0 = v$LEFT$SHIFT_9150_out0;
assign v$LEFT$SHIT_3308_out0 = v$LEFT$SHIFT_9150_out0;
assign v$LEFT$SHIT_3309_out0 = v$LEFT$SHIFT_9150_out0;
assign v$LEFT$SHIT_3310_out0 = v$LEFT$SHIFT_9150_out0;
assign v$_3322_out0 = v$_12388_out1[0:0];
assign v$_3322_out1 = v$_12388_out1[1:1];
assign v$_3323_out0 = v$_12389_out1[0:0];
assign v$_3323_out1 = v$_12389_out1[1:1];
assign v$_3864_out0 = v$_11306_out1[0:0];
assign v$_3864_out1 = v$_11306_out1[1:1];
assign v$_3865_out0 = v$_11307_out1[0:0];
assign v$_3865_out1 = v$_11307_out1[1:1];
assign v$XOR1_4124_out0 = v$A1_3146_out0 ^ v$C3_7297_out0;
assign v$XOR1_4125_out0 = v$A1_3147_out0 ^ v$C3_7298_out0;
assign v$SEL13_5054_out0 = v$IR2_1911_out0[9:8];
assign v$SEL13_5055_out0 = v$IR2_1912_out0[9:8];
assign v$CARRY_5219_out0 = v$CARRY_11411_out0;
assign v$CARRY_5220_out0 = v$CARRY_11412_out0;
assign v$_5293_out0 = v$_12388_out0[0:0];
assign v$_5293_out1 = v$_12388_out0[1:1];
assign v$_5294_out0 = v$_12389_out0[0:0];
assign v$_5294_out1 = v$_12389_out0[1:1];
assign v$_6707_out0 = v$_1683_out1[3:0];
assign v$_6707_out1 = v$_1683_out1[7:4];
assign v$_6708_out0 = v$_1684_out1[3:0];
assign v$_6708_out1 = v$_1684_out1[7:4];
assign v$_7264_out0 = v$_11306_out0[0:0];
assign v$_7264_out1 = v$_11306_out0[1:1];
assign v$_7265_out0 = v$_11307_out0[0:0];
assign v$_7265_out1 = v$_11307_out0[1:1];
assign v$SEL4_7339_out0 = v$IR2_1911_out0[15:15];
assign v$SEL4_7340_out0 = v$IR2_1912_out0[15:15];
assign v$CLK4_7347_out0 = v$CLK4_17354_out0;
assign v$CLK4_7348_out0 = v$CLK4_17355_out0;
assign v$INSTR$READ_7535_out0 = v$INSTR$READ1_12546_out0;
assign v$INSTR$READ_7536_out0 = v$INSTR$READ0_14785_out0;
assign v$SEL10_7597_out0 = v$IR2_1911_out0[9:9];
assign v$SEL10_7598_out0 = v$IR2_1912_out0[9:9];
assign v$NQ0_8120_out0 = v$G4_14607_out0;
assign v$NQ0_8121_out0 = v$G4_14608_out0;
assign v$RAMDOUT1_8627_out0 = v$DM1_8182_out1;
assign v$SEL11_8654_out0 = v$IR2_1911_out0[8:8];
assign v$SEL11_8655_out0 = v$IR2_1912_out0[8:8];
assign v$_8712_out0 = v$_1683_out0[3:0];
assign v$_8712_out1 = v$_1683_out0[7:4];
assign v$_8713_out0 = v$_1684_out0[3:0];
assign v$_8713_out1 = v$_1684_out0[7:4];
assign v$G65_9154_out0 = ! v$PHALT_15747_out0;
assign v$_9265_out0 = { v$_19129_out0,v$_18932_out0 };
assign v$_9266_out0 = { v$_19130_out0,v$_18933_out0 };
assign v$RAMDOUT0_9426_out0 = v$DM1_8182_out0;
assign v$G3_9809_out0 = ! v$RXDISABLE_8214_out0;
assign v$G3_9810_out0 = ! v$RXDISABLE_8215_out0;
assign v$_10354_out0 = v$AROM1_16768_out0[27:0];
assign v$_10354_out1 = v$AROM1_16768_out0[43:16];
assign v$_10355_out0 = v$AROM1_16769_out0[27:0];
assign v$_10355_out1 = v$AROM1_16769_out0[43:16];
assign v$_10703_out0 = { v$_1989_out0,v$_13995_out0 };
assign v$_10704_out0 = { v$_1990_out0,v$_13996_out0 };
assign v$G25_10727_out0 = ! v$CALCULATING_8122_out0;
assign v$G25_10728_out0 = ! v$CALCULATING_8123_out0;
assign v$Mode_11483_out0 = v$MODE_9454_out0;
assign v$Mode_11484_out0 = v$MODE_9455_out0;
assign v$G3_11496_out0 = ! v$OFF_4196_out0;
assign v$G3_11497_out0 = ! v$OFF_4197_out0;
assign v$NQ1_11550_out0 = v$G2_16361_out0;
assign v$NQ1_11551_out0 = v$G2_16362_out0;
assign v$G8_12863_out0 = ((v$G6_13585_out0 && !v$G7_14015_out0) || (!v$G6_13585_out0) && v$G7_14015_out0);
assign v$G8_12864_out0 = ((v$G6_13586_out0 && !v$G7_14016_out0) || (!v$G6_13586_out0) && v$G7_14016_out0);
assign v$SEL12_13371_out0 = v$IR2_1911_out0[15:12];
assign v$SEL12_13372_out0 = v$IR2_1912_out0[15:12];
assign v$Mode_13777_out0 = v$MODE_9454_out0;
assign v$Mode_13778_out0 = v$MODE_9455_out0;
assign v$EQ1_13938_out0 = v$_8414_out0 == 3'h0;
assign v$EQ1_13939_out0 = v$_8415_out0 == 3'h0;
assign v$COUT_14088_out0 = v$A1_3146_out1;
assign v$COUT_14089_out0 = v$A1_3147_out1;
assign v$G67_14340_out0 = ! v$PHALT_15747_out0;
assign v$G70_14638_out0 = v$PCHALT_17182_out0 && v$PHALT_15747_out0;
assign v$G67_14719_out0 = v$HALTED_12399_out0 && v$VALID$PREV_14013_out0;
assign v$G67_14720_out0 = v$HALTED_12400_out0 && v$VALID$PREV_14014_out0;
assign v$G4_14816_out0 = v$SOUT1_2082_out0 || v$INIT_11241_out0;
assign v$G4_14817_out0 = v$SOUT1_2088_out0 || v$INIT_11242_out0;
assign v$_15255_out0 = { v$_5715_out0,v$_7307_out0 };
assign v$_15256_out0 = { v$_5716_out0,v$_7308_out0 };
assign v$HALTSEL_15349_out0 = v$G2_7886_out0;
assign v$NQ0_15970_out0 = v$G9_17120_out0;
assign v$NQ0_15971_out0 = v$G9_17121_out0;
assign v$NQ0_16214_out0 = v$G1_1750_out0;
assign v$NQ0_16215_out0 = v$G1_1751_out0;
assign v$_16264_out0 = { v$_5759_out0,v$_16740_out0 };
assign v$_16265_out0 = { v$_5760_out0,v$_16741_out0 };
assign v$G69_16415_out0 = v$PCHALT_17182_out0 && v$PHALT_15747_out0;
assign v$G26_16633_out0 = ((v$G25_16715_out0 && !v$G22_7584_out0) || (!v$G25_16715_out0) && v$G22_7584_out0);
assign v$G26_16634_out0 = ((v$G25_16716_out0 && !v$G22_7585_out0) || (!v$G25_16716_out0) && v$G22_7585_out0);
assign v$CIN_16717_out0 = v$CIN_17983_out0;
assign v$CIN_16719_out0 = v$CIN_17985_out0;
assign v$CIN_16720_out0 = v$CIN_17986_out0;
assign v$CIN_16722_out0 = v$CIN_17988_out0;
assign v$NQ2_17316_out0 = v$G7_14914_out0;
assign v$NQ2_17317_out0 = v$G7_14915_out0;
assign v$NQ1_17350_out0 = v$G8_2473_out0;
assign v$NQ1_17351_out0 = v$G8_2474_out0;
assign v$PHALT_18124_out0 = v$G2_7886_out0;
assign v$CLEAR_19011_out0 = v$G1_34_out0;
assign v$CLEAR_19012_out0 = v$G1_35_out0;
assign v$RceivedParity_19151_out0 = v$RECIEVEDPARITY_6488_out0;
assign v$RceivedParity_19152_out0 = v$RECIEVEDPARITY_6489_out0;
assign v$NQ2_19175_out0 = v$G3_19021_out0;
assign v$NQ2_19176_out0 = v$G3_19022_out0;
assign v$PIPELINE$RESTART_19235_out0 = v$PIPELINE$RESTART_6348_out0;
assign v$PIPELINE$RESTART_19236_out0 = v$PIPELINE$RESTART_6349_out0;
assign v$_218_out0 = v$_8712_out1[1:0];
assign v$_218_out1 = v$_8712_out1[3:2];
assign v$_219_out0 = v$_8713_out1[1:0];
assign v$_219_out1 = v$_8713_out1[3:2];
assign v$G43_409_out0 = v$NQ2_19175_out0 && v$Q3_19033_out0;
assign v$G43_410_out0 = v$NQ2_19176_out0 && v$Q3_19034_out0;
assign v$G37_748_out0 = v$NQ0_8120_out0 || v$NQ1_263_out0;
assign v$G37_749_out0 = v$NQ0_8121_out0 || v$NQ1_264_out0;
assign v$S_1377_out0 = v$PHALT_18124_out0;
assign v$RXCLK_1393_out0 = v$EQ1_13938_out0;
assign v$RXCLK_1394_out0 = v$EQ1_13939_out0;
assign v$EQ12_1693_out0 = v$SEL12_13371_out0 == 4'h0;
assign v$EQ12_1694_out0 = v$SEL12_13372_out0 == 4'h0;
assign v$_1761_out0 = v$_6707_out1[1:0];
assign v$_1761_out1 = v$_6707_out1[3:2];
assign v$_1762_out0 = v$_6708_out1[1:0];
assign v$_1762_out1 = v$_6708_out1[3:2];
assign v$_1829_out0 = v$_10354_out1[7:0];
assign v$_1829_out1 = v$_10354_out1[15:8];
assign v$_1830_out0 = v$_10355_out1[7:0];
assign v$_1830_out1 = v$_10355_out1[15:8];
assign v$G54_2064_out0 = v$NQ1_263_out0 && v$NQ0_8120_out0;
assign v$G54_2065_out0 = v$NQ1_264_out0 && v$NQ0_8121_out0;
assign v$G23_2483_out0 = v$NQ3_1645_out0 || v$NQ2_3191_out0;
assign v$G23_2484_out0 = v$NQ3_1646_out0 || v$NQ2_3192_out0;
assign v$_2493_out0 = v$_2539_out0[1:0];
assign v$_2493_out1 = v$_2539_out0[3:2];
assign v$_2494_out0 = v$_2540_out0[1:0];
assign v$_2494_out1 = v$_2540_out0[3:2];
assign v$G19_2605_out0 = v$NQ1_263_out0 && v$NQ2_3191_out0;
assign v$G19_2606_out0 = v$NQ1_264_out0 && v$NQ2_3192_out0;
assign v$G51_3076_out0 = v$Q3_18893_out0 && v$NQ2_3191_out0;
assign v$G51_3077_out0 = v$Q3_18894_out0 && v$NQ2_3192_out0;
assign v$G16_3233_out0 = v$NQ1_17350_out0 && v$Q2_3367_out0;
assign v$G16_3234_out0 = v$NQ1_17351_out0 && v$Q2_3368_out0;
assign v$G56_3361_out0 = v$NQ3_1645_out0 && v$Q0_14284_out0;
assign v$G56_3362_out0 = v$NQ3_1646_out0 && v$Q0_14285_out0;
assign v$Write_3479_out0 = v$CLEAR_19011_out0;
assign v$Write_3480_out0 = v$CLEAR_19011_out0;
assign v$Write_3481_out0 = v$CLEAR_19011_out0;
assign v$Write_3482_out0 = v$CLEAR_19011_out0;
assign v$Write_3483_out0 = v$CLEAR_19011_out0;
assign v$Write_3484_out0 = v$CLEAR_19011_out0;
assign v$Write_3485_out0 = v$CLEAR_19012_out0;
assign v$Write_3486_out0 = v$CLEAR_19012_out0;
assign v$Write_3487_out0 = v$CLEAR_19012_out0;
assign v$Write_3488_out0 = v$CLEAR_19012_out0;
assign v$Write_3489_out0 = v$CLEAR_19012_out0;
assign v$Write_3490_out0 = v$CLEAR_19012_out0;
assign v$F1_3687_out0 = v$_5293_out1;
assign v$F1_3688_out0 = v$_5294_out1;
assign v$C_3832_out0 = v$CARRY_5219_out0;
assign v$C_3833_out0 = v$CARRY_5220_out0;
assign v$CLK4_3873_out0 = v$CLK4_7347_out0;
assign v$CLK4_3874_out0 = v$CLK4_7348_out0;
assign v$RXENABLE_3897_out0 = v$G3_9809_out0;
assign v$RXENABLE_3898_out0 = v$G3_9810_out0;
assign v$G59_4024_out0 = v$Q2_18125_out0 && v$NQ3_3209_out0;
assign v$G59_4025_out0 = v$Q2_18126_out0 && v$NQ3_3210_out0;
assign v$R2_4026_out0 = v$_3864_out0;
assign v$R2_4027_out0 = v$_3865_out0;
assign v$IR2_4118_out0 = v$IR2_2422_out0;
assign v$IR2_4119_out0 = v$IR2_2423_out0;
assign v$G26_4254_out0 = v$G27_12274_out0 && v$NQ2_3191_out0;
assign v$G26_4255_out0 = v$G27_12275_out0 && v$NQ2_3192_out0;
assign v$G15_4364_out0 = v$NQ0_16214_out0 && v$Q1_4619_out0;
assign v$G15_4365_out0 = v$NQ0_16215_out0 && v$Q1_4620_out0;
assign v$G11_5080_out0 = v$NQ2_3191_out0 && v$NQ1_263_out0;
assign v$G11_5081_out0 = v$NQ2_3192_out0 && v$NQ1_264_out0;
assign v$_5360_out0 = v$_2539_out1[1:0];
assign v$_5360_out1 = v$_2539_out1[3:2];
assign v$_5361_out0 = v$_2540_out1[1:0];
assign v$_5361_out1 = v$_2540_out1[3:2];
assign v$EQ13_5469_out0 = v$SEL12_13371_out0 == 4'h1;
assign v$EQ13_5470_out0 = v$SEL12_13372_out0 == 4'h1;
assign v$_6352_out0 = v$Mode_11483_out0[0:0];
assign v$_6352_out1 = v$Mode_11483_out0[2:2];
assign v$_6353_out0 = v$Mode_11484_out0[0:0];
assign v$_6353_out1 = v$Mode_11484_out0[2:2];
assign v$Q_6418_out0 = v$_10703_out0;
assign v$Q_6419_out0 = v$_10704_out0;
assign v$IR2$REG$IMMEDIATE_6456_out0 = v$SEL10_7597_out0;
assign v$IR2$REG$IMMEDIATE_6457_out0 = v$SEL10_7598_out0;
assign v$G16_6650_out0 = v$NQ3_1645_out0 && v$Q2_5696_out0;
assign v$G16_6651_out0 = v$NQ3_1646_out0 && v$Q2_5697_out0;
assign v$_7687_out0 = v$_3104_out0[1:0];
assign v$_7687_out1 = v$_3104_out0[3:2];
assign v$_7688_out0 = v$_3105_out0[1:0];
assign v$_7688_out1 = v$_3105_out0[3:2];
assign v$G29_7784_out0 = v$NQ1_263_out0 || v$NQ0_8120_out0;
assign v$G29_7785_out0 = v$NQ1_264_out0 || v$NQ0_8121_out0;
assign v$IR2$FPU$OP_7868_out0 = v$SEL13_5054_out0;
assign v$IR2$FPU$OP_7869_out0 = v$SEL13_5055_out0;
assign v$_8517_out0 = v$_8712_out0[1:0];
assign v$_8517_out1 = v$_8712_out0[3:2];
assign v$_8518_out0 = v$_8713_out0[1:0];
assign v$_8518_out1 = v$_8713_out0[3:2];
assign v$G11_8539_out0 = v$NQ1_17350_out0 && v$NQ0_15970_out0;
assign v$G11_8540_out0 = v$NQ1_17351_out0 && v$NQ0_15971_out0;
assign v$F3_8557_out0 = v$_3322_out1;
assign v$F3_8558_out0 = v$_3323_out1;
assign v$CINA_8774_out0 = v$CIN_16717_out0;
assign v$CINA_8856_out0 = v$CIN_16719_out0;
assign v$CINA_8897_out0 = v$CIN_16720_out0;
assign v$CINA_8979_out0 = v$CIN_16722_out0;
assign v$G66_9263_out0 = v$PCHALT_17182_out0 && v$G65_9154_out0;
assign v$G32_9441_out0 = v$NQ1_11550_out0 || v$NQ0_16214_out0;
assign v$G32_9442_out0 = v$NQ1_11551_out0 || v$NQ0_16215_out0;
assign v$_9795_out0 = v$_3104_out1[1:0];
assign v$_9795_out1 = v$_3104_out1[3:2];
assign v$_9796_out0 = v$_3105_out1[1:0];
assign v$_9796_out1 = v$_3105_out1[3:2];
assign v$G42_9958_out0 = v$Q2_18125_out0 && v$NQ3_3209_out0;
assign v$G42_9959_out0 = v$Q2_18126_out0 && v$NQ3_3210_out0;
assign v$MUX1_10337_out0 = v$CLEAR_19011_out0 ? v$C3_13741_out0 : v$A1_4168_out0;
assign v$MUX1_10338_out0 = v$CLEAR_19012_out0 ? v$C3_13742_out0 : v$A1_4169_out0;
assign v$_10356_out0 = v$_1369_out1[2:0];
assign v$_10356_out1 = v$_1369_out1[5:3];
assign v$_10359_out0 = v$_1372_out1[2:0];
assign v$_10359_out1 = v$_1372_out1[5:3];
assign v$IS$IR2$DATA$PROCESSING_10368_out0 = v$SEL4_7339_out0;
assign v$IS$IR2$DATA$PROCESSING_10369_out0 = v$SEL4_7340_out0;
assign v$G49_10904_out0 = v$NQ3_1645_out0 && v$Q1_11427_out0;
assign v$G49_10905_out0 = v$NQ3_1646_out0 && v$Q1_11428_out0;
assign v$G5_11186_out0 = v$NQ2_17316_out0 && v$G6_3580_out0;
assign v$G5_11187_out0 = v$NQ2_17317_out0 && v$G6_3581_out0;
assign v$G36_11364_out0 = v$NQ2_3191_out0 && v$Q3_18893_out0;
assign v$G36_11365_out0 = v$NQ2_3192_out0 && v$Q3_18894_out0;
assign v$G17_12250_out0 = v$NQ2_3191_out0 && v$Q1_11427_out0;
assign v$G17_12251_out0 = v$NQ2_3192_out0 && v$Q1_11428_out0;
assign v$F2_12662_out0 = v$_3322_out0;
assign v$F2_12663_out0 = v$_3323_out0;
assign v$DATA$OUT0_12867_out0 = v$RAMDOUT0_9426_out0;
assign v$Q_13552_out0 = v$_9265_out0;
assign v$Q_13553_out0 = v$_9266_out0;
assign v$_13561_out0 = v$_1677_out1[2:0];
assign v$_13561_out1 = v$_1677_out1[5:3];
assign v$_13564_out0 = v$_1680_out1[2:0];
assign v$_13564_out1 = v$_1680_out1[5:3];
assign v$G50_13791_out0 = v$NQ3_1645_out0 && v$Q2_5696_out0;
assign v$G50_13792_out0 = v$NQ3_1646_out0 && v$Q2_5697_out0;
assign v$_13867_out0 = v$_6707_out0[1:0];
assign v$_13867_out1 = v$_6707_out0[3:2];
assign v$_13868_out0 = v$_6708_out0[1:0];
assign v$_13868_out1 = v$_6708_out0[3:2];
assign v$_13873_out0 = v$Mode_13777_out0[0:0];
assign v$_13873_out1 = v$Mode_13777_out0[2:2];
assign v$_13874_out0 = v$Mode_13778_out0[0:0];
assign v$_13874_out1 = v$Mode_13778_out0[2:2];
assign v$G9_14031_out0 = v$NQ2_19175_out0 && v$NQ1_11550_out0;
assign v$G9_14032_out0 = v$NQ2_19176_out0 && v$NQ1_11551_out0;
assign v$MUX6_14134_out0 = v$PIPELINE$RESTART_19235_out0 ? v$C2_14082_out0 : v$FF9_11158_out0;
assign v$MUX6_14135_out0 = v$PIPELINE$RESTART_19236_out0 ? v$C2_14083_out0 : v$FF9_11159_out0;
assign v$POut_14269_out0 = v$_16264_out0;
assign v$POut_14270_out0 = v$_16265_out0;
assign v$_14324_out0 = v$_1677_out0[2:0];
assign v$_14324_out1 = v$_1677_out0[5:3];
assign v$_14327_out0 = v$_1680_out0[2:0];
assign v$_14327_out1 = v$_1680_out0[5:3];
assign v$G68_15429_out0 = v$PCHALT_17182_out0 && v$G67_14340_out0;
assign v$INSTR$READ_15505_out0 = v$INSTR$READ_7535_out0;
assign v$INSTR$READ_15506_out0 = v$INSTR$READ_7536_out0;
assign v$G62_15602_out0 = v$Q3_19033_out0 && v$NQ2_19175_out0;
assign v$G62_15603_out0 = v$Q3_19034_out0 && v$NQ2_19176_out0;
assign v$R1_15628_out0 = v$_7264_out1;
assign v$R1_15629_out0 = v$_7265_out1;
assign v$R0_15792_out0 = v$_7264_out0;
assign v$R0_15793_out0 = v$_7265_out0;
assign v$R3_15899_out0 = v$_3864_out1;
assign v$R3_15900_out0 = v$_3865_out1;
assign v$DATA$OUT1_16195_out0 = v$RAMDOUT1_8627_out0;
assign v$F0_16438_out0 = v$_5293_out0;
assign v$F0_16439_out0 = v$_5294_out0;
assign v$G3_16702_out0 = ! v$PHALT_18124_out0;
assign v$IR2$RD_16976_out0 = v$SEL5_704_out0;
assign v$IR2$RD_16977_out0 = v$SEL5_705_out0;
assign v$_16985_out0 = v$_10354_out0[11:0];
assign v$_16985_out1 = v$_10354_out0[27:16];
assign v$_16986_out0 = v$_10355_out0[11:0];
assign v$_16986_out1 = v$_10355_out0[27:16];
assign v$G50_17963_out0 = v$Q2_18125_out0 && v$NQ3_3209_out0;
assign v$G50_17964_out0 = v$Q2_18126_out0 && v$NQ3_3210_out0;
assign v$EQ1_18042_out0 = v$XOR1_4124_out0 == 5'h0;
assign v$EQ1_18043_out0 = v$XOR1_4125_out0 == 5'h0;
assign v$IR2$S$WB_18080_out0 = v$SEL11_8654_out0;
assign v$IR2$S$WB_18081_out0 = v$SEL11_8655_out0;
assign v$_18118_out0 = { v$G1_1343_out0,v$C2_18617_out0 };
assign v$_18119_out0 = { v$G1_1344_out0,v$C2_18618_out0 };
assign v$_18340_out0 = v$_1369_out0[2:0];
assign v$_18340_out1 = v$_1369_out0[5:3];
assign v$_18343_out0 = v$_1372_out0[2:0];
assign v$_18343_out1 = v$_1372_out0[5:3];
assign v$CLK4_18601_out0 = v$CLK4_7347_out0;
assign v$CLK4_18602_out0 = v$CLK4_7348_out0;
assign v$G68_18717_out0 = v$HALT$PREV$PREV_18681_out0 || v$G67_14719_out0;
assign v$G68_18718_out0 = v$HALT$PREV$PREV_18682_out0 || v$G67_14720_out0;
assign v$TX_18860_out0 = v$G4_14816_out0;
assign v$TX_18861_out0 = v$G4_14817_out0;
assign v$_18901_out0 = v$MODE_1773_out0[0:0];
assign v$_18901_out1 = v$MODE_1773_out0[2:2];
assign v$_18902_out0 = v$MODE_1774_out0[0:0];
assign v$_18902_out1 = v$MODE_1774_out0[2:2];
assign v$G14_19043_out0 = v$NQ0_15970_out0 && v$NQ2_17316_out0;
assign v$G14_19044_out0 = v$NQ0_15971_out0 && v$NQ2_17317_out0;
assign v$G42_19085_out0 = v$Q0_14284_out0 && v$NQ3_1645_out0;
assign v$G42_19086_out0 = v$Q0_14285_out0 && v$NQ3_1646_out0;
assign v$G60_19369_out0 = v$NQ3_3209_out0 && v$Q1_4619_out0;
assign v$G60_19370_out0 = v$NQ3_3210_out0 && v$Q1_4620_out0;
assign v$R_60_out0 = v$INSTR$READ_15505_out0;
assign v$R_61_out0 = v$INSTR$READ_15506_out0;
assign v$EQ7_239_out0 = v$Q_6418_out0 == 4'hc;
assign v$EQ7_240_out0 = v$Q_6419_out0 == 4'hc;
assign v$END_407_out0 = v$_13873_out1;
assign v$END_408_out0 = v$_13874_out1;
assign v$8_1341_out0 = v$IR2_4118_out0[11:10];
assign v$8_1342_out0 = v$IR2_4119_out0[11:10];
assign v$SEL12_1513_out0 = v$IR2_4118_out0[6:6];
assign v$SEL12_1514_out0 = v$IR2_4119_out0[6:6];
assign v$EQ6_1723_out0 = v$Q_6418_out0 == 4'hb;
assign v$EQ6_1724_out0 = v$Q_6419_out0 == 4'hb;
assign v$6_2112_out0 = v$IR2_4118_out0[15:15];
assign v$6_2113_out0 = v$IR2_4119_out0[15:15];
assign v$G48_2487_out0 = v$G51_3076_out0 && v$G54_2064_out0;
assign v$G48_2488_out0 = v$G51_3077_out0 && v$G54_2065_out0;
assign v$EQ3_2808_out0 = v$Q_6418_out0 == 4'hb;
assign v$EQ3_2809_out0 = v$Q_6419_out0 == 4'hb;
assign v$EQ4_2813_out0 = v$Q_13552_out0 == 4'h9;
assign v$EQ4_2814_out0 = v$Q_13553_out0 == 4'h9;
assign v$_3129_out0 = v$_14324_out0[0:0];
assign v$_3129_out1 = v$_14324_out0[2:2];
assign v$_3132_out0 = v$_14327_out0[0:0];
assign v$_3132_out1 = v$_14327_out0[2:2];
assign v$IR2_3511_out0 = v$IR2_4118_out0;
assign v$IR2_3512_out0 = v$IR2_4119_out0;
assign v$_3969_out0 = v$_7687_out0[0:0];
assign v$_3969_out1 = v$_7687_out0[1:1];
assign v$_3970_out0 = v$_7688_out0[0:0];
assign v$_3970_out1 = v$_7688_out0[1:1];
assign v$_4148_out0 = v$_6352_out1[0:0];
assign v$_4148_out1 = v$_6352_out1[1:1];
assign v$_4149_out0 = v$_6353_out1[0:0];
assign v$_4149_out1 = v$_6353_out1[1:1];
assign v$_4172_out0 = v$_8517_out0[0:0];
assign v$_4172_out1 = v$_8517_out0[1:1];
assign v$_4173_out0 = v$_8518_out0[0:0];
assign v$_4173_out1 = v$_8518_out0[1:1];
assign v$SEL10_4311_out0 = v$IR2_4118_out0[5:5];
assign v$SEL10_4312_out0 = v$IR2_4119_out0[5:5];
assign v$EQ3_4362_out0 = v$Q_13552_out0 == 4'hb;
assign v$EQ3_4363_out0 = v$Q_13553_out0 == 4'hb;
assign v$IR2$IS$LDST_4560_out0 = v$EQ12_1693_out0;
assign v$IR2$IS$LDST_4561_out0 = v$EQ12_1694_out0;
assign v$_4987_out0 = v$_218_out1[0:0];
assign v$_4987_out1 = v$_218_out1[1:1];
assign v$_4988_out0 = v$_219_out1[0:0];
assign v$_4988_out1 = v$_219_out1[1:1];
assign v$G47_5660_out0 = v$G49_10904_out0 || v$G50_13791_out0;
assign v$G47_5661_out0 = v$G49_10905_out0 || v$G50_13792_out0;
assign v$EQ14_5729_out0 = v$IR2$FPU$OP_7868_out0 == 2'h3;
assign v$EQ14_5730_out0 = v$IR2$FPU$OP_7869_out0 == 2'h3;
assign v$_6074_out0 = v$_218_out0[0:0];
assign v$_6074_out1 = v$_218_out0[1:1];
assign v$_6075_out0 = v$_219_out0[0:0];
assign v$_6075_out1 = v$_219_out0[1:1];
assign v$RX_6447_out0 = v$TX_18860_out0;
assign v$RX_6448_out0 = v$TX_18861_out0;
assign v$PIN_6871_out0 = v$_1829_out1;
assign v$PIN_6874_out0 = v$_1829_out0;
assign v$PIN_6877_out0 = v$_1830_out1;
assign v$PIN_6880_out0 = v$_1830_out0;
assign v$G58_7333_out0 = v$G60_19369_out0 || v$G59_4024_out0;
assign v$G58_7334_out0 = v$G60_19370_out0 || v$G59_4025_out0;
assign v$IR2$IS$FPU_7335_out0 = v$EQ13_5469_out0;
assign v$IR2$IS$FPU_7336_out0 = v$EQ13_5470_out0;
assign v$_7605_out0 = v$_13867_out1[0:0];
assign v$_7605_out1 = v$_13867_out1[1:1];
assign v$_7606_out0 = v$_13868_out1[0:0];
assign v$_7606_out1 = v$_13868_out1[1:1];
assign v$EQ1_7756_out0 = v$Q_6418_out0 == 4'h9;
assign v$EQ1_7757_out0 = v$Q_6419_out0 == 4'h9;
assign v$5_7828_out0 = v$IR2_4118_out0[1:0];
assign v$5_7829_out0 = v$IR2_4119_out0[1:0];
assign v$STP$SAVED_7884_out0 = v$MUX6_14134_out0;
assign v$STP$SAVED_7885_out0 = v$MUX6_14135_out0;
assign v$DATA$OUT_7936_out0 = v$DATA$OUT1_16195_out0;
assign v$DATA$OUT_7937_out0 = v$DATA$OUT0_12867_out0;
assign v$_8088_out0 = v$_18340_out0[0:0];
assign v$_8088_out1 = v$_18340_out0[2:2];
assign v$_8091_out0 = v$_18343_out0[0:0];
assign v$_8091_out1 = v$_18343_out0[2:2];
assign v$_8297_out0 = v$_2493_out1[0:0];
assign v$_8297_out1 = v$_2493_out1[1:1];
assign v$_8298_out0 = v$_2494_out1[0:0];
assign v$_8298_out1 = v$_2494_out1[1:1];
assign v$S_8341_out0 = v$S_1377_out0;
assign v$G61_8592_out0 = v$G62_15602_out0 && v$NQ1_11550_out0;
assign v$G61_8593_out0 = v$G62_15603_out0 && v$NQ1_11551_out0;
assign v$P_8621_out0 = v$_13873_out0;
assign v$P_8622_out0 = v$_13874_out0;
assign v$_9125_out0 = v$_1761_out0[0:0];
assign v$_9125_out1 = v$_1761_out0[1:1];
assign v$_9126_out0 = v$_1762_out0[0:0];
assign v$_9126_out1 = v$_1762_out0[1:1];
assign v$_9157_out0 = v$_5360_out1[0:0];
assign v$_9157_out1 = v$_5360_out1[1:1];
assign v$_9158_out0 = v$_5361_out1[0:0];
assign v$_9158_out1 = v$_5361_out1[1:1];
assign v$_9389_out0 = v$_10356_out1[0:0];
assign v$_9389_out1 = v$_10356_out1[2:2];
assign v$_9392_out0 = v$_10359_out1[0:0];
assign v$_9392_out1 = v$_10359_out1[2:2];
assign v$EQ5_9433_out0 = v$Q_6418_out0 == 4'ha;
assign v$EQ5_9434_out0 = v$Q_6419_out0 == 4'ha;
assign v$SEL4_9817_out0 = v$IR2_4118_out0[9:8];
assign v$SEL4_9818_out0 = v$IR2_4119_out0[9:8];
assign v$G60_9841_out0 = v$G61_17069_out0 && v$G68_18717_out0;
assign v$G60_9842_out0 = v$G61_17070_out0 && v$G68_18718_out0;
assign v$_9857_out0 = v$_9795_out0[0:0];
assign v$_9857_out1 = v$_9795_out0[1:1];
assign v$_9858_out0 = v$_9796_out0[0:0];
assign v$_9858_out1 = v$_9796_out0[1:1];
assign v$EQ4_10007_out0 = v$Q_6418_out0 == 4'hc;
assign v$EQ4_10008_out0 = v$Q_6419_out0 == 4'hc;
assign v$RXBYTE_10010_out0 = v$POut_14269_out0;
assign v$RXBYTE_10011_out0 = v$POut_14270_out0;
assign v$_11264_out0 = v$_13561_out1[0:0];
assign v$_11264_out1 = v$_13561_out1[2:2];
assign v$_11267_out0 = v$_13564_out1[0:0];
assign v$_11267_out1 = v$_13564_out1[2:2];
assign v$EQ2_12176_out0 = v$Q_13552_out0 == 4'ha;
assign v$EQ2_12177_out0 = v$Q_13553_out0 == 4'ha;
assign v$G28_12513_out0 = v$Q2_5696_out0 && v$G29_7784_out0;
assign v$G28_12514_out0 = v$Q2_5697_out0 && v$G29_7785_out0;
assign v$PARITY_12637_out0 = v$_18901_out0;
assign v$PARITY_12638_out0 = v$_18902_out0;
assign v$_12641_out0 = v$_8517_out1[0:0];
assign v$_12641_out1 = v$_8517_out1[1:1];
assign v$_12642_out0 = v$_8518_out1[0:0];
assign v$_12642_out1 = v$_8518_out1[1:1];
assign v$G35_13219_out0 = v$G36_11364_out0 && v$G37_748_out0;
assign v$G35_13220_out0 = v$G36_11365_out0 && v$G37_749_out0;
assign v$_13473_out0 = v$_16985_out0[3:0];
assign v$_13473_out1 = v$_16985_out0[11:8];
assign v$_13474_out0 = v$_16986_out0[3:0];
assign v$_13474_out1 = v$_16986_out0[11:8];
assign v$G40_14259_out0 = v$G41_19089_out0 && v$G42_9958_out0;
assign v$G40_14260_out0 = v$G41_19090_out0 && v$G42_9959_out0;
assign {v$A1_14282_out1,v$A1_14282_out0 } = v$REG1_14166_out0 + v$_18118_out0 + v$C1_6703_out0;
assign {v$A1_14283_out1,v$A1_14283_out0 } = v$REG1_14167_out0 + v$_18119_out0 + v$C1_6704_out0;
assign v$_14431_out0 = v$_7687_out1[0:0];
assign v$_14431_out1 = v$_7687_out1[1:1];
assign v$_14432_out0 = v$_7688_out1[0:0];
assign v$_14432_out1 = v$_7688_out1[1:1];
assign v$9_14775_out0 = v$IR2_4118_out0[14:12];
assign v$9_14776_out0 = v$IR2_4119_out0[14:12];
assign v$_14849_out0 = v$_1761_out1[0:0];
assign v$_14849_out1 = v$_1761_out1[1:1];
assign v$_14850_out0 = v$_1762_out1[0:0];
assign v$_14850_out1 = v$_1762_out1[1:1];
assign v$EQ1_14926_out0 = v$Q_13552_out0 == 4'h1;
assign v$EQ1_14927_out0 = v$Q_13553_out0 == 4'h1;
assign v$_15108_out0 = v$_2493_out0[0:0];
assign v$_15108_out1 = v$_2493_out0[1:1];
assign v$_15109_out0 = v$_2494_out0[0:0];
assign v$_15109_out1 = v$_2494_out0[1:1];
assign v$G2_15651_out0 = ! v$Write_3479_out0;
assign v$G2_15652_out0 = ! v$Write_3480_out0;
assign v$G2_15653_out0 = ! v$Write_3481_out0;
assign v$G2_15654_out0 = ! v$Write_3482_out0;
assign v$G2_15655_out0 = ! v$Write_3483_out0;
assign v$G2_15656_out0 = ! v$Write_3484_out0;
assign v$G2_15657_out0 = ! v$Write_3485_out0;
assign v$G2_15658_out0 = ! v$Write_3486_out0;
assign v$G2_15659_out0 = ! v$Write_3487_out0;
assign v$G2_15660_out0 = ! v$Write_3488_out0;
assign v$G2_15661_out0 = ! v$Write_3489_out0;
assign v$G2_15662_out0 = ! v$Write_3490_out0;
assign v$_15758_out0 = v$_10356_out0[0:0];
assign v$_15758_out1 = v$_10356_out0[2:2];
assign v$_15761_out0 = v$_10359_out0[0:0];
assign v$_15761_out1 = v$_10359_out0[2:2];
assign v$_15786_out0 = v$_13867_out0[0:0];
assign v$_15786_out1 = v$_13867_out0[1:1];
assign v$_15787_out0 = v$_13868_out0[0:0];
assign v$_15787_out1 = v$_13868_out0[1:1];
assign v$7_15947_out0 = v$IR2_4118_out0[8:8];
assign v$7_15948_out0 = v$IR2_4119_out0[8:8];
assign v$ParityEN_16385_out0 = v$_6352_out0;
assign v$ParityEN_16386_out0 = v$_6353_out0;
assign v$_16443_out0 = v$_9795_out1[0:0];
assign v$_16443_out1 = v$_9795_out1[1:1];
assign v$_16444_out0 = v$_9796_out1[0:0];
assign v$_16444_out1 = v$_9796_out1[1:1];
assign v$RXCLK_16448_out0 = v$RXCLK_1393_out0;
assign v$RXCLK_16449_out0 = v$RXCLK_1394_out0;
assign v$SEL11_16493_out0 = v$IR2_4118_out0[7:7];
assign v$SEL11_16494_out0 = v$IR2_4119_out0[7:7];
assign v$C_16498_out0 = v$C_3832_out0;
assign v$C_16499_out0 = v$C_3833_out0;
assign v$_16876_out0 = v$_18340_out1[0:0];
assign v$_16876_out1 = v$_18340_out1[2:2];
assign v$_16879_out0 = v$_18343_out1[0:0];
assign v$_16879_out1 = v$_18343_out1[2:2];
assign v$_17361_out0 = v$_14324_out1[0:0];
assign v$_17361_out1 = v$_14324_out1[2:2];
assign v$_17364_out0 = v$_14327_out1[0:0];
assign v$_17364_out1 = v$_14327_out1[2:2];
assign v$R_17367_out0 = v$G3_16702_out0;
assign v$_17381_out0 = v$_16985_out1[7:0];
assign v$_17381_out1 = v$_16985_out1[15:8];
assign v$_17382_out0 = v$_16986_out1[7:0];
assign v$_17382_out1 = v$_16986_out1[15:8];
assign v$G39_17501_out0 = v$Q2_5696_out0 && v$G42_19085_out0;
assign v$G39_17502_out0 = v$Q2_5697_out0 && v$G42_19086_out0;
assign v$_17577_out0 = v$_5360_out0[0:0];
assign v$_17577_out1 = v$_5360_out0[1:1];
assign v$_17578_out0 = v$_5361_out0[0:0];
assign v$_17578_out1 = v$_5361_out0[1:1];
assign v$G21_18276_out0 = v$G23_2483_out0 && v$G22_4474_out0;
assign v$G21_18277_out0 = v$G23_2484_out0 && v$G22_4475_out0;
assign v$_18599_out0 = v$_18901_out1[0:0];
assign v$_18599_out1 = v$_18901_out1[1:1];
assign v$_18600_out0 = v$_18902_out1[0:0];
assign v$_18600_out1 = v$_18902_out1[1:1];
assign v$_18787_out0 = v$_13561_out0[0:0];
assign v$_18787_out1 = v$_13561_out0[2:2];
assign v$_18790_out0 = v$_13564_out0[0:0];
assign v$_18790_out1 = v$_13564_out0[2:2];
assign v$MUX1_19207_out0 = v$EQ1_18042_out0 ? v$C4_15259_out0 : v$A1_3146_out0;
assign v$MUX1_19208_out0 = v$EQ1_18043_out0 ? v$C4_15260_out0 : v$A1_3147_out0;
assign v$G31_19245_out0 = v$G32_9441_out0 && v$NQ3_3209_out0;
assign v$G31_19246_out0 = v$G32_9442_out0 && v$NQ3_3210_out0;
assign v$EQ2_19266_out0 = v$Q_6418_out0 == 4'h0;
assign v$EQ2_19267_out0 = v$Q_6419_out0 == 4'h0;
assign v$G56_708_out0 = v$EQ3_2808_out0 || v$EQ4_10007_out0;
assign v$G56_709_out0 = v$EQ3_2809_out0 || v$EQ4_10008_out0;
assign v$IR2$S_1315_out0 = v$7_15947_out0;
assign v$IR2$S_1316_out0 = v$7_15948_out0;
assign v$G9_1331_out0 = ((v$_7605_out1 && !v$_14431_out1) || (!v$_7605_out1) && v$_14431_out1);
assign v$G9_1332_out0 = ((v$_7606_out1 && !v$_14432_out1) || (!v$_7606_out1) && v$_14432_out1);
assign v$DATA$OUT_1468_out0 = v$DATA$OUT_7936_out0;
assign v$DATA$OUT_1469_out0 = v$DATA$OUT_7937_out0;
assign v$G4_1491_out0 = ((v$_12641_out1 && !v$_8297_out1) || (!v$_12641_out1) && v$_8297_out1);
assign v$G4_1492_out0 = ((v$_12642_out1 && !v$_8298_out1) || (!v$_12642_out1) && v$_8298_out1);
assign v$G47_1685_out0 = v$PARITY_12637_out0 && v$EQ1_7756_out0;
assign v$G47_1686_out0 = v$PARITY_12638_out0 && v$EQ1_7757_out0;
assign v$R_1749_out0 = v$R_17367_out0;
assign v$_1827_out0 = { v$C8_7599_out0,v$_13473_out0 };
assign v$_1828_out0 = { v$C8_7600_out0,v$_13474_out0 };
assign v$IR2$FPU$OP_1845_out0 = v$SEL4_9817_out0;
assign v$IR2$FPU$OP_1846_out0 = v$SEL4_9818_out0;
assign v$G12_1981_out0 = ((v$_9125_out1 && !v$_9857_out1) || (!v$_9125_out1) && v$_9857_out1);
assign v$G12_1982_out0 = ((v$_9126_out1 && !v$_9858_out1) || (!v$_9126_out1) && v$_9858_out1);
assign v$G15_2030_out0 = ((v$_9125_out0 && !v$_9857_out0) || (!v$_9125_out0) && v$_9857_out0);
assign v$G15_2031_out0 = ((v$_9126_out0 && !v$_9858_out0) || (!v$_9126_out0) && v$_9858_out0);
assign v$B12_2114_out0 = v$_8088_out0;
assign v$B12_2117_out0 = v$_8091_out0;
assign v$G10_2161_out0 = ((v$_14849_out1 && !v$_16443_out1) || (!v$_14849_out1) && v$_16443_out1);
assign v$G10_2162_out0 = ((v$_14850_out1 && !v$_16444_out1) || (!v$_14850_out1) && v$_16444_out1);
assign v$G25_2658_out0 = v$IR2$IS$LDST_4560_out0 && v$IR2$S$WB_18080_out0;
assign v$G25_2659_out0 = v$IR2$IS$LDST_4561_out0 && v$IR2$S$WB_18081_out0;
assign v$G30_2660_out0 = v$G31_19245_out0 && v$Q2_18125_out0;
assign v$G30_2661_out0 = v$G31_19246_out0 && v$Q2_18126_out0;
assign v$B0_3421_out0 = v$_3129_out0;
assign v$B0_3424_out0 = v$_3132_out0;
assign v$2StopBits_3683_out0 = v$_4148_out1;
assign v$2StopBits_3684_out0 = v$_4149_out1;
assign v$G16_3720_out0 = ((v$_7605_out0 && !v$_14431_out0) || (!v$_7605_out0) && v$_14431_out0);
assign v$G16_3721_out0 = ((v$_7606_out0 && !v$_14432_out0) || (!v$_7606_out0) && v$_14432_out0);
assign v$S_4182_out0 = v$_18599_out1;
assign v$S_4183_out0 = v$_18600_out1;
assign v$B9_4220_out0 = v$_11264_out0;
assign v$B9_4223_out0 = v$_11267_out0;
assign v$IR2$FPU$LOAD_4390_out0 = v$SEL11_16493_out0;
assign v$IR2$FPU$LOAD_4391_out0 = v$SEL11_16494_out0;
assign v$G8_5032_out0 = ((v$_4987_out1 && !v$_9157_out1) || (!v$_4987_out1) && v$_9157_out1);
assign v$G8_5033_out0 = ((v$_4988_out1 && !v$_9158_out1) || (!v$_4988_out1) && v$_9158_out1);
assign v$_5212_out0 = v$IR2_3511_out0[14:12];
assign v$_5213_out0 = v$IR2_3512_out0[14:12];
assign v$OUT_5217_out0 = v$MUX1_19207_out0;
assign v$OUT_5218_out0 = v$MUX1_19208_out0;
assign v$G55_5265_out0 = v$G56_3361_out0 || v$G48_2487_out0;
assign v$G55_5266_out0 = v$G56_3362_out0 || v$G48_2488_out0;
assign v$G2_5670_out0 = ((v$_4172_out1 && !v$_15108_out1) || (!v$_4172_out1) && v$_15108_out1);
assign v$G2_5671_out0 = ((v$_4173_out1 && !v$_15109_out1) || (!v$_4173_out1) && v$_15109_out1);
assign v$G39_6326_out0 = v$G40_14259_out0 || v$G43_409_out0;
assign v$G39_6327_out0 = v$G40_14260_out0 || v$G43_410_out0;
assign v$G6_6428_out0 = ((v$_6074_out1 && !v$_17577_out1) || (!v$_6074_out1) && v$_17577_out1);
assign v$G6_6429_out0 = ((v$_6075_out1 && !v$_17578_out1) || (!v$_6075_out1) && v$_17578_out1);
assign v$PIN_6869_out0 = v$_17381_out1;
assign v$PIN_6870_out0 = v$_17381_out0;
assign v$PIN_6873_out0 = v$_13473_out1;
assign v$PIN_6875_out0 = v$_17382_out1;
assign v$PIN_6876_out0 = v$_17382_out0;
assign v$PIN_6879_out0 = v$_13474_out1;
assign v$_7176_out0 = v$_18787_out1[0:0];
assign v$_7176_out1 = v$_18787_out1[1:1];
assign v$_7179_out0 = v$_18790_out1[0:0];
assign v$_7179_out1 = v$_18790_out1[1:1];
assign v$_7258_out0 = v$_17361_out1[0:0];
assign v$_7258_out1 = v$_17361_out1[1:1];
assign v$_7261_out0 = v$_17364_out1[0:0];
assign v$_7261_out1 = v$_17364_out1[1:1];
assign v$_7272_out0 = v$IR2_3511_out0[7:4];
assign v$_7273_out0 = v$IR2_3512_out0[7:4];
assign v$_7591_out0 = v$IR2_3511_out0[4:0];
assign v$_7592_out0 = v$IR2_3512_out0[4:0];
assign v$IR2$15_7754_out0 = v$6_2112_out0;
assign v$IR2$15_7755_out0 = v$6_2113_out0;
assign v$IR2_8094_out0 = v$IR2_3511_out0;
assign v$IR2_8095_out0 = v$IR2_3512_out0;
assign v$G64_8104_out0 = v$EQ3_4362_out0 && v$G63_10444_out0;
assign v$G64_8105_out0 = v$EQ3_4363_out0 && v$G63_10445_out0;
assign v$G11_8572_out0 = ((v$_15786_out1 && !v$_3969_out1) || (!v$_15786_out1) && v$_3969_out1);
assign v$G11_8573_out0 = ((v$_15787_out1 && !v$_3970_out1) || (!v$_15787_out1) && v$_3970_out1);
assign v$CLK4_9180_out0 = v$RXCLK_16448_out0;
assign v$CLK4_9181_out0 = v$RXCLK_16449_out0;
assign v$RXBIT_9243_out0 = v$RX_6447_out0;
assign v$RXBIT_9244_out0 = v$RX_6448_out0;
assign v$G57_9305_out0 = v$EQ2_12176_out0 && v$G58_168_out0;
assign v$G57_9306_out0 = v$EQ2_12177_out0 && v$G58_169_out0;
assign v$_9753_out0 = v$_9389_out1[0:0];
assign v$_9753_out1 = v$_9389_out1[1:1];
assign v$_9756_out0 = v$_9392_out1[0:0];
assign v$_9756_out1 = v$_9392_out1[1:1];
assign v$B3_9845_out0 = v$_17361_out0;
assign v$B3_9848_out0 = v$_17364_out0;
assign v$_9873_out0 = v$_11264_out1[0:0];
assign v$_9873_out1 = v$_11264_out1[1:1];
assign v$_9876_out0 = v$_11267_out1[0:0];
assign v$_9876_out1 = v$_11267_out1[1:1];
assign v$B15_10446_out0 = v$_16876_out0;
assign v$B15_10449_out0 = v$_16879_out0;
assign v$G1_10773_out0 = ((v$_4172_out0 && !v$_15108_out0) || (!v$_4172_out0) && v$_15108_out0);
assign v$G1_10774_out0 = ((v$_4173_out0 && !v$_15109_out0) || (!v$_4173_out0) && v$_15109_out0);
assign v$OddParity_11182_out0 = v$_4148_out0;
assign v$OddParity_11183_out0 = v$_4149_out0;
assign v$B18_11368_out0 = v$_15758_out0;
assign v$B18_11371_out0 = v$_15761_out0;
assign v$Q1P_11515_out0 = v$G21_18276_out0;
assign v$Q1P_11516_out0 = v$G21_18277_out0;
assign v$_11531_out0 = v$_3129_out1[0:0];
assign v$_11531_out1 = v$_3129_out1[1:1];
assign v$_11534_out0 = v$_3132_out1[0:0];
assign v$_11534_out1 = v$_3132_out1[1:1];
assign v$_11920_out0 = v$IR2_3511_out0[9:9];
assign v$_11921_out0 = v$IR2_3512_out0[9:9];
assign v$G61_12174_out0 = v$EQ4_2813_out0 && v$P_8621_out0;
assign v$G61_12175_out0 = v$EQ4_2814_out0 && v$P_8622_out0;
assign v$IR2$FPU$32BIT_12372_out0 = v$SEL10_4311_out0;
assign v$IR2$FPU$32BIT_12373_out0 = v$SEL10_4312_out0;
assign v$G14_12611_out0 = ((v$_14849_out0 && !v$_16443_out0) || (!v$_14849_out0) && v$_16443_out0);
assign v$G14_12612_out0 = ((v$_14850_out0 && !v$_16444_out0) || (!v$_14850_out0) && v$_16444_out0);
assign v$G7_13231_out0 = ((v$_4987_out0 && !v$_9157_out0) || (!v$_4987_out0) && v$_9157_out0);
assign v$G7_13232_out0 = ((v$_4988_out0 && !v$_9158_out0) || (!v$_4988_out0) && v$_9158_out0);
assign v$G53_13284_out0 = v$EQ1_14926_out0 && v$G52_16544_out0;
assign v$G53_13285_out0 = v$EQ1_14927_out0 && v$G52_16545_out0;
assign v$_13433_out0 = v$PIN_6871_out0[3:0];
assign v$_13433_out1 = v$PIN_6871_out0[7:4];
assign v$_13436_out0 = v$PIN_6874_out0[3:0];
assign v$_13436_out1 = v$PIN_6874_out0[7:4];
assign v$_13439_out0 = v$PIN_6877_out0[3:0];
assign v$_13439_out1 = v$PIN_6877_out0[7:4];
assign v$_13442_out0 = v$PIN_6880_out0[3:0];
assign v$_13442_out1 = v$PIN_6880_out0[7:4];
assign v$IR2$M_13567_out0 = v$5_7828_out0;
assign v$IR2$M_13568_out0 = v$5_7829_out0;
assign v$_13758_out0 = v$_16876_out1[0:0];
assign v$_13758_out1 = v$_16876_out1[1:1];
assign v$_13761_out0 = v$_16879_out1[0:0];
assign v$_13761_out1 = v$_16879_out1[1:1];
assign v$B6_13883_out0 = v$_18787_out0;
assign v$B6_13886_out0 = v$_18790_out0;
assign v$G13_14029_out0 = ((v$_15786_out0 && !v$_3969_out0) || (!v$_15786_out0) && v$_3969_out0);
assign v$G13_14030_out0 = ((v$_15787_out0 && !v$_3970_out0) || (!v$_15787_out0) && v$_3970_out0);
assign v$G57_14037_out0 = v$G61_8592_out0 || v$G58_7333_out0;
assign v$G57_14038_out0 = v$G61_8593_out0 || v$G58_7334_out0;
assign v$G18_14086_out0 = ! v$C_16498_out0;
assign v$G18_14087_out0 = ! v$C_16499_out0;
assign v$IR2$D_15090_out0 = v$8_1341_out0;
assign v$IR2$D_15091_out0 = v$8_1342_out0;
assign v$G28_15272_out0 = v$IR2$IS$FPU_7335_out0 && v$EQ14_5729_out0;
assign v$G28_15273_out0 = v$IR2$IS$FPU_7336_out0 && v$EQ14_5730_out0;
assign v$G59_15731_out0 = v$G58_2714_out0 || v$G60_9841_out0;
assign v$G59_15732_out0 = v$G58_2715_out0 || v$G60_9842_out0;
assign v$G40_15739_out0 = v$Q1_11427_out0 && v$G39_17501_out0;
assign v$G40_15740_out0 = v$Q1_11428_out0 && v$G39_17502_out0;
assign v$G5_15815_out0 = ((v$_6074_out0 && !v$_17577_out0) || (!v$_6074_out0) && v$_17577_out0);
assign v$G5_15816_out0 = ((v$_6075_out0 && !v$_17578_out0) || (!v$_6075_out0) && v$_17578_out0);
assign v$IR2$FPU$LOADA_15851_out0 = v$SEL12_1513_out0;
assign v$IR2$FPU$LOADA_15852_out0 = v$SEL12_1514_out0;
assign v$G22_15929_out0 = ! v$C_16498_out0;
assign v$G22_15930_out0 = ! v$C_16499_out0;
assign v$G28_16226_out0 = v$STALL$PREV$CYCLE_6059_out0 || v$STP$SAVED_7884_out0;
assign v$G28_16227_out0 = v$STALL$PREV$CYCLE_6060_out0 || v$STP$SAVED_7885_out0;
assign v$END_16336_out0 = v$A1_14282_out1;
assign v$END_16337_out0 = v$A1_14283_out1;
assign v$ODDPARITY_16534_out0 = v$_18599_out0;
assign v$ODDPARITY_16535_out0 = v$_18600_out0;
assign v$_17208_out0 = v$_15758_out1[0:0];
assign v$_17208_out1 = v$_15758_out1[1:1];
assign v$_17211_out0 = v$_15761_out1[0:0];
assign v$_17211_out1 = v$_15761_out1[1:1];
assign v$SEL3_17270_out0 = v$IR2_3511_out0[15:12];
assign v$SEL3_17271_out0 = v$IR2_3512_out0[15:12];
assign v$_17358_out0 = v$IR2_3511_out0[3:2];
assign v$_17359_out0 = v$IR2_3512_out0[3:2];
assign v$G45_17511_out0 = ! v$P_8621_out0;
assign v$G45_17512_out0 = ! v$P_8622_out0;
assign v$_17965_out0 = v$_8088_out1[0:0];
assign v$_17965_out1 = v$_8088_out1[1:1];
assign v$_17968_out0 = v$_8091_out1[0:0];
assign v$_17968_out1 = v$_8091_out1[1:1];
assign v$G3_18094_out0 = ((v$_12641_out0 && !v$_8297_out0) || (!v$_12641_out0) && v$_8297_out0);
assign v$G3_18095_out0 = ((v$_12642_out0 && !v$_8298_out0) || (!v$_12642_out0) && v$_8298_out0);
assign v$_18623_out0 = v$IR2_3511_out0[8:8];
assign v$_18624_out0 = v$IR2_3512_out0[8:8];
assign v$IR2$OP_18625_out0 = v$9_14775_out0;
assign v$IR2$OP_18626_out0 = v$9_14776_out0;
assign v$B21_18689_out0 = v$_9389_out0;
assign v$B21_18692_out0 = v$_9392_out0;
assign v$G25_18703_out0 = v$G26_4254_out0 || v$G28_12513_out0;
assign v$G25_18704_out0 = v$G26_4255_out0 || v$G28_12514_out0;
assign v$R_18958_out0 = v$R_60_out0;
assign v$R_18959_out0 = v$R_61_out0;
assign v$G35_19105_out0 = ! v$IR2$IS$LDST_4560_out0;
assign v$G35_19106_out0 = ! v$IR2$IS$LDST_4561_out0;
assign v$G33_19227_out0 = v$IR2$IS$LDST_4560_out0 && v$IR2$S$WB_18080_out0;
assign v$G33_19228_out0 = v$IR2$IS$LDST_4561_out0 && v$IR2$S$WB_18081_out0;
assign v$EQ7_19241_out0 = v$IR2_3511_out0 == 16'h7000;
assign v$EQ7_19242_out0 = v$IR2_3512_out0 == 16'h7000;
assign v$G2_19310_out0 = v$RXENABLE_3897_out0 && v$RXCLK_16448_out0;
assign v$G2_19311_out0 = v$RXENABLE_3898_out0 && v$RXCLK_16449_out0;
assign v$RX_44_out0 = v$RXBIT_9243_out0;
assign v$RX_45_out0 = v$RXBIT_9244_out0;
assign v$G27_269_out0 = v$G1_10773_out0 || v$G2_5670_out0;
assign v$G27_270_out0 = v$G1_10774_out0 || v$G2_5671_out0;
assign v$K_313_out0 = v$_7591_out0;
assign v$K_314_out0 = v$_7592_out0;
assign v$G17_381_out0 = v$S_4182_out0 && v$NQ2_19175_out0;
assign v$G17_382_out0 = v$S_4183_out0 && v$NQ2_19176_out0;
assign v$B23_1441_out0 = v$_9753_out1;
assign v$B23_1444_out0 = v$_9756_out1;
assign v$G25_1470_out0 = v$G5_15815_out0 || v$G6_6428_out0;
assign v$G25_1471_out0 = v$G5_15816_out0 || v$G6_6429_out0;
assign v$OP_2034_out0 = v$IR2$OP_18625_out0;
assign v$OP_2035_out0 = v$IR2$OP_18626_out0;
assign v$B_2896_out0 = v$B6_13883_out0;
assign v$B_2897_out0 = v$B3_9845_out0;
assign v$B_2898_out0 = v$B21_18689_out0;
assign v$B_2899_out0 = v$B9_4220_out0;
assign v$B_2900_out0 = v$B15_10446_out0;
assign v$B_2904_out0 = v$B12_2114_out0;
assign v$B_2908_out0 = v$B0_3421_out0;
assign v$B_2913_out0 = v$B18_11368_out0;
assign v$B_2968_out0 = v$B6_13886_out0;
assign v$B_2969_out0 = v$B3_9848_out0;
assign v$B_2970_out0 = v$B21_18692_out0;
assign v$B_2971_out0 = v$B9_4223_out0;
assign v$B_2972_out0 = v$B15_10449_out0;
assign v$B_2976_out0 = v$B12_2117_out0;
assign v$B_2980_out0 = v$B0_3424_out0;
assign v$B_2985_out0 = v$B18_11371_out0;
assign v$RX_3176_out0 = v$RXBIT_9243_out0;
assign v$RX_3177_out0 = v$RXBIT_9244_out0;
assign v$G52_3181_out0 = v$S_4182_out0 || v$NQ0_16214_out0;
assign v$G52_3182_out0 = v$S_4183_out0 || v$NQ0_16215_out0;
assign v$B2_3326_out0 = v$_11531_out1;
assign v$B2_3329_out0 = v$_11534_out1;
assign v$C_3419_out0 = v$_11920_out0;
assign v$C_3420_out0 = v$_11921_out0;
assign v$G12_3804_out0 = ! v$IR2$FPU$LOADA_15851_out0;
assign v$G12_3805_out0 = ! v$IR2$FPU$LOADA_15852_out0;
assign v$B20_4112_out0 = v$_17208_out1;
assign v$B20_4115_out0 = v$_17211_out1;
assign v$B14_4158_out0 = v$_17965_out1;
assign v$B14_4161_out0 = v$_17968_out1;
assign v$IR1_4315_out0 = v$R_18958_out0;
assign v$IR1_4316_out0 = v$R_18959_out0;
assign v$IR2$VALID_4376_out0 = v$G59_15731_out0;
assign v$IR2$VALID_4377_out0 = v$G59_15732_out0;
assign v$RX_5021_out0 = v$RXBIT_9243_out0;
assign v$RX_5022_out0 = v$RXBIT_9244_out0;
assign v$G34_5096_out0 = v$G33_19227_out0 || v$G35_19105_out0;
assign v$G34_5097_out0 = v$G33_19228_out0 || v$G35_19106_out0;
assign v$LOADA_5363_out0 = v$IR2$FPU$LOADA_15851_out0;
assign v$LOADA_5364_out0 = v$IR2$FPU$LOADA_15852_out0;
assign v$S_6017_out0 = v$_18623_out0;
assign v$S_6018_out0 = v$_18624_out0;
assign v$G9_6588_out0 = ((v$G8_12863_out0 && !v$OddParity_11182_out0) || (!v$G8_12863_out0) && v$OddParity_11182_out0);
assign v$G9_6589_out0 = ((v$G8_12864_out0 && !v$OddParity_11183_out0) || (!v$G8_12864_out0) && v$OddParity_11183_out0);
assign v$PIN_6872_out0 = v$_1827_out0;
assign v$PIN_6878_out0 = v$_1828_out0;
assign v$NP_7574_out0 = v$G45_17511_out0;
assign v$NP_7575_out0 = v$G45_17512_out0;
assign v$EQ1_8110_out0 = v$OUT_5217_out0 == 5'h0;
assign v$EQ1_8111_out0 = v$OUT_5218_out0 == 5'h0;
assign v$OPCODE_8218_out0 = v$_5212_out0;
assign v$OPCODE_8219_out0 = v$_5213_out0;
assign v$SHIFT_8348_out0 = v$_17358_out0;
assign v$SHIFT_8349_out0 = v$_17359_out0;
assign v$B1_8426_out0 = v$_11531_out0;
assign v$B1_8429_out0 = v$_11534_out0;
assign v$_8760_out0 = v$_13433_out1[1:0];
assign v$_8760_out1 = v$_13433_out1[3:2];
assign v$_8763_out0 = v$_13436_out1[1:0];
assign v$_8763_out1 = v$_13436_out1[3:2];
assign v$_8766_out0 = v$_13439_out1[1:0];
assign v$_8766_out1 = v$_13439_out1[3:2];
assign v$_8769_out0 = v$_13442_out1[1:0];
assign v$_8769_out1 = v$_13442_out1[3:2];
assign v$B13_9022_out0 = v$_17965_out0;
assign v$B13_9025_out0 = v$_17968_out0;
assign v$G17_9176_out0 = v$G13_14029_out0 || v$G11_8572_out0;
assign v$G17_9177_out0 = v$G13_14030_out0 || v$G11_8573_out0;
assign v$RXFlagSet_9435_out0 = v$G53_13284_out0;
assign v$RXFlagSet_9436_out0 = v$G53_13285_out0;
assign v$B11_9443_out0 = v$_9873_out1;
assign v$B11_9446_out0 = v$_9876_out1;
assign v$G24_10000_out0 = v$NQ3_1645_out0 && v$G25_18703_out0;
assign v$G24_10001_out0 = v$NQ3_1646_out0 && v$G25_18704_out0;
assign v$EQ10_10285_out0 = v$IR2$FPU$OP_1845_out0 == 2'h3;
assign v$EQ10_10286_out0 = v$IR2$FPU$OP_1846_out0 == 2'h3;
assign v$B10_10297_out0 = v$_9873_out0;
assign v$B10_10300_out0 = v$_9876_out0;
assign v$G27_10687_out0 = v$S_4182_out0 && v$NQ2_19175_out0;
assign v$G27_10688_out0 = v$S_4183_out0 && v$NQ2_19176_out0;
assign v$G18_10707_out0 = v$G16_3720_out0 || v$G9_1331_out0;
assign v$G18_10708_out0 = v$G16_3721_out0 || v$G9_1332_out0;
assign v$G70_10735_out0 = v$S_4182_out0 && v$EQ6_1723_out0;
assign v$G70_10736_out0 = v$S_4183_out0 && v$EQ6_1724_out0;
assign v$G24_10805_out0 = v$G7_13231_out0 || v$G8_5032_out0;
assign v$G24_10806_out0 = v$G7_13232_out0 || v$G8_5033_out0;
assign v$IR15_11184_out0 = v$IR2$15_7754_out0;
assign v$IR15_11185_out0 = v$IR2$15_7755_out0;
assign v$B22_11300_out0 = v$_9753_out0;
assign v$B22_11303_out0 = v$_9756_out0;
assign v$G46_11405_out0 = ! v$S_4182_out0;
assign v$G46_11406_out0 = ! v$S_4183_out0;
assign v$LOAD_12270_out0 = v$IR2$FPU$LOAD_4390_out0;
assign v$LOAD_12271_out0 = v$IR2$FPU$LOAD_4391_out0;
assign v$IR2$FULL$OP$CODE_12392_out0 = v$SEL3_17270_out0;
assign v$IR2$FULL$OP$CODE_12393_out0 = v$SEL3_17271_out0;
assign v$CLK4_12779_out0 = v$G2_19310_out0;
assign v$CLK4_12780_out0 = v$G2_19311_out0;
assign v$G20_13310_out0 = v$G15_2030_out0 || v$G12_1981_out0;
assign v$G20_13311_out0 = v$G15_2031_out0 || v$G12_1982_out0;
assign v$SHIFTEN_13335_out0 = v$G57_14037_out0;
assign v$SHIFTEN_13336_out0 = v$G57_14038_out0;
assign v$_13413_out0 = v$_13433_out0[1:0];
assign v$_13413_out1 = v$_13433_out0[3:2];
assign v$_13416_out0 = v$_13436_out0[1:0];
assign v$_13416_out1 = v$_13436_out0[3:2];
assign v$_13419_out0 = v$_13439_out0[1:0];
assign v$_13419_out1 = v$_13439_out0[3:2];
assign v$_13422_out0 = v$_13442_out0[1:0];
assign v$_13422_out1 = v$_13442_out0[3:2];
assign v$_13431_out0 = v$PIN_6869_out0[3:0];
assign v$_13431_out1 = v$PIN_6869_out0[7:4];
assign v$_13432_out0 = v$PIN_6870_out0[3:0];
assign v$_13432_out1 = v$PIN_6870_out0[7:4];
assign v$_13435_out0 = v$PIN_6873_out0[3:0];
assign v$_13435_out1 = v$PIN_6873_out0[7:4];
assign v$_13437_out0 = v$PIN_6875_out0[3:0];
assign v$_13437_out1 = v$PIN_6875_out0[7:4];
assign v$_13438_out0 = v$PIN_6876_out0[3:0];
assign v$_13438_out1 = v$PIN_6876_out0[7:4];
assign v$_13441_out0 = v$PIN_6879_out0[3:0];
assign v$_13441_out1 = v$PIN_6879_out0[7:4];
assign v$B8_13715_out0 = v$_7176_out1;
assign v$B8_13718_out0 = v$_7179_out1;
assign v$B_13793_out0 = v$_7272_out0;
assign v$B_13794_out0 = v$_7273_out0;
assign v$G54_14798_out0 = v$G28_16226_out0 || v$HALT$PREV_10837_out0;
assign v$G54_14799_out0 = v$G28_16227_out0 || v$HALT$PREV_10838_out0;
assign v$G21_14847_out0 = v$G14_12611_out0 || v$G10_2161_out0;
assign v$G21_14848_out0 = v$G14_12612_out0 || v$G10_2162_out0;
assign v$B4_15266_out0 = v$_7258_out0;
assign v$B4_15269_out0 = v$_7261_out0;
assign v$G26_15513_out0 = v$G3_18094_out0 || v$G4_1491_out0;
assign v$G26_15514_out0 = v$G3_18095_out0 || v$G4_1492_out0;
assign v$G66_15853_out0 = ((v$ODDPARITY_16534_out0 && !v$EVENPARITY_14162_out0) || (!v$ODDPARITY_16534_out0) && v$EVENPARITY_14162_out0);
assign v$G66_15854_out0 = ((v$ODDPARITY_16535_out0 && !v$EVENPARITY_14163_out0) || (!v$ODDPARITY_16535_out0) && v$EVENPARITY_14163_out0);
assign v$B17_16125_out0 = v$_13758_out1;
assign v$B17_16128_out0 = v$_13761_out1;
assign v$G46_16729_out0 = v$G55_5265_out0 || v$G47_5660_out0;
assign v$G46_16730_out0 = v$G55_5266_out0 || v$G47_5661_out0;
assign v$ParityCheck_16733_out0 = v$G57_9305_out0;
assign v$ParityCheck_16734_out0 = v$G57_9306_out0;
assign v$G32_16952_out0 = v$G35_13219_out0 || v$G40_15739_out0;
assign v$G32_16953_out0 = v$G35_13220_out0 || v$G40_15740_out0;
assign v$B16_17034_out0 = v$_13758_out0;
assign v$B16_17037_out0 = v$_13761_out0;
assign v$RXReset_17150_out0 = v$G64_8104_out0;
assign v$RXReset_17151_out0 = v$G64_8105_out0;
assign v$G55_17278_out0 = v$EQ2_19266_out0 || v$G56_708_out0;
assign v$G55_17279_out0 = v$EQ2_19267_out0 || v$G56_709_out0;
assign v$RAMDOUT_17399_out0 = v$DATA$OUT_1468_out0;
assign v$RAMDOUT_17400_out0 = v$DATA$OUT_1469_out0;
assign v$B19_17410_out0 = v$_17208_out0;
assign v$B19_17413_out0 = v$_17211_out0;
assign v$G63_17433_out0 = v$G57_14037_out0 && v$SERIALIN_6011_out0;
assign v$G63_17434_out0 = v$G57_14038_out0 && v$SERIALIN_6012_out0;
assign v$B7_17634_out0 = v$_7176_out0;
assign v$B7_17637_out0 = v$_7179_out0;
assign v$MUX4_17682_out0 = v$G47_1685_out0 ? v$C4_3127_out0 : v$G39_6326_out0;
assign v$MUX4_17683_out0 = v$G47_1686_out0 ? v$C4_3128_out0 : v$G39_6327_out0;
assign v$G3_18299_out0 = ! v$R_1749_out0;
assign v$G9_18316_out0 = ! v$EQ7_19241_out0;
assign v$G9_18317_out0 = ! v$EQ7_19242_out0;
assign v$IR2_18567_out0 = v$IR2_8094_out0;
assign v$IR2_18568_out0 = v$IR2_8095_out0;
assign v$B5_18978_out0 = v$_7258_out1;
assign v$B5_18981_out0 = v$_7261_out1;
assign v$CHECKPARITY_1489_out0 = v$ParityCheck_16733_out0;
assign v$CHECKPARITY_1490_out0 = v$ParityCheck_16734_out0;
assign v$1_1687_out0 = v$IR2_18567_out0[8:8];
assign v$1_1688_out0 = v$IR2_18568_out0[8:8];
assign v$_1799_out0 = v$_13413_out1[0:0];
assign v$_1799_out1 = v$_13413_out1[1:1];
assign v$_1802_out0 = v$_13416_out1[0:0];
assign v$_1802_out1 = v$_13416_out1[1:1];
assign v$_1805_out0 = v$_13419_out1[0:0];
assign v$_1805_out1 = v$_13419_out1[1:1];
assign v$_1808_out0 = v$_13422_out1[0:0];
assign v$_1808_out1 = v$_13422_out1[1:1];
assign v$G65_2654_out0 = v$EQ5_9433_out0 && v$G66_15853_out0;
assign v$G65_2655_out0 = v$EQ5_9434_out0 && v$G66_15854_out0;
assign v$CLK4_2728_out0 = v$CLK4_12779_out0;
assign v$CLK4_2729_out0 = v$CLK4_12780_out0;
assign v$B_2901_out0 = v$B7_17634_out0;
assign v$B_2902_out0 = v$B1_8426_out0;
assign v$B_2903_out0 = v$B14_4158_out0;
assign v$B_2905_out0 = v$B8_13715_out0;
assign v$B_2906_out0 = v$B17_16125_out0;
assign v$B_2907_out0 = v$B23_1441_out0;
assign v$B_2909_out0 = v$B13_9022_out0;
assign v$B_2910_out0 = v$B4_15266_out0;
assign v$B_2911_out0 = v$B19_17410_out0;
assign v$B_2912_out0 = v$B22_11300_out0;
assign v$B_2914_out0 = v$B10_10297_out0;
assign v$B_2915_out0 = v$B20_4112_out0;
assign v$B_2916_out0 = v$B2_3326_out0;
assign v$B_2917_out0 = v$B11_9443_out0;
assign v$B_2918_out0 = v$B5_18978_out0;
assign v$B_2919_out0 = v$B16_17034_out0;
assign v$B_2973_out0 = v$B7_17637_out0;
assign v$B_2974_out0 = v$B1_8429_out0;
assign v$B_2975_out0 = v$B14_4161_out0;
assign v$B_2977_out0 = v$B8_13718_out0;
assign v$B_2978_out0 = v$B17_16128_out0;
assign v$B_2979_out0 = v$B23_1444_out0;
assign v$B_2981_out0 = v$B13_9025_out0;
assign v$B_2982_out0 = v$B4_15269_out0;
assign v$B_2983_out0 = v$B19_17413_out0;
assign v$B_2984_out0 = v$B22_11303_out0;
assign v$B_2986_out0 = v$B10_10300_out0;
assign v$B_2987_out0 = v$B20_4115_out0;
assign v$B_2988_out0 = v$B2_3329_out0;
assign v$B_2989_out0 = v$B11_9446_out0;
assign v$B_2990_out0 = v$B5_18981_out0;
assign v$B_2991_out0 = v$B16_17037_out0;
assign v$G10_3112_out0 = ((v$G9_6588_out0 && !v$RceivedParity_19151_out0) || (!v$G9_6588_out0) && v$RceivedParity_19151_out0);
assign v$G10_3113_out0 = ((v$G9_6589_out0 && !v$RceivedParity_19152_out0) || (!v$G9_6589_out0) && v$RceivedParity_19152_out0);
assign v$SEL6_3219_out0 = v$IR1_4315_out0[1:0];
assign v$SEL6_3220_out0 = v$IR1_4316_out0[1:0];
assign v$G11_3475_out0 = v$IR2$FPU$LOAD_4390_out0 && v$G12_3804_out0;
assign v$G11_3476_out0 = v$IR2$FPU$LOAD_4391_out0 && v$G12_3805_out0;
assign v$SEL2_3895_out0 = v$IR1_4315_out0[8:8];
assign v$SEL2_3896_out0 = v$IR1_4316_out0[8:8];
assign v$Q2P_4318_out0 = v$G24_10000_out0;
assign v$Q2P_4319_out0 = v$G24_10001_out0;
assign v$S_4400_out0 = v$S_6017_out0;
assign v$S_4401_out0 = v$S_6018_out0;
assign v$LOADA_5295_out0 = v$LOADA_5363_out0;
assign v$LOADA_5296_out0 = v$LOADA_5364_out0;
assign v$C_6338_out0 = v$C_3419_out0;
assign v$C_6339_out0 = v$C_3420_out0;
assign v$LOAD_6451_out0 = v$LOAD_12270_out0;
assign v$LOAD_6452_out0 = v$LOAD_12271_out0;
assign v$EQ6_6654_out0 = v$IR2$FULL$OP$CODE_12392_out0 == 4'h7;
assign v$EQ6_6655_out0 = v$IR2$FULL$OP$CODE_12393_out0 == 4'h7;
assign v$SHIFT_7303_out0 = v$SHIFT_8348_out0;
assign v$SHIFT_7304_out0 = v$SHIFT_8349_out0;
assign v$_7987_out0 = v$_13413_out0[0:0];
assign v$_7987_out1 = v$_13413_out0[1:1];
assign v$_7990_out0 = v$_13416_out0[0:0];
assign v$_7990_out1 = v$_13416_out0[1:1];
assign v$_7993_out0 = v$_13419_out0[0:0];
assign v$_7993_out1 = v$_13419_out0[1:1];
assign v$_7996_out0 = v$_13422_out0[0:0];
assign v$_7996_out1 = v$_13422_out0[1:1];
assign v$SEL9_8299_out0 = v$IR1_4315_out0[11:10];
assign v$SEL9_8300_out0 = v$IR1_4316_out0[11:10];
assign v$G54_8437_out0 = v$G55_17278_out0 || v$G63_17433_out0;
assign v$G54_8438_out0 = v$G55_17279_out0 || v$G63_17434_out0;
assign v$_8758_out0 = v$_13431_out1[1:0];
assign v$_8758_out1 = v$_13431_out1[3:2];
assign v$_8759_out0 = v$_13432_out1[1:0];
assign v$_8759_out1 = v$_13432_out1[3:2];
assign v$_8762_out0 = v$_13435_out1[1:0];
assign v$_8762_out1 = v$_13435_out1[3:2];
assign v$_8764_out0 = v$_13437_out1[1:0];
assign v$_8764_out1 = v$_13437_out1[3:2];
assign v$_8765_out0 = v$_13438_out1[1:0];
assign v$_8765_out1 = v$_13438_out1[3:2];
assign v$_8768_out0 = v$_13441_out1[1:0];
assign v$_8768_out1 = v$_13441_out1[3:2];
assign v$R_9127_out0 = v$RX_5021_out0;
assign v$R_9128_out0 = v$RX_5022_out0;
assign v$SEL1_9141_out0 = v$IR1_4315_out0[15:12];
assign v$SEL1_9142_out0 = v$IR1_4316_out0[15:12];
assign v$6_10287_out0 = v$IR2_18567_out0[7:7];
assign v$6_10288_out0 = v$IR2_18568_out0[7:7];
assign v$SHIFTEN_10737_out0 = v$SHIFTEN_13335_out0;
assign v$SHIFTEN_10738_out0 = v$SHIFTEN_13336_out0;
assign v$G28_11298_out0 = v$G27_269_out0 || v$G26_15513_out0;
assign v$G28_11299_out0 = v$G27_270_out0 || v$G26_15514_out0;
assign v$FINISHED_11360_out0 = v$EQ1_8110_out0;
assign v$FINISHED_11361_out0 = v$EQ1_8111_out0;
assign v$IR15_11494_out0 = v$IR15_11184_out0;
assign v$IR15_11495_out0 = v$IR15_11185_out0;
assign v$G18_11539_out0 = v$IR2$FPU$LOAD_4390_out0 && v$EQ10_10285_out0;
assign v$G18_11540_out0 = v$IR2$FPU$LOAD_4391_out0 && v$EQ10_10286_out0;
assign v$Q3P_12238_out0 = v$MUX4_17682_out0;
assign v$Q3P_12239_out0 = v$MUX4_17683_out0;
assign v$IR2$VALID_12366_out0 = v$IR2$VALID_4376_out0;
assign v$IR2$VALID_12367_out0 = v$IR2$VALID_4377_out0;
assign v$G11_12417_out0 = v$Q3_19033_out0 && v$G52_3181_out0;
assign v$G11_12418_out0 = v$Q3_19034_out0 && v$G52_3182_out0;
assign v$_12433_out0 = v$_8760_out1[0:0];
assign v$_12433_out1 = v$_8760_out1[1:1];
assign v$_12436_out0 = v$_8763_out1[0:0];
assign v$_12436_out1 = v$_8763_out1[1:1];
assign v$_12439_out0 = v$_8766_out1[0:0];
assign v$_12439_out1 = v$_8766_out1[1:1];
assign v$_12442_out0 = v$_8769_out1[0:0];
assign v$_12442_out1 = v$_8769_out1[1:1];
assign v$EQ11_12455_out0 = v$IR2$FULL$OP$CODE_12392_out0 == 4'h1;
assign v$EQ11_12456_out0 = v$IR2$FULL$OP$CODE_12393_out0 == 4'h1;
assign v$SEL11_12766_out0 = v$IR2_18567_out0[7:7];
assign v$SEL11_12767_out0 = v$IR2_18568_out0[7:7];
assign v$_12795_out0 = { v$K_313_out0,v$C1_16407_out0 };
assign v$_12796_out0 = { v$K_314_out0,v$C1_16408_out0 };
assign v$5_12857_out0 = v$IR2_18567_out0[9:9];
assign v$5_12858_out0 = v$IR2_18568_out0[9:9];
assign v$EQ4_13295_out0 = v$IR2_18567_out0 == 16'h7000;
assign v$EQ4_13296_out0 = v$IR2_18568_out0 == 16'h7000;
assign v$2_13308_out0 = v$IR2_18567_out0[11:10];
assign v$2_13309_out0 = v$IR2_18568_out0[11:10];
assign v$SEL10_13393_out0 = v$IR2_18567_out0[9:8];
assign v$SEL10_13394_out0 = v$IR2_18568_out0[9:8];
assign v$_13411_out0 = v$_13431_out0[1:0];
assign v$_13411_out1 = v$_13431_out0[3:2];
assign v$_13412_out0 = v$_13432_out0[1:0];
assign v$_13412_out1 = v$_13432_out0[3:2];
assign v$_13415_out0 = v$_13435_out0[1:0];
assign v$_13415_out1 = v$_13435_out0[3:2];
assign v$_13417_out0 = v$_13437_out0[1:0];
assign v$_13417_out1 = v$_13437_out0[3:2];
assign v$_13418_out0 = v$_13438_out0[1:0];
assign v$_13418_out1 = v$_13438_out0[3:2];
assign v$_13421_out0 = v$_13441_out0[1:0];
assign v$_13421_out1 = v$_13441_out0[3:2];
assign v$_13434_out0 = v$PIN_6872_out0[3:0];
assign v$_13434_out1 = v$PIN_6872_out0[7:4];
assign v$_13440_out0 = v$PIN_6878_out0[3:0];
assign v$_13440_out1 = v$PIN_6878_out0[7:4];
assign v$G1_13560_out0 = v$STATE_16630_out0 && v$G3_18299_out0;
assign v$EQ12_13843_out0 = v$IR2$FULL$OP$CODE_12392_out0 == 4'h1;
assign v$EQ12_13844_out0 = v$IR2$FULL$OP$CODE_12393_out0 == 4'h1;
assign v$3_13980_out0 = v$IR2_18567_out0[5:2];
assign v$3_13981_out0 = v$IR2_18568_out0[5:2];
assign v$Q3P_14397_out0 = v$G32_16952_out0;
assign v$Q3P_14398_out0 = v$G32_16953_out0;
assign v$G29_14601_out0 = v$G25_1470_out0 || v$G24_10805_out0;
assign v$G29_14602_out0 = v$G25_1471_out0 || v$G24_10806_out0;
assign v$7_14618_out0 = v$IR2_18567_out0[1:0];
assign v$7_14619_out0 = v$IR2_18568_out0[1:0];
assign v$9_14918_out0 = v$IR2_18567_out0[15:12];
assign v$9_14919_out0 = v$IR2_18568_out0[15:12];
assign v$G2_15098_out0 = ((v$RX_44_out0 && !v$FF3_7649_out0) || (!v$RX_44_out0) && v$FF3_7649_out0);
assign v$G2_15099_out0 = ((v$RX_45_out0 && !v$FF3_7650_out0) || (!v$RX_45_out0) && v$FF3_7650_out0);
assign v$_15112_out0 = v$_8760_out0[0:0];
assign v$_15112_out1 = v$_8760_out0[1:1];
assign v$_15115_out0 = v$_8763_out0[0:0];
assign v$_15115_out1 = v$_8763_out0[1:1];
assign v$_15118_out0 = v$_8766_out0[0:0];
assign v$_15118_out1 = v$_8766_out0[1:1];
assign v$_15121_out0 = v$_8769_out0[0:0];
assign v$_15121_out1 = v$_8769_out0[1:1];
assign v$B_15227_out0 = v$B_13793_out0;
assign v$B_15228_out0 = v$B_13794_out0;
assign v$RXSET_15291_out0 = v$RXFlagSet_9435_out0;
assign v$RXSET_15292_out0 = v$RXFlagSet_9436_out0;
assign v$RXINTERRUPT_15456_out0 = v$RXReset_17150_out0;
assign v$RXINTERRUPT_15457_out0 = v$RXReset_17151_out0;
assign v$SEL8_15723_out0 = v$IR1_4315_out0[9:8];
assign v$SEL8_15724_out0 = v$IR1_4316_out0[9:8];
assign v$4_15776_out0 = v$IR2_18567_out0[6:6];
assign v$4_15777_out0 = v$IR2_18568_out0[6:6];
assign v$MUX1_15845_out0 = v$G54_14798_out0 ? v$REG3_3046_out0 : v$R_18958_out0;
assign v$MUX1_15846_out0 = v$G54_14799_out0 ? v$REG3_3047_out0 : v$R_18959_out0;
assign v$8_16131_out0 = v$IR2_18567_out0[15:15];
assign v$8_16132_out0 = v$IR2_18568_out0[15:15];
assign v$SEL7_16208_out0 = v$IR1_4315_out0[9:9];
assign v$SEL7_16209_out0 = v$IR1_4316_out0[9:9];
assign v$G53_16434_out0 = v$G17_381_out0 || v$NQ3_3209_out0;
assign v$G53_16435_out0 = v$G17_382_out0 || v$NQ3_3210_out0;
assign v$G22_16456_out0 = v$G20_13310_out0 || v$G21_14847_out0;
assign v$G22_16457_out0 = v$G20_13311_out0 || v$G21_14848_out0;
assign v$G19_16556_out0 = v$G17_9176_out0 || v$G18_10707_out0;
assign v$G19_16557_out0 = v$G17_9177_out0 || v$G18_10708_out0;
assign v$G26_16639_out0 = v$NQ3_3209_out0 || v$G27_10687_out0;
assign v$G26_16640_out0 = v$NQ3_3210_out0 || v$G27_10688_out0;
assign v$EQ1_16735_out0 = v$OPCODE_8218_out0 == 3'h4;
assign v$EQ1_16736_out0 = v$OPCODE_8219_out0 == 3'h4;
assign v$ShiftOut_16960_out0 = v$G46_16729_out0;
assign v$ShiftOut_16961_out0 = v$G46_16730_out0;
assign v$OP_18253_out0 = v$OP_2034_out0;
assign v$OP_18254_out0 = v$OP_2035_out0;
assign v$G10_18785_out0 = v$NP_7574_out0 && v$G11_5080_out0;
assign v$G10_18786_out0 = v$NP_7575_out0 && v$G11_5081_out0;
assign v$NS_18801_out0 = v$G46_11405_out0;
assign v$NS_18802_out0 = v$G46_11406_out0;
assign v$EQ9_18887_out0 = v$IR2$FULL$OP$CODE_12392_out0 == 4'h1;
assign v$EQ9_18888_out0 = v$IR2$FULL$OP$CODE_12393_out0 == 4'h1;
assign v$EQ1_19203_out0 = v$IR2$FULL$OP$CODE_12392_out0 == 4'h1;
assign v$EQ1_19204_out0 = v$IR2$FULL$OP$CODE_12393_out0 == 4'h1;
assign v$IR1$S$WB_336_out0 = v$SEL2_3895_out0;
assign v$IR1$S$WB_337_out0 = v$SEL2_3896_out0;
assign v$RXSHIFT_736_out0 = v$ShiftOut_16960_out0;
assign v$RXSHIFT_737_out0 = v$ShiftOut_16961_out0;
assign v$G69_1355_out0 = ! v$R_9127_out0;
assign v$G69_1356_out0 = ! v$R_9128_out0;
assign v$R_1639_out0 = v$FINISHED_11360_out0;
assign v$R_1642_out0 = v$FINISHED_11361_out0;
assign v$_1797_out0 = v$_13411_out1[0:0];
assign v$_1797_out1 = v$_13411_out1[1:1];
assign v$_1798_out0 = v$_13412_out1[0:0];
assign v$_1798_out1 = v$_13412_out1[1:1];
assign v$_1801_out0 = v$_13415_out1[0:0];
assign v$_1801_out1 = v$_13415_out1[1:1];
assign v$_1803_out0 = v$_13417_out1[0:0];
assign v$_1803_out1 = v$_13417_out1[1:1];
assign v$_1804_out0 = v$_13418_out1[0:0];
assign v$_1804_out1 = v$_13418_out1[1:1];
assign v$_1807_out0 = v$_13421_out1[0:0];
assign v$_1807_out1 = v$_13421_out1[1:1];
assign v$EQ1_2712_out0 = v$OP_18253_out0 == 3'h4;
assign v$EQ1_2713_out0 = v$OP_18254_out0 == 3'h4;
assign v$IR2$OPCODE_2761_out0 = v$9_14918_out0;
assign v$IR2$OPCODE_2762_out0 = v$9_14919_out0;
assign v$MUX1_2778_out0 = v$G2_15653_out0 ? v$SIN_94_out0 : v$_7987_out0;
assign v$MUX1_2781_out0 = v$G2_15656_out0 ? v$SIN_97_out0 : v$_7990_out0;
assign v$MUX1_2784_out0 = v$G2_15659_out0 ? v$SIN_100_out0 : v$_7993_out0;
assign v$MUX1_2787_out0 = v$G2_15662_out0 ? v$SIN_103_out0 : v$_7996_out0;
assign v$_2849_out0 = v$OP_18253_out0[0:0];
assign v$_2850_out0 = v$OP_18254_out0[0:0];
assign v$IR2$FPU$OP_3088_out0 = v$SEL10_13393_out0;
assign v$IR2$FPU$OP_3089_out0 = v$SEL10_13394_out0;
assign v$IR2$IS$FPU_3137_out0 = v$EQ12_13843_out0;
assign v$IR2$IS$FPU_3138_out0 = v$EQ12_13844_out0;
assign v$_3193_out0 = v$OP_18253_out0[2:2];
assign v$_3194_out0 = v$OP_18254_out0[2:2];
assign v$IR2$N_3195_out0 = v$3_13980_out0;
assign v$IR2$N_3196_out0 = v$3_13981_out0;
assign v$MUX8_3794_out0 = v$G2_15653_out0 ? v$FF2_15392_out0 : v$_15112_out0;
assign v$MUX8_3797_out0 = v$G2_15656_out0 ? v$FF2_15395_out0 : v$_15115_out0;
assign v$MUX8_3800_out0 = v$G2_15659_out0 ? v$FF2_15398_out0 : v$_15118_out0;
assign v$MUX8_3803_out0 = v$G2_15662_out0 ? v$FF2_15401_out0 : v$_15121_out0;
assign v$B_3885_out0 = v$B_15227_out0;
assign v$B_3886_out0 = v$B_15228_out0;
assign v$G23_4550_out0 = v$G19_16556_out0 || v$G22_16456_out0;
assign v$G23_4551_out0 = v$G19_16557_out0 || v$G22_16457_out0;
assign v$IR2$D_5114_out0 = v$2_13308_out0;
assign v$IR2$D_5115_out0 = v$2_13309_out0;
assign v$RXset_5317_out0 = v$RXSET_15291_out0;
assign v$RXset_5318_out0 = v$RXSET_15292_out0;
assign v$MUX1_5354_out0 = v$FINISHED_11360_out0 ? v$C1_16272_out0 : v$OUT_5217_out0;
assign v$MUX1_5355_out0 = v$FINISHED_11361_out0 ? v$C1_16273_out0 : v$OUT_5218_out0;
assign v$EQ4_5656_out0 = v$SEL8_15723_out0 == 2'h2;
assign v$EQ4_5657_out0 = v$SEL8_15724_out0 == 2'h2;
assign v$IR1$RD_5731_out0 = v$SEL9_8299_out0;
assign v$IR1$RD_5732_out0 = v$SEL9_8300_out0;
assign v$IR2$U_6182_out0 = v$4_15776_out0;
assign v$IR2$U_6183_out0 = v$4_15777_out0;
assign v$G14_6392_out0 = v$G15_4364_out0 && v$G53_16434_out0;
assign v$G14_6393_out0 = v$G15_4365_out0 && v$G53_16435_out0;
assign v$ISMOV_6907_out0 = v$EQ1_16735_out0;
assign v$ISMOV_6908_out0 = v$EQ1_16736_out0;
assign v$FINISHED_7284_out0 = v$FINISHED_11360_out0;
assign v$FINISHED_7285_out0 = v$FINISHED_11361_out0;
assign v$SHIFTEN_7382_out0 = v$SHIFTEN_10737_out0;
assign v$SHIFTEN_7383_out0 = v$SHIFTEN_10738_out0;
assign v$G2_7905_out0 = v$G1_13560_out0 || v$S_8341_out0;
assign v$_7985_out0 = v$_13411_out0[0:0];
assign v$_7985_out1 = v$_13411_out0[1:1];
assign v$_7986_out0 = v$_13412_out0[0:0];
assign v$_7986_out1 = v$_13412_out0[1:1];
assign v$_7989_out0 = v$_13415_out0[0:0];
assign v$_7989_out1 = v$_13415_out0[1:1];
assign v$_7991_out0 = v$_13417_out0[0:0];
assign v$_7991_out1 = v$_13417_out0[1:1];
assign v$_7992_out0 = v$_13418_out0[0:0];
assign v$_7992_out1 = v$_13418_out0[1:1];
assign v$_7995_out0 = v$_13421_out0[0:0];
assign v$_7995_out1 = v$_13421_out0[1:1];
assign v$EQ2_8279_out0 = v$OP_18253_out0 == 3'h5;
assign v$EQ2_8280_out0 = v$OP_18254_out0 == 3'h5;
assign v$S_8475_out0 = v$S_4400_out0;
assign v$S_8476_out0 = v$S_4401_out0;
assign v$G69_8519_out0 = v$EQ7_239_out0 && v$NS_18801_out0;
assign v$G69_8520_out0 = v$EQ7_240_out0 && v$NS_18802_out0;
assign v$_8541_out0 = v$OP_18253_out0[1:1];
assign v$_8542_out0 = v$OP_18254_out0[1:1];
assign v$STOP$2_8543_out0 = v$EQ4_13295_out0;
assign v$STOP$2_8544_out0 = v$EQ4_13296_out0;
assign v$_8761_out0 = v$_13434_out1[1:0];
assign v$_8761_out1 = v$_13434_out1[3:2];
assign v$_8767_out0 = v$_13440_out1[1:0];
assign v$_8767_out1 = v$_13440_out1[3:2];
assign v$IR2$M_9178_out0 = v$7_14618_out0;
assign v$IR2$M_9179_out0 = v$7_14619_out0;
assign v$G8_9881_out0 = v$G9_14031_out0 && v$G11_12417_out0;
assign v$G8_9882_out0 = v$G9_14032_out0 && v$G11_12418_out0;
assign v$MUX5_9904_out0 = v$G2_15653_out0 ? v$FF5_1917_out0 : v$_7987_out1;
assign v$MUX5_9907_out0 = v$G2_15656_out0 ? v$FF5_1920_out0 : v$_7990_out1;
assign v$MUX5_9910_out0 = v$G2_15659_out0 ? v$FF5_1923_out0 : v$_7993_out1;
assign v$MUX5_9913_out0 = v$G2_15662_out0 ? v$FF5_1926_out0 : v$_7996_out1;
assign v$IR1$OPCODE_9944_out0 = v$SEL1_9141_out0;
assign v$IR1$OPCODE_9945_out0 = v$SEL1_9142_out0;
assign v$_9960_out0 = v$OP_18253_out0[2:2];
assign v$_9961_out0 = v$OP_18254_out0[2:2];
assign v$C_9990_out0 = v$C_6338_out0;
assign v$C_9991_out0 = v$C_6339_out0;
assign v$MUX3_10376_out0 = v$G2_15653_out0 ? v$FF7_8611_out0 : v$_15112_out1;
assign v$MUX3_10379_out0 = v$G2_15656_out0 ? v$FF7_8614_out0 : v$_15115_out1;
assign v$MUX3_10382_out0 = v$G2_15659_out0 ? v$FF7_8617_out0 : v$_15118_out1;
assign v$MUX3_10385_out0 = v$G2_15662_out0 ? v$FF7_8620_out0 : v$_15121_out1;
assign v$IR1$C$L_10480_out0 = v$SEL7_16208_out0;
assign v$IR1$C$L_10481_out0 = v$SEL7_16209_out0;
assign v$G10_10725_out0 = v$EQ6_6654_out0 && v$G9_18316_out0;
assign v$G10_10726_out0 = v$EQ6_6655_out0 && v$G9_18317_out0;
assign v$_10733_out0 = v$OP_18253_out0[1:1];
assign v$_10734_out0 = v$OP_18254_out0[1:1];
assign v$MUX6_10841_out0 = v$G2_15653_out0 ? v$FF1_16689_out0 : v$_1799_out1;
assign v$MUX6_10844_out0 = v$G2_15656_out0 ? v$FF1_16692_out0 : v$_1802_out1;
assign v$MUX6_10847_out0 = v$G2_15659_out0 ? v$FF1_16695_out0 : v$_1805_out1;
assign v$MUX6_10850_out0 = v$G2_15662_out0 ? v$FF1_16698_out0 : v$_1808_out1;
assign v$IR2$FPU$L_11232_out0 = v$SEL11_12766_out0;
assign v$IR2$FPU$L_11233_out0 = v$SEL11_12767_out0;
assign v$G62_12324_out0 = v$G61_12174_out0 && v$CLK4_2728_out0;
assign v$G62_12325_out0 = v$G61_12175_out0 && v$CLK4_2729_out0;
assign v$_12431_out0 = v$_8758_out1[0:0];
assign v$_12431_out1 = v$_8758_out1[1:1];
assign v$_12432_out0 = v$_8759_out1[0:0];
assign v$_12432_out1 = v$_8759_out1[1:1];
assign v$_12435_out0 = v$_8762_out1[0:0];
assign v$_12435_out1 = v$_8762_out1[1:1];
assign v$_12437_out0 = v$_8764_out1[0:0];
assign v$_12437_out1 = v$_8764_out1[1:1];
assign v$_12438_out0 = v$_8765_out1[0:0];
assign v$_12438_out1 = v$_8765_out1[1:1];
assign v$_12441_out0 = v$_8768_out1[0:0];
assign v$_12441_out1 = v$_8768_out1[1:1];
assign v$G1_12789_out0 = v$FINISHED_11360_out0 || v$CALCULATING_1647_out0;
assign v$G1_12790_out0 = v$FINISHED_11361_out0 || v$CALCULATING_1648_out0;
assign v$G20_12859_out0 = ! v$LOAD_6451_out0;
assign v$G20_12860_out0 = ! v$LOAD_6452_out0;
assign v$IR2$L_13058_out0 = v$5_12857_out0;
assign v$IR2$L_13059_out0 = v$5_12858_out0;
assign v$_13414_out0 = v$_13434_out0[1:0];
assign v$_13414_out1 = v$_13434_out0[3:2];
assign v$_13420_out0 = v$_13440_out0[1:0];
assign v$_13420_out1 = v$_13440_out0[3:2];
assign v$_13641_out0 = { v$Q2P_4318_out0,v$Q3P_14397_out0 };
assign v$_13642_out0 = { v$Q2P_4319_out0,v$Q3P_14398_out0 };
assign v$G11_13991_out0 = ! v$LOAD_6451_out0;
assign v$G11_13992_out0 = ! v$LOAD_6452_out0;
assign v$_14272_out0 = v$OP_18253_out0[0:0];
assign v$_14273_out0 = v$OP_18254_out0[0:0];
assign v$MUX2_14409_out0 = v$G2_15653_out0 ? v$FF8_15066_out0 : v$_12433_out1;
assign v$MUX2_14412_out0 = v$G2_15656_out0 ? v$FF8_15069_out0 : v$_12436_out1;
assign v$MUX2_14415_out0 = v$G2_15659_out0 ? v$FF8_15072_out0 : v$_12439_out1;
assign v$MUX2_14418_out0 = v$G2_15662_out0 ? v$FF8_15075_out0 : v$_12442_out1;
assign v$B$IS$RD_14695_out0 = v$G11_3475_out0;
assign v$B$IS$RD_14696_out0 = v$G11_3476_out0;
assign v$_15110_out0 = v$_8758_out0[0:0];
assign v$_15110_out1 = v$_8758_out0[1:1];
assign v$_15111_out0 = v$_8759_out0[0:0];
assign v$_15111_out1 = v$_8759_out0[1:1];
assign v$_15114_out0 = v$_8762_out0[0:0];
assign v$_15114_out1 = v$_8762_out0[1:1];
assign v$_15116_out0 = v$_8764_out0[0:0];
assign v$_15116_out1 = v$_8764_out0[1:1];
assign v$_15117_out0 = v$_8765_out0[0:0];
assign v$_15117_out1 = v$_8765_out0[1:1];
assign v$_15120_out0 = v$_8768_out0[0:0];
assign v$_15120_out1 = v$_8768_out0[1:1];
assign v$G10_15189_out0 = ! v$LOADA_5295_out0;
assign v$G10_15190_out0 = ! v$LOADA_5296_out0;
assign v$IR2$W_15717_out0 = v$1_1687_out0;
assign v$IR2$W_15718_out0 = v$1_1688_out0;
assign v$G64_15843_out0 = v$G54_8437_out0 || v$G65_2654_out0;
assign v$G64_15844_out0 = v$G54_8438_out0 || v$G65_2655_out0;
assign v$RXINTERRUPT_15935_out0 = v$RXINTERRUPT_15456_out0;
assign v$RXINTERRUPT_15936_out0 = v$RXINTERRUPT_15457_out0;
assign v$EQ3_16095_out0 = v$OP_18253_out0 == 3'h7;
assign v$EQ3_16096_out0 = v$OP_18254_out0 == 3'h7;
assign v$IR2$LS_16436_out0 = v$8_16131_out0;
assign v$IR2$LS_16437_out0 = v$8_16132_out0;
assign v$G19_16657_out0 = v$EQ9_18887_out0 && v$G18_11539_out0;
assign v$G19_16658_out0 = v$EQ9_18888_out0 && v$G18_11540_out0;
assign v$G12_16862_out0 = ! v$R_9127_out0;
assign v$G12_16863_out0 = ! v$R_9128_out0;
assign v$IR1_17302_out0 = v$MUX1_15845_out0;
assign v$IR1_17303_out0 = v$MUX1_15846_out0;
assign v$MUX4_17460_out0 = v$G2_15653_out0 ? v$FF6_2819_out0 : v$_12433_out0;
assign v$MUX4_17463_out0 = v$G2_15656_out0 ? v$FF6_2822_out0 : v$_12436_out0;
assign v$MUX4_17466_out0 = v$G2_15659_out0 ? v$FF6_2825_out0 : v$_12439_out0;
assign v$MUX4_17469_out0 = v$G2_15662_out0 ? v$FF6_2828_out0 : v$_12442_out0;
assign v$IR2$P_17955_out0 = v$6_10287_out0;
assign v$IR2$P_17956_out0 = v$6_10288_out0;
assign v$E_17993_out0 = v$G2_15098_out0;
assign v$E_17994_out0 = v$G2_15099_out0;
assign v$MUX7_18519_out0 = v$G2_15653_out0 ? v$FF3_10398_out0 : v$_1799_out0;
assign v$MUX7_18522_out0 = v$G2_15656_out0 ? v$FF3_10401_out0 : v$_1802_out0;
assign v$MUX7_18525_out0 = v$G2_15659_out0 ? v$FF3_10404_out0 : v$_1805_out0;
assign v$MUX7_18528_out0 = v$G2_15662_out0 ? v$FF3_10407_out0 : v$_1808_out0;
assign v$IR1$RM_18905_out0 = v$SEL6_3219_out0;
assign v$IR1$RM_18906_out0 = v$SEL6_3220_out0;
assign v$IR1$FPU$OP$CODE_18922_out0 = v$SEL8_15723_out0;
assign v$IR1$FPU$OP$CODE_18923_out0 = v$SEL8_15724_out0;
assign v$G24_18994_out0 = v$G25_14641_out0 && v$G26_16639_out0;
assign v$G24_18995_out0 = v$G25_14642_out0 && v$G26_16640_out0;
assign v$G37_19073_out0 = v$Q3_19033_out0 && v$NS_18801_out0;
assign v$G37_19074_out0 = v$Q3_19034_out0 && v$NS_18802_out0;
assign v$G30_19215_out0 = v$G28_11298_out0 || v$G29_14601_out0;
assign v$G30_19216_out0 = v$G28_11299_out0 || v$G29_14602_out0;
assign v$CheckParity_19290_out0 = v$CHECKPARITY_1489_out0;
assign v$CheckParity_19291_out0 = v$CHECKPARITY_1490_out0;
assign v$IR2$VALID_19367_out0 = v$IR2$VALID_12366_out0;
assign v$IR2$VALID_19368_out0 = v$IR2$VALID_12367_out0;
assign v$_316_out0 = v$IR1_17302_out0[15:12];
assign v$_317_out0 = v$IR1_17303_out0[15:12];
assign v$S_1004_out0 = v$S_8475_out0;
assign v$S_1005_out0 = v$S_8476_out0;
assign v$TX_1458_out0 = v$G64_15843_out0;
assign v$TX_1459_out0 = v$G64_15844_out0;
assign v$EQ16_1739_out0 = v$IR1$FPU$OP$CODE_18922_out0 == 2'h3;
assign v$EQ16_1740_out0 = v$IR1$FPU$OP$CODE_18923_out0 == 2'h3;
assign v$R_1743_out0 = v$R_1639_out0;
assign v$R_1746_out0 = v$R_1642_out0;
assign v$_1800_out0 = v$_13414_out1[0:0];
assign v$_1800_out1 = v$_13414_out1[1:1];
assign v$_1806_out0 = v$_13420_out1[0:0];
assign v$_1806_out1 = v$_13420_out1[1:1];
assign v$RXset_1859_out0 = v$RXset_5317_out0;
assign v$RXset_1860_out0 = v$RXset_5318_out0;
assign v$S_2636_out0 = v$S_8475_out0;
assign v$S_2637_out0 = v$S_8476_out0;
assign v$MUX1_2776_out0 = v$G2_15651_out0 ? v$SIN_92_out0 : v$_7985_out0;
assign v$MUX1_2777_out0 = v$G2_15652_out0 ? v$SIN_93_out0 : v$_7986_out0;
assign v$MUX1_2780_out0 = v$G2_15655_out0 ? v$SIN_96_out0 : v$_7989_out0;
assign v$MUX1_2782_out0 = v$G2_15657_out0 ? v$SIN_98_out0 : v$_7991_out0;
assign v$MUX1_2783_out0 = v$G2_15658_out0 ? v$SIN_99_out0 : v$_7992_out0;
assign v$MUX1_2786_out0 = v$G2_15661_out0 ? v$SIN_102_out0 : v$_7995_out0;
assign v$G6_3383_out0 = v$G8_9881_out0 || v$G14_6392_out0;
assign v$G6_3384_out0 = v$G8_9882_out0 || v$G14_6393_out0;
assign v$EQ7_3706_out0 = v$IR2$OPCODE_2761_out0 == 4'h1;
assign v$EQ7_3707_out0 = v$IR2$OPCODE_2762_out0 == 4'h1;
assign v$MUX8_3792_out0 = v$G2_15651_out0 ? v$FF2_15390_out0 : v$_15110_out0;
assign v$MUX8_3793_out0 = v$G2_15652_out0 ? v$FF2_15391_out0 : v$_15111_out0;
assign v$MUX8_3796_out0 = v$G2_15655_out0 ? v$FF2_15394_out0 : v$_15114_out0;
assign v$MUX8_3798_out0 = v$G2_15657_out0 ? v$FF2_15396_out0 : v$_15116_out0;
assign v$MUX8_3799_out0 = v$G2_15658_out0 ? v$FF2_15397_out0 : v$_15117_out0;
assign v$MUX8_3802_out0 = v$G2_15661_out0 ? v$FF2_15400_out0 : v$_15120_out0;
assign v$XOR3_4194_out0 = v$IR2$RD_16976_out0 ^ v$IR1$RM_18905_out0;
assign v$XOR3_4195_out0 = v$IR2$RD_16977_out0 ^ v$IR1$RM_18906_out0;
assign v$G20_5691_out0 = ! v$G19_16657_out0;
assign v$G20_5692_out0 = ! v$G19_16658_out0;
assign v$ShiftEN_6115_out0 = v$RXSHIFT_736_out0;
assign v$ShiftEN_6116_out0 = v$RXSHIFT_737_out0;
assign v$G6_6224_out0 = v$_9960_out0 && v$_8541_out0;
assign v$G6_6225_out0 = v$_9961_out0 && v$_8542_out0;
assign v$G9_6490_out0 = v$EQ2_8279_out0 || v$EQ3_16095_out0;
assign v$G9_6491_out0 = v$EQ2_8280_out0 || v$EQ3_16096_out0;
assign v$MUX2_6922_out0 = v$G47_1685_out0 ? v$C2_16851_out0 : v$G24_18994_out0;
assign v$MUX2_6923_out0 = v$G47_1686_out0 ? v$C2_16852_out0 : v$G24_18995_out0;
assign v$IR2$VALID_7739_out0 = v$IR2$VALID_19367_out0;
assign v$IR2$VALID_7740_out0 = v$IR2$VALID_19368_out0;
assign v$_7988_out0 = v$_13414_out0[0:0];
assign v$_7988_out1 = v$_13414_out0[1:1];
assign v$_7994_out0 = v$_13420_out0[0:0];
assign v$_7994_out1 = v$_13420_out0[1:1];
assign v$_8037_out0 = v$IR1_17302_out0[11:0];
assign v$_8038_out0 = v$IR1_17303_out0[11:0];
assign v$EQ9_8295_out0 = v$IR1_17302_out0 == 16'h7000;
assign v$EQ9_8296_out0 = v$IR1_17303_out0 == 16'h7000;
assign v$G19_8570_out0 = v$SHIFTEN_7382_out0 && v$CLK4_3873_out0;
assign v$G19_8571_out0 = v$SHIFTEN_7383_out0 && v$CLK4_3874_out0;
assign v$B_8628_out0 = v$B_3885_out0;
assign v$B_8629_out0 = v$B_3886_out0;
assign v$XOR1_8639_out0 = v$IR1$RM_18905_out0 ^ v$IR2$RD_16976_out0;
assign v$XOR1_8640_out0 = v$IR1$RM_18906_out0 ^ v$IR2$RD_16977_out0;
assign v$MUX1_8649_out0 = v$C_9990_out0 ? v$C1_14855_out0 : v$SHIFT_7303_out0;
assign v$MUX1_8650_out0 = v$C_9991_out0 ? v$C1_14856_out0 : v$SHIFT_7304_out0;
assign v$S_9799_out0 = v$S_8475_out0;
assign v$S_9800_out0 = v$S_8476_out0;
assign v$MUX5_9902_out0 = v$G2_15651_out0 ? v$FF5_1915_out0 : v$_7985_out1;
assign v$MUX5_9903_out0 = v$G2_15652_out0 ? v$FF5_1916_out0 : v$_7986_out1;
assign v$MUX5_9906_out0 = v$G2_15655_out0 ? v$FF5_1919_out0 : v$_7989_out1;
assign v$MUX5_9908_out0 = v$G2_15657_out0 ? v$FF5_1921_out0 : v$_7991_out1;
assign v$MUX5_9909_out0 = v$G2_15658_out0 ? v$FF5_1922_out0 : v$_7992_out1;
assign v$MUX5_9912_out0 = v$G2_15661_out0 ? v$FF5_1925_out0 : v$_7995_out1;
assign v$MUX3_10374_out0 = v$G2_15651_out0 ? v$FF7_8609_out0 : v$_15110_out1;
assign v$MUX3_10375_out0 = v$G2_15652_out0 ? v$FF7_8610_out0 : v$_15111_out1;
assign v$MUX3_10378_out0 = v$G2_15655_out0 ? v$FF7_8613_out0 : v$_15114_out1;
assign v$MUX3_10380_out0 = v$G2_15657_out0 ? v$FF7_8615_out0 : v$_15116_out1;
assign v$MUX3_10381_out0 = v$G2_15658_out0 ? v$FF7_8616_out0 : v$_15117_out1;
assign v$MUX3_10384_out0 = v$G2_15661_out0 ? v$FF7_8619_out0 : v$_15120_out1;
assign v$G3_10685_out0 = ! v$E_17993_out0;
assign v$G3_10686_out0 = ! v$E_17994_out0;
assign v$MUX6_10839_out0 = v$G2_15651_out0 ? v$FF1_16687_out0 : v$_1797_out1;
assign v$MUX6_10840_out0 = v$G2_15652_out0 ? v$FF1_16688_out0 : v$_1798_out1;
assign v$MUX6_10843_out0 = v$G2_15655_out0 ? v$FF1_16691_out0 : v$_1801_out1;
assign v$MUX6_10845_out0 = v$G2_15657_out0 ? v$FF1_16693_out0 : v$_1803_out1;
assign v$MUX6_10846_out0 = v$G2_15658_out0 ? v$FF1_16694_out0 : v$_1804_out1;
assign v$MUX6_10849_out0 = v$G2_15661_out0 ? v$FF1_16697_out0 : v$_1807_out1;
assign v$IR2$IS$FPU_12415_out0 = v$IR2$IS$FPU_3137_out0;
assign v$IR2$IS$FPU_12416_out0 = v$IR2$IS$FPU_3138_out0;
assign v$_12434_out0 = v$_8761_out1[0:0];
assign v$_12434_out1 = v$_8761_out1[1:1];
assign v$_12440_out0 = v$_8767_out1[0:0];
assign v$_12440_out1 = v$_8767_out1[1:1];
assign v$G32_12457_out0 = !(v$G30_19215_out0 || v$G23_4550_out0);
assign v$G32_12458_out0 = !(v$G30_19216_out0 || v$G23_4551_out0);
assign v$MUX5_12517_out0 = v$STP$SAVED_7884_out0 ? v$IR1_17302_out0 : v$R_18958_out0;
assign v$MUX5_12518_out0 = v$STP$SAVED_7885_out0 ? v$IR1_17303_out0 : v$R_18959_out0;
assign v$G4_12565_out0 = ! v$_3193_out0;
assign v$G4_12566_out0 = ! v$_3194_out0;
assign v$MUX2_12801_out0 = v$_10733_out0 ? v$FF1_10761_out0 : v$_14272_out0;
assign v$MUX2_12802_out0 = v$_10734_out0 ? v$FF1_10762_out0 : v$_14273_out0;
assign v$RXINT_13139_out0 = v$RXINTERRUPT_15935_out0;
assign v$RXINT_13140_out0 = v$RXINTERRUPT_15936_out0;
assign v$ISMOV_13213_out0 = v$ISMOV_6907_out0;
assign v$ISMOV_13214_out0 = v$ISMOV_6908_out0;
assign v$S_13389_out0 = v$S_8475_out0;
assign v$S_13390_out0 = v$S_8476_out0;
assign v$EQ2_13445_out0 = v$IR1$OPCODE_9944_out0 == 4'h1;
assign v$EQ2_13446_out0 = v$IR1$OPCODE_9945_out0 == 4'h1;
assign v$EQ1_13516_out0 = v$IR1$OPCODE_9944_out0 == 4'h0;
assign v$EQ1_13517_out0 = v$IR1$OPCODE_9945_out0 == 4'h0;
assign v$IR1_13974_out0 = v$IR1_17302_out0;
assign v$IR1_13975_out0 = v$IR1_17303_out0;
assign v$NEXTSTATE_14116_out0 = v$G2_7905_out0;
assign v$MUX2_14407_out0 = v$G2_15651_out0 ? v$FF8_15064_out0 : v$_12431_out1;
assign v$MUX2_14408_out0 = v$G2_15652_out0 ? v$FF8_15065_out0 : v$_12432_out1;
assign v$MUX2_14411_out0 = v$G2_15655_out0 ? v$FF8_15068_out0 : v$_12435_out1;
assign v$MUX2_14413_out0 = v$G2_15657_out0 ? v$FF8_15070_out0 : v$_12437_out1;
assign v$MUX2_14414_out0 = v$G2_15658_out0 ? v$FF8_15071_out0 : v$_12438_out1;
assign v$MUX2_14417_out0 = v$G2_15661_out0 ? v$FF8_15074_out0 : v$_12441_out1;
assign v$G36_14715_out0 = v$G37_19073_out0 && v$G38_10705_out0;
assign v$G36_14716_out0 = v$G37_19074_out0 && v$G38_10706_out0;
assign v$_15113_out0 = v$_8761_out0[0:0];
assign v$_15113_out1 = v$_8761_out0[1:1];
assign v$_15119_out0 = v$_8767_out0[0:0];
assign v$_15119_out1 = v$_8767_out0[1:1];
assign v$G68_15784_out0 = v$G69_8519_out0 || v$G70_10735_out0;
assign v$G68_15785_out0 = v$G69_8520_out0 || v$G70_10736_out0;
assign v$EQ6_16480_out0 = v$IR2$FPU$OP_3088_out0 == 2'h3;
assign v$EQ6_16481_out0 = v$IR2$FPU$OP_3089_out0 == 2'h3;
assign v$G9_16651_out0 = ! v$IR1$C$L_10480_out0;
assign v$G9_16652_out0 = ! v$IR1$C$L_10481_out0;
assign v$G10_17126_out0 = v$E_17993_out0 && v$NQ2_17316_out0;
assign v$G10_17127_out0 = v$E_17994_out0 && v$NQ2_17317_out0;
assign v$NR_17276_out0 = v$G12_16862_out0;
assign v$NR_17277_out0 = v$G12_16863_out0;
assign v$MUX4_17458_out0 = v$G2_15651_out0 ? v$FF6_2817_out0 : v$_12431_out0;
assign v$MUX4_17459_out0 = v$G2_15652_out0 ? v$FF6_2818_out0 : v$_12432_out0;
assign v$MUX4_17462_out0 = v$G2_15655_out0 ? v$FF6_2821_out0 : v$_12435_out0;
assign v$MUX4_17464_out0 = v$G2_15657_out0 ? v$FF6_2823_out0 : v$_12437_out0;
assign v$MUX4_17465_out0 = v$G2_15658_out0 ? v$FF6_2824_out0 : v$_12438_out0;
assign v$MUX4_17468_out0 = v$G2_15661_out0 ? v$FF6_2827_out0 : v$_12441_out0;
assign v$EQ15_17642_out0 = v$IR1$OPCODE_9944_out0 == 4'h1;
assign v$EQ15_17643_out0 = v$IR1$OPCODE_9945_out0 == 4'h1;
assign v$G2_18263_out0 = ! v$C_9990_out0;
assign v$G2_18264_out0 = ! v$C_9991_out0;
assign v$MUX1_18336_out0 = v$_2849_out0 ? v$C2_10434_out0 : v$C1_16938_out0;
assign v$MUX1_18337_out0 = v$_2850_out0 ? v$C2_10435_out0 : v$C1_16939_out0;
assign v$MUX7_18517_out0 = v$G2_15651_out0 ? v$FF3_10396_out0 : v$_1797_out0;
assign v$MUX7_18518_out0 = v$G2_15652_out0 ? v$FF3_10397_out0 : v$_1798_out0;
assign v$MUX7_18521_out0 = v$G2_15655_out0 ? v$FF3_10400_out0 : v$_1801_out0;
assign v$MUX7_18523_out0 = v$G2_15657_out0 ? v$FF3_10402_out0 : v$_1803_out0;
assign v$MUX7_18524_out0 = v$G2_15658_out0 ? v$FF3_10403_out0 : v$_1804_out0;
assign v$MUX7_18527_out0 = v$G2_15661_out0 ? v$FF3_10406_out0 : v$_1807_out0;
assign v$G11_18621_out0 = v$G10_3112_out0 && v$CheckParity_19290_out0;
assign v$G11_18622_out0 = v$G10_3113_out0 && v$CheckParity_19291_out0;
assign v$XOR2_19103_out0 = v$IR1$RD_5731_out0 ^ v$IR2$RD_16976_out0;
assign v$XOR2_19104_out0 = v$IR1$RD_5732_out0 ^ v$IR2$RD_16977_out0;
assign v$FINISHED_19280_out0 = v$FINISHED_7284_out0;
assign v$FINISHED_19281_out0 = v$FINISHED_7285_out0;
assign v$IR1_22_out0 = v$IR1_13974_out0;
assign v$IR1_23_out0 = v$IR1_13975_out0;
assign v$G29_744_out0 = ! v$EQ16_1739_out0;
assign v$G29_745_out0 = ! v$EQ16_1740_out0;
assign v$_996_out0 = v$B_8628_out0[2:2];
assign v$_997_out0 = v$B_8629_out0[2:2];
assign v$G34_1727_out0 = v$G35_4476_out0 || v$G36_14715_out0;
assign v$G34_1728_out0 = v$G35_4477_out0 || v$G36_14716_out0;
assign v$FINISHED_2461_out0 = v$FINISHED_19280_out0;
assign v$FINISHED_2462_out0 = v$FINISHED_19281_out0;
assign v$G8_2607_out0 = ! v$G9_6490_out0;
assign v$G8_2608_out0 = ! v$G9_6491_out0;
assign v$MUX1_2779_out0 = v$G2_15654_out0 ? v$SIN_95_out0 : v$_7988_out0;
assign v$MUX1_2785_out0 = v$G2_15660_out0 ? v$SIN_101_out0 : v$_7994_out0;
assign v$NE_3637_out0 = v$G3_10685_out0;
assign v$NE_3638_out0 = v$G3_10686_out0;
assign v$RXErrorSet_3679_out0 = v$G11_18621_out0;
assign v$RXErrorSet_3680_out0 = v$G11_18622_out0;
assign v$MUX8_3795_out0 = v$G2_15654_out0 ? v$FF2_15393_out0 : v$_15113_out0;
assign v$MUX8_3801_out0 = v$G2_15660_out0 ? v$FF2_15399_out0 : v$_15119_out0;
assign v$EQ6_4128_out0 = v$XOR2_19103_out0 == 2'h0;
assign v$EQ6_4129_out0 = v$XOR2_19104_out0 == 2'h0;
assign v$ISMOV_4234_out0 = v$ISMOV_13213_out0;
assign v$ISMOV_4235_out0 = v$ISMOV_13214_out0;
assign v$EQ5_5070_out0 = v$XOR3_4194_out0 == 2'h0;
assign v$EQ5_5071_out0 = v$XOR3_4195_out0 == 2'h0;
assign v$G1_5662_out0 = v$G10_17126_out0 && v$G11_8539_out0;
assign v$G1_5663_out0 = v$G10_17127_out0 && v$G11_8540_out0;
assign v$Q1P_6027_out0 = v$MUX2_6922_out0;
assign v$Q1P_6028_out0 = v$MUX2_6923_out0;
assign v$G21_7802_out0 = v$EQ6_16480_out0 && v$IR2$FPU$L_11232_out0;
assign v$G21_7803_out0 = v$EQ6_16481_out0 && v$IR2$FPU$L_11233_out0;
assign v$INTERRUPT1_8595_out0 = v$RXINT_13139_out0;
assign v$INTERRUPT1_8596_out0 = v$RXINT_13140_out0;
assign v$ISMOV_9117_out0 = v$ISMOV_13213_out0;
assign v$ISMOV_9118_out0 = v$ISMOV_13214_out0;
assign v$MUX5_9905_out0 = v$G2_15654_out0 ? v$FF5_1918_out0 : v$_7988_out1;
assign v$MUX5_9911_out0 = v$G2_15660_out0 ? v$FF5_1924_out0 : v$_7994_out1;
assign v$SR_10350_out0 = v$MUX1_8649_out0;
assign v$SR_10351_out0 = v$MUX1_8650_out0;
assign v$MUX3_10377_out0 = v$G2_15654_out0 ? v$FF7_8612_out0 : v$_15113_out1;
assign v$MUX3_10383_out0 = v$G2_15660_out0 ? v$FF7_8618_out0 : v$_15119_out1;
assign v$S_10809_out0 = v$S_13389_out0;
assign v$S_10810_out0 = v$S_13390_out0;
assign v$MUX6_10842_out0 = v$G2_15654_out0 ? v$FF1_16690_out0 : v$_1800_out1;
assign v$MUX6_10848_out0 = v$G2_15660_out0 ? v$FF1_16696_out0 : v$_1806_out1;
assign v$_11282_out0 = v$B_8628_out0[1:1];
assign v$_11283_out0 = v$B_8629_out0[1:1];
assign v$G67_11571_out0 = v$G71_15857_out0 && v$G68_15784_out0;
assign v$G67_11572_out0 = v$G71_15858_out0 && v$G68_15785_out0;
assign v$EQUAL_12184_out0 = v$G32_12457_out0;
assign v$EQUAL_12185_out0 = v$G32_12458_out0;
assign v$TX_12248_out0 = v$TX_1458_out0;
assign v$TX_12249_out0 = v$TX_1459_out0;
assign v$IR1$IS$LDST_13783_out0 = v$EQ1_13516_out0;
assign v$IR1$IS$LDST_13784_out0 = v$EQ1_13517_out0;
assign v$MUX2_14410_out0 = v$G2_15654_out0 ? v$FF8_15067_out0 : v$_12434_out1;
assign v$MUX2_14416_out0 = v$G2_15660_out0 ? v$FF8_15073_out0 : v$_12440_out1;
assign v$_14928_out0 = v$B_8628_out0[3:3];
assign v$_14929_out0 = v$B_8629_out0[3:3];
assign v$N_15106_out0 = v$_8037_out0;
assign v$N_15107_out0 = v$_8038_out0;
assign v$G10_15166_out0 = v$EQ2_13445_out0 && v$EQ4_5656_out0;
assign v$G10_15167_out0 = v$EQ2_13446_out0 && v$EQ4_5657_out0;
assign v$IR2$VALID_15430_out0 = v$IR2$VALID_7739_out0;
assign v$IR2$VALID_15431_out0 = v$IR2$VALID_7740_out0;
assign v$_15748_out0 = v$B_8628_out0[0:0];
assign v$_15749_out0 = v$B_8629_out0[0:0];
assign v$EQ3_15864_out0 = v$XOR1_8639_out0 == 2'h0;
assign v$EQ3_15865_out0 = v$XOR1_8640_out0 == 2'h0;
assign v$STP$DECODED_17154_out0 = v$EQ9_8295_out0;
assign v$STP$DECODED_17155_out0 = v$EQ9_8296_out0;
assign v$MUX4_17461_out0 = v$G2_15654_out0 ? v$FF6_2820_out0 : v$_12434_out0;
assign v$MUX4_17467_out0 = v$G2_15660_out0 ? v$FF6_2826_out0 : v$_12440_out0;
assign v$S_17544_out0 = v$RXset_1859_out0;
assign v$S_17555_out0 = v$RXset_1860_out0;
assign v$G16_17588_out0 = v$RXset_1859_out0 && v$RXlast_13391_out0;
assign v$G16_17589_out0 = v$RXset_1860_out0 && v$RXlast_13392_out0;
assign v$G9_17602_out0 = v$NQ2_3191_out0 && v$NR_17276_out0;
assign v$G9_17603_out0 = v$NQ2_3192_out0 && v$NR_17277_out0;
assign v$G3_18293_out0 = ! v$R_1743_out0;
assign v$G3_18296_out0 = ! v$R_1746_out0;
assign v$OP_18409_out0 = v$_316_out0;
assign v$OP_18410_out0 = v$_317_out0;
assign v$MUX7_18520_out0 = v$G2_15654_out0 ? v$FF3_10399_out0 : v$_1800_out0;
assign v$MUX7_18526_out0 = v$G2_15660_out0 ? v$FF3_10405_out0 : v$_1806_out0;
assign v$S_18561_out0 = v$S_9799_out0;
assign v$S_18562_out0 = v$S_9800_out0;
assign v$G20_18885_out0 = v$NR_17276_out0 || v$Q3_18893_out0;
assign v$G20_18886_out0 = v$NR_17277_out0 || v$Q3_18894_out0;
assign v$G1_19257_out0 = v$ShiftEN_6115_out0 && v$CLK4_9180_out0;
assign v$G1_19258_out0 = v$ShiftEN_6116_out0 && v$CLK4_9181_out0;
assign v$G1_166_out0 = v$S_2636_out0 && v$ISMOV_9117_out0;
assign v$G1_167_out0 = v$S_2637_out0 && v$ISMOV_9118_out0;
assign v$G1_1403_out0 = v$S_1004_out0 && v$ISMOV_4234_out0;
assign v$G1_1404_out0 = v$S_1005_out0 && v$ISMOV_4235_out0;
assign v$G30_1877_out0 = v$EQ15_17642_out0 && v$G29_744_out0;
assign v$G30_1878_out0 = v$EQ15_17643_out0 && v$G29_745_out0;
assign v$G2_2620_out0 = v$EQUAL_12184_out0 && v$G3_11496_out0;
assign v$G2_2621_out0 = v$EQUAL_12185_out0 && v$G3_11497_out0;
assign v$G15_2874_out0 = v$IR1$IS$LDST_13783_out0 && v$IR1$S$WB_336_out0;
assign v$G15_2875_out0 = v$IR1$IS$LDST_13784_out0 && v$IR1$S$WB_337_out0;
assign v$IS$IR1$FMUL_3174_out0 = v$G10_15166_out0;
assign v$IS$IR1$FMUL_3175_out0 = v$G10_15167_out0;
assign v$G24_3609_out0 = v$IR1$IS$LDST_13783_out0 && v$IR1$S$WB_336_out0;
assign v$G24_3610_out0 = v$IR1$IS$LDST_13784_out0 && v$IR1$S$WB_337_out0;
assign v$SR_4532_out0 = v$SR_10350_out0;
assign v$SR_4533_out0 = v$SR_10350_out0;
assign v$SR_4534_out0 = v$SR_10350_out0;
assign v$SR_4535_out0 = v$SR_10350_out0;
assign v$SR_4536_out0 = v$SR_10351_out0;
assign v$SR_4537_out0 = v$SR_10351_out0;
assign v$SR_4538_out0 = v$SR_10351_out0;
assign v$SR_4539_out0 = v$SR_10351_out0;
assign v$OP_5253_out0 = v$OP_18409_out0;
assign v$OP_5254_out0 = v$OP_18410_out0;
assign v$G33_5348_out0 = v$NQ2_19175_out0 && v$G34_1727_out0;
assign v$G33_5349_out0 = v$NQ2_19176_out0 && v$G34_1728_out0;
assign v$IR2$VALID_6701_out0 = v$IR2$VALID_15430_out0;
assign v$IR2$VALID_6702_out0 = v$IR2$VALID_15431_out0;
assign v$G1_7643_out0 = v$G2_18263_out0 && v$_15748_out0;
assign v$G1_7644_out0 = v$G2_18264_out0 && v$_15749_out0;
assign v$IR1_7941_out0 = v$IR1_22_out0;
assign v$IR1_7942_out0 = v$IR1_23_out0;
assign v$G18_8726_out0 = v$G20_18885_out0 && v$G19_2605_out0;
assign v$G18_8727_out0 = v$G20_18886_out0 && v$G19_2606_out0;
assign v$G11_9984_out0 = v$EQ6_4128_out0 || v$EQ5_5070_out0;
assign v$G11_9985_out0 = v$EQ6_4129_out0 || v$EQ5_5071_out0;
assign v$Shift_9986_out0 = v$G1_19257_out0;
assign v$Shift_9987_out0 = v$G1_19258_out0;
assign v$EXEC2_10281_out0 = v$IR2$VALID_15430_out0;
assign v$EXEC2_10282_out0 = v$IR2$VALID_15431_out0;
assign v$IR2$VALID_11160_out0 = v$IR2$VALID_15430_out0;
assign v$IR2$VALID_11161_out0 = v$IR2$VALID_15431_out0;
assign v$G8_11581_out0 = v$Q1_11427_out0 && v$G9_17602_out0;
assign v$G8_11582_out0 = v$Q1_11428_out0 && v$G9_17603_out0;
assign v$FINISHED_12202_out0 = v$FINISHED_2461_out0;
assign v$FINISHED_12203_out0 = v$FINISHED_2462_out0;
assign v$G13_12722_out0 = v$G14_19043_out0 && v$NE_3637_out0;
assign v$G13_12723_out0 = v$G14_19044_out0 && v$NE_3638_out0;
assign v$ERR_13343_out0 = v$RXErrorSet_3679_out0;
assign v$ERR_13344_out0 = v$RXErrorSet_3680_out0;
assign v$G1_13554_out0 = v$STATE_16624_out0 && v$G3_18293_out0;
assign v$G1_13557_out0 = v$STATE_16627_out0 && v$G3_18296_out0;
assign v$G15_14180_out0 = v$NE_3637_out0 && v$G16_3233_out0;
assign v$G15_14181_out0 = v$NE_3638_out0 && v$G16_3234_out0;
assign v$G32_14802_out0 = v$IR1$IS$LDST_13783_out0 && v$G34_5096_out0;
assign v$G32_14803_out0 = v$IR1$IS$LDST_13784_out0 && v$G34_5097_out0;
assign v$G25_15262_out0 = v$G21_7802_out0 && v$EQ7_3706_out0;
assign v$G25_15263_out0 = v$G21_7803_out0 && v$EQ7_3707_out0;
assign v$G4_15287_out0 = v$NE_3637_out0 && v$G5_11186_out0;
assign v$G4_15288_out0 = v$NE_3638_out0 && v$G5_11187_out0;
assign v$G17_15402_out0 = v$IR2$VALID_15430_out0 && v$G20_5691_out0;
assign v$G17_15403_out0 = v$IR2$VALID_15431_out0 && v$G20_5692_out0;
assign v$N_15454_out0 = v$N_15106_out0;
assign v$N_15455_out0 = v$N_15107_out0;
assign v$EQUAL_16432_out0 = v$EQUAL_12184_out0;
assign v$EQUAL_16433_out0 = v$EQUAL_12185_out0;
assign v$EXEC2_16486_out0 = v$IR2$VALID_15430_out0;
assign v$EXEC2_16487_out0 = v$IR2$VALID_15431_out0;
assign v$TXRST_16998_out0 = v$G67_11571_out0;
assign v$TXRST_16999_out0 = v$G67_11572_out0;
assign v$EN_17005_out0 = v$_11282_out0;
assign v$EN_17006_out0 = v$_996_out0;
assign v$EN_17007_out0 = v$_14928_out0;
assign v$EN_17009_out0 = v$_11283_out0;
assign v$EN_17010_out0 = v$_997_out0;
assign v$EN_17011_out0 = v$_14929_out0;
assign v$S_17546_out0 = v$G16_17588_out0;
assign v$S_17557_out0 = v$G16_17589_out0;
assign v$G14_17632_out0 = v$IR1$IS$LDST_13783_out0 && v$G9_16651_out0;
assign v$G14_17633_out0 = v$IR1$IS$LDST_13784_out0 && v$G9_16652_out0;
assign v$G36_17991_out0 = ! v$STP$DECODED_17154_out0;
assign v$G36_17992_out0 = ! v$STP$DECODED_17155_out0;
assign v$EDGE1_18050_out0 = v$INTERRUPT1_8595_out0;
assign v$EDGE1_18051_out0 = v$INTERRUPT1_8596_out0;
assign v$EXEC2_448_out0 = v$EXEC2_16486_out0;
assign v$EXEC2_449_out0 = v$EXEC2_16487_out0;
assign v$IR1$IS$FPU$ARITHMETIC_1533_out0 = v$G30_1877_out0;
assign v$IR1$IS$FPU$ARITHMETIC_1534_out0 = v$G30_1878_out0;
assign v$G1_2078_out0 = v$EXEC2_16486_out0 && v$IR15_11494_out0;
assign v$G1_2079_out0 = v$EXEC2_16487_out0 && v$IR15_11495_out0;
assign v$EXEC2_2109_out0 = v$EXEC2_10281_out0;
assign v$EXEC2_2110_out0 = v$EXEC2_10282_out0;
assign v$G12_2420_out0 = v$G13_12722_out0 || v$G15_14180_out0;
assign v$G12_2421_out0 = v$G13_12723_out0 || v$G15_14181_out0;
assign v$G3_2634_out0 = v$G15_2874_out0 && v$IS$IR2$DATA$PROCESSING_10368_out0;
assign v$G3_2635_out0 = v$G15_2875_out0 && v$IS$IR2$DATA$PROCESSING_10369_out0;
assign v$G29_3814_out0 = v$G30_2660_out0 || v$G33_5348_out0;
assign v$G29_3815_out0 = v$G30_2661_out0 || v$G33_5349_out0;
assign v$G3_4110_out0 = v$G8_11581_out0 || v$G10_18785_out0;
assign v$G3_4111_out0 = v$G8_11582_out0 || v$G10_18786_out0;
assign v$SEL1_5457_out0 = v$IR1_7941_out0[9:8];
assign v$SEL1_5458_out0 = v$IR1_7942_out0[9:8];
assign v$G12_6432_out0 = v$IS$IR1$FMUL_3174_out0 && v$G11_9984_out0;
assign v$G12_6433_out0 = v$IS$IR1$FMUL_3175_out0 && v$G11_9985_out0;
assign v$_6443_out0 = v$IR1_7941_out0[1:0];
assign v$_6444_out0 = v$IR1_7942_out0[1:0];
assign v$IR2$VALID$AND$NOT$FLOAD_7603_out0 = v$G17_15402_out0;
assign v$IR2$VALID$AND$NOT$FLOAD_7604_out0 = v$G17_15403_out0;
assign v$FINISHED_8327_out0 = v$FINISHED_12202_out0;
assign v$FINISHED_8328_out0 = v$FINISHED_12203_out0;
assign v$TXRST_8358_out0 = v$TXRST_16998_out0;
assign v$TXRST_8359_out0 = v$TXRST_16999_out0;
assign v$N_8578_out0 = v$N_15454_out0;
assign v$N_8579_out0 = v$N_15455_out0;
assign v$S_10894_out0 = v$G1_1403_out0;
assign v$S_10895_out0 = v$G1_1404_out0;
assign v$S_11196_out0 = v$G1_166_out0;
assign v$S_11197_out0 = v$G1_167_out0;
assign v$N_12539_out0 = v$N_15454_out0;
assign v$N_12540_out0 = v$N_15455_out0;
assign v$_13341_out0 = v$IR1_7941_out0[15:15];
assign v$_13342_out0 = v$IR1_7942_out0[15:15];
assign v$G26_13755_out0 = v$G24_3609_out0 && v$G25_2658_out0;
assign v$G26_13756_out0 = v$G24_3610_out0 && v$G25_2659_out0;
assign v$SEL13_13831_out0 = v$IR1_7941_out0[5:5];
assign v$SEL13_13832_out0 = v$IR1_7942_out0[5:5];
assign v$IR2$VALID_13833_out0 = v$IR2$VALID_6701_out0;
assign v$IR2$VALID_13834_out0 = v$IR2$VALID_6702_out0;
assign v$_14119_out0 = v$IR1_7941_out0[8:8];
assign v$_14120_out0 = v$IR1_7942_out0[8:8];
assign v$G23_14691_out0 = ! v$G25_15262_out0;
assign v$G23_14692_out0 = ! v$G25_15263_out0;
assign v$G37_14699_out0 = v$IS$IR1$FMUL_3174_out0 && v$IS$IR2$DATA$PROCESSING_10368_out0;
assign v$G37_14700_out0 = v$IS$IR1$FMUL_3175_out0 && v$IS$IR2$DATA$PROCESSING_10369_out0;
assign v$OP_15388_out0 = v$OP_5253_out0;
assign v$OP_15389_out0 = v$OP_5254_out0;
assign v$COUNTERINTERRUPT_15460_out0 = v$G2_2620_out0;
assign v$COUNTERINTERRUPT_15461_out0 = v$G2_2621_out0;
assign v$IR2$VALID_16482_out0 = v$IR2$VALID_11160_out0;
assign v$IR2$VALID_16483_out0 = v$IR2$VALID_11161_out0;
assign v$_16528_out0 = v$IR1_7941_out0[11:10];
assign v$_16529_out0 = v$IR1_7942_out0[11:10];
assign v$EN_17004_out0 = v$G1_7643_out0;
assign v$EN_17008_out0 = v$G1_7644_out0;
assign v$_17304_out0 = v$IR1_7941_out0[14:12];
assign v$_17305_out0 = v$IR1_7942_out0[14:12];
assign v$SR_17424_out0 = v$SR_4532_out0;
assign v$SR_17425_out0 = v$SR_4533_out0;
assign v$SR_17426_out0 = v$SR_4534_out0;
assign v$SR_17427_out0 = v$SR_4535_out0;
assign v$SR_17428_out0 = v$SR_4536_out0;
assign v$SR_17429_out0 = v$SR_4537_out0;
assign v$SR_17430_out0 = v$SR_4538_out0;
assign v$SR_17431_out0 = v$SR_4539_out0;
assign v$EN_17562_out0 = v$EN_17005_out0;
assign v$EN_17563_out0 = v$EN_17006_out0;
assign v$EN_17564_out0 = v$EN_17007_out0;
assign v$EN_17566_out0 = v$EN_17009_out0;
assign v$EN_17567_out0 = v$EN_17010_out0;
assign v$EN_17568_out0 = v$EN_17011_out0;
assign v$G16_17575_out0 = v$EQ3_15864_out0 && v$G32_14802_out0;
assign v$G16_17576_out0 = v$EQ3_15865_out0 && v$G32_14803_out0;
assign v$INTERRUPT1_18306_out0 = v$EDGE1_18050_out0;
assign v$INTERRUPT1_18307_out0 = v$EDGE1_18051_out0;
assign v$G15_18435_out0 = v$G17_12250_out0 || v$G18_8726_out0;
assign v$G15_18436_out0 = v$G17_12251_out0 || v$G18_8727_out0;
assign v$IR1_18639_out0 = v$IR1_7941_out0;
assign v$IR1_18640_out0 = v$IR1_7942_out0;
assign v$IR1_706_out0 = v$IR1_18639_out0;
assign v$IR1_707_out0 = v$IR1_18640_out0;
assign v$R_1640_out0 = v$FINISHED_8327_out0;
assign v$R_1643_out0 = v$FINISHED_8328_out0;
assign v$G31_1983_out0 = v$G28_15272_out0 && v$IR1$IS$FPU$ARITHMETIC_1533_out0;
assign v$G31_1984_out0 = v$G28_15273_out0 && v$IR1$IS$FPU$ARITHMETIC_1534_out0;
assign v$SEL2_2628_out0 = v$IR1_18639_out0[15:12];
assign v$SEL2_2629_out0 = v$IR1_18640_out0[15:12];
assign v$EQ1_3042_out0 = v$SR_17425_out0 == 2'h1;
assign v$EQ1_3043_out0 = v$SR_17429_out0 == 2'h1;
assign v$EQ2_3431_out0 = v$SR_17427_out0 == 2'h2;
assign v$EQ2_3432_out0 = v$SR_17431_out0 == 2'h2;
assign v$G18_3607_out0 = v$INTERRUPT1_18306_out0 && v$G17_5717_out0;
assign v$G18_3608_out0 = v$INTERRUPT1_18307_out0 && v$G17_5718_out0;
assign v$TXINTERRUPT_3824_out0 = v$TXRST_8358_out0;
assign v$TXINTERRUPT_3825_out0 = v$TXRST_8359_out0;
assign v$IR1$FPU$OP_4019_out0 = v$SEL1_5457_out0;
assign v$IR1$FPU$OP_4020_out0 = v$SEL1_5458_out0;
assign v$IR1$D_4378_out0 = v$_16528_out0;
assign v$IR1$D_4379_out0 = v$_16529_out0;
assign v$G2_5263_out0 = v$Q3_18893_out0 && v$G3_4110_out0;
assign v$G2_5264_out0 = v$Q3_18894_out0 && v$G3_4111_out0;
assign v$EQ1_5291_out0 = v$SR_17426_out0 == 2'h1;
assign v$EQ1_5292_out0 = v$SR_17430_out0 == 2'h1;
assign v$EQ1_5299_out0 = v$SR_17424_out0 == 2'h3;
assign v$EQ1_5300_out0 = v$SR_17428_out0 == 2'h3;
assign v$G26_5343_out0 = v$G25_10727_out0 || v$FINISHED_8327_out0;
assign v$G26_5344_out0 = v$G25_10728_out0 || v$FINISHED_8328_out0;
assign v$G14_5626_out0 = v$G16_6650_out0 || v$G15_18435_out0;
assign v$G14_5627_out0 = v$G16_6651_out0 || v$G15_18436_out0;
assign v$EQ3_5676_out0 = v$SR_17426_out0 == 2'h3;
assign v$EQ3_5677_out0 = v$SR_17430_out0 == 2'h3;
assign v$IR1$OP_5761_out0 = v$_17304_out0;
assign v$IR1$OP_5762_out0 = v$_17305_out0;
assign v$IR1$15_6043_out0 = v$_13341_out0;
assign v$IR1$15_6044_out0 = v$_13342_out0;
assign v$MUX3_6396_out0 = v$G47_1685_out0 ? v$C3_19163_out0 : v$G29_3814_out0;
assign v$MUX3_6397_out0 = v$G47_1686_out0 ? v$C3_19164_out0 : v$G29_3815_out0;
assign v$G4_7870_out0 = v$G3_2634_out0 || v$G16_17575_out0;
assign v$G4_7871_out0 = v$G3_2635_out0 || v$G16_17576_out0;
assign v$IR1$S_8164_out0 = v$_14119_out0;
assign v$IR1$S_8165_out0 = v$_14120_out0;
assign v$IR1$32$BITS_8191_out0 = v$SEL13_13831_out0;
assign v$IR1$32$BITS_8192_out0 = v$SEL13_13832_out0;
assign v$EQ3_8225_out0 = v$SR_17424_out0 == 2'h1;
assign v$EQ3_8226_out0 = v$SR_17428_out0 == 2'h1;
assign v$EQ1_10860_out0 = v$SR_17427_out0 == 2'h3;
assign v$EQ1_10861_out0 = v$SR_17431_out0 == 2'h3;
assign v$OP_11500_out0 = v$OP_15388_out0;
assign v$OP_11501_out0 = v$OP_15389_out0;
assign v$_12326_out0 = { v$N_12539_out0,v$C1_5654_out0 };
assign v$_12327_out0 = { v$N_12540_out0,v$C1_5655_out0 };
assign v$G6_12509_out0 = v$IR2$VALID_13833_out0 && v$IR2$L_13058_out0;
assign v$G6_12510_out0 = v$IR2$VALID_13834_out0 && v$IR2$L_13059_out0;
assign v$EQ3_12702_out0 = v$SR_17427_out0 == 2'h1;
assign v$EQ3_12703_out0 = v$SR_17431_out0 == 2'h1;
assign v$IR1$M_13829_out0 = v$_6443_out0;
assign v$IR1$M_13830_out0 = v$_6444_out0;
assign v$G7_14136_out0 = v$G1_2078_out0 && v$G8_2607_out0;
assign v$G7_14137_out0 = v$G1_2079_out0 && v$G8_2608_out0;
assign v$EQ2_14201_out0 = v$SR_17425_out0 == 2'h2;
assign v$EQ2_14202_out0 = v$SR_17429_out0 == 2'h2;
assign v$EQ2_14904_out0 = v$SR_17424_out0 == 2'h2;
assign v$EQ2_14905_out0 = v$SR_17428_out0 == 2'h2;
assign v$FMUL$FINISHED_15076_out0 = v$FINISHED_8327_out0;
assign v$FMUL$FINISHED_15077_out0 = v$FINISHED_8328_out0;
assign v$G14_15285_out0 = ! v$INTERRUPT1_18306_out0;
assign v$G14_15286_out0 = ! v$INTERRUPT1_18307_out0;
assign v$EXEC2_16981_out0 = v$EXEC2_2109_out0;
assign v$EXEC2_16982_out0 = v$EXEC2_2110_out0;
assign v$EQ2_17012_out0 = v$SR_17426_out0 == 2'h2;
assign v$EQ2_17013_out0 = v$SR_17430_out0 == 2'h2;
assign v$G32_17032_out0 = v$INTERRUPT3_3708_out0 || v$COUNTERINTERRUPT_15460_out0;
assign v$G32_17033_out0 = v$INTERRUPT3_3709_out0 || v$COUNTERINTERRUPT_15461_out0;
assign v$EQ3_17164_out0 = v$SR_17425_out0 == 2'h3;
assign v$EQ3_17165_out0 = v$SR_17429_out0 == 2'h3;
assign v$EN_17561_out0 = v$EN_17004_out0;
assign v$EN_17565_out0 = v$EN_17008_out0;
assign v$TXReset_18441_out0 = v$TXRST_8358_out0;
assign v$TXReset_18442_out0 = v$TXRST_8359_out0;
assign v$G24_18545_out0 = v$IR2$VALID_13833_out0 && v$G23_14691_out0;
assign v$G24_18546_out0 = v$IR2$VALID_13834_out0 && v$G23_14692_out0;
assign v$N_18899_out0 = v$N_8578_out0;
assign v$N_18900_out0 = v$N_8579_out0;
assign v$G21_19292_out0 = v$IR2$VALID$AND$NOT$FLOAD_7603_out0 && v$EQ11_12455_out0;
assign v$G21_19293_out0 = v$IR2$VALID$AND$NOT$FLOAD_7604_out0 && v$EQ11_12456_out0;
assign v$R_1744_out0 = v$R_1640_out0;
assign v$R_1747_out0 = v$R_1643_out0;
assign v$N_1777_out0 = v$N_18899_out0;
assign v$N_1778_out0 = v$N_18900_out0;
assign v$G8_2050_out0 = v$EQ1_5299_out0 && v$EN_17561_out0;
assign v$G8_2051_out0 = v$EQ3_17164_out0 && v$EN_17562_out0;
assign v$G8_2052_out0 = v$EQ3_5676_out0 && v$EN_17563_out0;
assign v$G8_2053_out0 = v$EQ1_10860_out0 && v$EN_17564_out0;
assign v$G8_2054_out0 = v$EQ1_5300_out0 && v$EN_17565_out0;
assign v$G8_2055_out0 = v$EQ3_17165_out0 && v$EN_17566_out0;
assign v$G8_2056_out0 = v$EQ3_5677_out0 && v$EN_17567_out0;
assign v$G8_2057_out0 = v$EQ1_10861_out0 && v$EN_17568_out0;
assign v$NEXTENDED_2072_out0 = v$_12326_out0;
assign v$NEXTENDED_2073_out0 = v$_12327_out0;
assign v$G3_2800_out0 = v$EQ3_8225_out0 && v$EN_17561_out0;
assign v$G3_2801_out0 = v$EQ1_3042_out0 && v$EN_17562_out0;
assign v$G3_2802_out0 = v$EQ1_5291_out0 && v$EN_17563_out0;
assign v$G3_2803_out0 = v$EQ3_12702_out0 && v$EN_17564_out0;
assign v$G3_2804_out0 = v$EQ3_8226_out0 && v$EN_17565_out0;
assign v$G3_2805_out0 = v$EQ1_3043_out0 && v$EN_17566_out0;
assign v$G3_2806_out0 = v$EQ1_5292_out0 && v$EN_17567_out0;
assign v$G3_2807_out0 = v$EQ3_12703_out0 && v$EN_17568_out0;
assign v$MUX2_3090_out0 = v$IR2$VALID$AND$NOT$FLOAD_7603_out0 ? v$IR2$D_15090_out0 : v$IR1$M_13829_out0;
assign v$MUX2_3091_out0 = v$IR2$VALID$AND$NOT$FLOAD_7604_out0 ? v$IR2$D_15091_out0 : v$IR1$M_13830_out0;
assign v$OP_3869_out0 = v$OP_11500_out0;
assign v$OP_3870_out0 = v$OP_11501_out0;
assign v$EXEC2_4154_out0 = v$EXEC2_16981_out0;
assign v$EXEC2_4155_out0 = v$EXEC2_16982_out0;
assign v$G4_4186_out0 = v$EQ2_14904_out0 && v$EN_17561_out0;
assign v$G4_4187_out0 = v$EQ2_14201_out0 && v$EN_17562_out0;
assign v$G4_4188_out0 = v$EQ2_17012_out0 && v$EN_17563_out0;
assign v$G4_4189_out0 = v$EQ2_3431_out0 && v$EN_17564_out0;
assign v$G4_4190_out0 = v$EQ2_14905_out0 && v$EN_17565_out0;
assign v$G4_4191_out0 = v$EQ2_14202_out0 && v$EN_17566_out0;
assign v$G4_4192_out0 = v$EQ2_17013_out0 && v$EN_17567_out0;
assign v$G4_4193_out0 = v$EQ2_3432_out0 && v$EN_17568_out0;
assign v$EXEC2_4552_out0 = v$EXEC2_16981_out0;
assign v$EXEC2_4553_out0 = v$EXEC2_16982_out0;
assign v$G16_4639_out0 = v$FF2_17272_out0 && v$G14_15285_out0;
assign v$G16_4640_out0 = v$FF2_17273_out0 && v$G14_15286_out0;
assign v$TXINT_5126_out0 = v$TXINTERRUPT_3824_out0;
assign v$TXINT_5127_out0 = v$TXINTERRUPT_3825_out0;
assign v$Q2P_6320_out0 = v$MUX3_6396_out0;
assign v$Q2P_6321_out0 = v$MUX3_6397_out0;
assign v$G8_6340_out0 = v$G4_7870_out0 || v$G14_17632_out0;
assign v$G8_6341_out0 = v$G4_7871_out0 || v$G14_17633_out0;
assign v$EQ3_7548_out0 = v$IR1$FPU$OP_4019_out0 == 2'h2;
assign v$EQ3_7549_out0 = v$IR1$FPU$OP_4020_out0 == 2'h2;
assign v$EXEC2_8333_out0 = v$EXEC2_16981_out0;
assign v$EXEC2_8334_out0 = v$EXEC2_16982_out0;
assign v$G36_8364_out0 = v$G31_1983_out0 || v$G37_14699_out0;
assign v$G36_8365_out0 = v$G31_1984_out0 || v$G37_14700_out0;
assign v$EQ16_11237_out0 = v$IR1$FPU$OP_4019_out0 == 2'h3;
assign v$EQ16_11238_out0 = v$IR1$FPU$OP_4020_out0 == 2'h3;
assign v$RD_12364_out0 = v$IR1$D_4378_out0;
assign v$RD_12365_out0 = v$IR1$D_4379_out0;
assign v$S_13233_out0 = v$IR1$S_8164_out0;
assign v$S_13234_out0 = v$IR1$S_8165_out0;
assign v$G15_13976_out0 = v$G18_3607_out0 && v$R1_15628_out0;
assign v$G15_13977_out0 = v$G18_3608_out0 && v$R1_15629_out0;
assign v$FINISHED_14451_out0 = v$FMUL$FINISHED_15076_out0;
assign v$FINISHED_14452_out0 = v$FMUL$FINISHED_15077_out0;
assign v$INT3_14645_out0 = v$G32_17032_out0;
assign v$INT3_14646_out0 = v$G32_17033_out0;
assign v$G13_15713_out0 = v$NQ0_8120_out0 && v$G14_5626_out0;
assign v$G13_15714_out0 = v$NQ0_8121_out0 && v$G14_5627_out0;
assign v$G4_16428_out0 = ! v$IR1$15_6043_out0;
assign v$G4_16429_out0 = ! v$IR1$15_6044_out0;
assign v$IR1_16608_out0 = v$IR1_706_out0;
assign v$IR1_16609_out0 = v$IR1_707_out0;
assign v$EQ4_17130_out0 = v$IR1$FPU$OP_4019_out0 == 2'h2;
assign v$EQ4_17131_out0 = v$IR1$FPU$OP_4020_out0 == 2'h2;
assign v$IR1$FULL$OP$CODE_17650_out0 = v$SEL2_2628_out0;
assign v$IR1$FULL$OP$CODE_17651_out0 = v$SEL2_2629_out0;
assign v$EXEC2_18249_out0 = v$EXEC2_16981_out0;
assign v$EXEC2_18250_out0 = v$EXEC2_16982_out0;
assign v$N_18551_out0 = v$N_18899_out0;
assign v$N_18552_out0 = v$N_18900_out0;
assign v$R_18942_out0 = v$TXReset_18441_out0;
assign v$R_18953_out0 = v$TXReset_18442_out0;
assign v$WENALU_19270_out0 = v$G7_14136_out0;
assign v$WENALU_19271_out0 = v$G7_14137_out0;
assign v$_42_out0 = v$IR1_16608_out0[8:8];
assign v$_43_out0 = v$IR1_16609_out0[8:8];
assign v$FMUL$FINISHED_202_out0 = v$FINISHED_14451_out0;
assign v$FMUL$FINISHED_203_out0 = v$FINISHED_14452_out0;
assign v$EQ8_261_out0 = v$IR1$FULL$OP$CODE_17650_out0 == 4'h0;
assign v$EQ8_262_out0 = v$IR1$FULL$OP$CODE_17651_out0 == 4'h0;
assign v$_1012_out0 = v$IR1_16608_out0[11:10];
assign v$_1013_out0 = v$IR1_16609_out0[11:10];
assign v$EXEC2_1313_out0 = v$EXEC2_4552_out0;
assign v$EXEC2_1314_out0 = v$EXEC2_4553_out0;
assign v$EXEC2_1621_out0 = v$EXEC2_8333_out0;
assign v$EXEC2_1622_out0 = v$EXEC2_8334_out0;
assign v$EQ5_1657_out0 = v$IR1$FULL$OP$CODE_17650_out0 == 4'h1;
assign v$EQ5_1658_out0 = v$IR1$FULL$OP$CODE_17651_out0 == 4'h1;
assign v$INTERRUPT0_1967_out0 = v$TXINT_5126_out0;
assign v$INTERRUPT0_1968_out0 = v$TXINT_5127_out0;
assign v$_1999_out0 = v$IR1_16608_out0[5:2];
assign v$_2000_out0 = v$IR1_16609_out0[5:2];
assign v$EQ5_2074_out0 = v$OP_3869_out0 == 4'h6;
assign v$EQ5_2075_out0 = v$OP_3870_out0 == 4'h6;
assign v$_2130_out0 = v$IR1_16608_out0[6:6];
assign v$_2131_out0 = v$IR1_16609_out0[6:6];
assign v$EDGE3_2446_out0 = v$INT3_14645_out0;
assign v$EDGE3_2447_out0 = v$INT3_14646_out0;
assign v$_2640_out0 = v$IR1_16608_out0[9:9];
assign v$_2641_out0 = v$IR1_16609_out0[9:9];
assign v$_2866_out0 = { v$Q2P_6320_out0,v$Q3P_12238_out0 };
assign v$_2867_out0 = { v$Q2P_6321_out0,v$Q3P_12239_out0 };
assign v$WENALU_4228_out0 = v$WENALU_19270_out0;
assign v$WENALU_4229_out0 = v$WENALU_19271_out0;
assign v$EQ1_4267_out0 = v$OP_3869_out0 == 4'h2;
assign v$EQ1_4268_out0 = v$OP_3870_out0 == 4'h2;
assign v$EQ3_6015_out0 = v$OP_3869_out0 == 4'h4;
assign v$EQ3_6016_out0 = v$OP_3870_out0 == 4'h4;
assign v$_7607_out0 = v$IR1_16608_out0[7:7];
assign v$_7608_out0 = v$IR1_16609_out0[7:7];
assign v$EXEC2_8362_out0 = v$EXEC2_18249_out0;
assign v$EXEC2_8363_out0 = v$EXEC2_18250_out0;
assign v$MUX16_9038_out0 = v$FINISHED_14451_out0 ? v$RD$FPU_13518_out0 : v$MUX2_3090_out0;
assign v$MUX16_9039_out0 = v$FINISHED_14452_out0 ? v$RD$FPU_13519_out0 : v$MUX2_3091_out0;
assign v$EQ13_9710_out0 = v$IR1$FULL$OP$CODE_17650_out0 == 4'h1;
assign v$EQ13_9711_out0 = v$IR1$FULL$OP$CODE_17651_out0 == 4'h1;
assign v$EQ4_9727_out0 = v$OP_3869_out0 == 4'h5;
assign v$EQ4_9728_out0 = v$OP_3870_out0 == 4'h5;
assign v$EXEC2_9813_out0 = v$EXEC2_4154_out0;
assign v$EXEC2_9814_out0 = v$EXEC2_4155_out0;
assign v$_11286_out0 = v$IR1_16608_out0[1:0];
assign v$_11287_out0 = v$IR1_16609_out0[1:0];
assign v$EQ2_11292_out0 = v$OP_3869_out0 == 4'h3;
assign v$EQ2_11293_out0 = v$OP_3870_out0 == 4'h3;
assign v$N_12322_out0 = v$N_18551_out0;
assign v$N_12323_out0 = v$N_18552_out0;
assign v$EQ14_12688_out0 = v$IR1$FULL$OP$CODE_17650_out0 == 4'h1;
assign v$EQ14_12689_out0 = v$IR1$FULL$OP$CODE_17651_out0 == 4'h1;
assign v$_13333_out0 = v$IR1_16608_out0[15:15];
assign v$_13334_out0 = v$IR1_16609_out0[15:15];
assign v$NEXTENDED_14977_out0 = v$NEXTENDED_2072_out0;
assign v$NEXTENDED_14978_out0 = v$NEXTENDED_2073_out0;
assign v$G13_15463_out0 = v$G8_6340_out0 || v$G12_6432_out0;
assign v$G13_15464_out0 = v$G8_6341_out0 || v$G12_6433_out0;
assign v$G1_15877_out0 = v$G2_5263_out0 || v$G13_15713_out0;
assign v$G1_15878_out0 = v$G2_5264_out0 || v$G13_15714_out0;
assign v$G6_16157_out0 = ! v$R_18942_out0;
assign v$G6_16168_out0 = ! v$R_18953_out0;
assign v$EQ15_16391_out0 = v$IR1$FULL$OP$CODE_17650_out0 == 4'h1;
assign v$EQ15_16392_out0 = v$IR1$FULL$OP$CODE_17651_out0 == 4'h1;
assign v$EQ2_16405_out0 = v$IR1_16608_out0 == 16'h7000;
assign v$EQ2_16406_out0 = v$IR1_16609_out0 == 16'h7000;
assign v$_16655_out0 = v$IR1_16608_out0[15:12];
assign v$_16656_out0 = v$IR1_16609_out0[15:12];
assign v$EQ6_16860_out0 = v$OP_3869_out0 == 4'h7;
assign v$EQ6_16861_out0 = v$OP_3870_out0 == 4'h7;
assign v$S_17002_out0 = v$S_13233_out0;
assign v$S_17003_out0 = v$S_13234_out0;
assign v$G13_17152_out0 = v$G16_4639_out0 && v$F1_3687_out0;
assign v$G13_17153_out0 = v$G16_4640_out0 && v$F1_3688_out0;
assign v$END_17218_out0 = v$N_1777_out0;
assign v$END_17219_out0 = v$N_1778_out0;
assign v$G3_18294_out0 = ! v$R_1744_out0;
assign v$G3_18297_out0 = ! v$R_1747_out0;
assign v$JMI_72_out0 = v$EQ4_9727_out0;
assign v$JMI_73_out0 = v$EQ4_9728_out0;
assign v$G5_1267_out0 = v$FF2_13621_out0 && v$G6_16157_out0;
assign v$G5_1272_out0 = v$FF2_13632_out0 && v$G6_16168_out0;
assign v$JMP_1825_out0 = v$EQ3_6015_out0;
assign v$JMP_1826_out0 = v$EQ3_6016_out0;
assign v$JLS_2120_out0 = v$EQ2_11292_out0;
assign v$JLS_2121_out0 = v$EQ2_11293_out0;
assign v$INTERRUPT3_3040_out0 = v$EDGE3_2446_out0;
assign v$INTERRUPT3_3041_out0 = v$EDGE3_2447_out0;
assign v$IR1$OPCODE_3102_out0 = v$_16655_out0;
assign v$IR1$OPCODE_3103_out0 = v$_16656_out0;
assign v$INT2_3379_out0 = v$FMUL$FINISHED_202_out0;
assign v$INT2_3380_out0 = v$FMUL$FINISHED_203_out0;
assign v$G25_3750_out0 = ! v$EQ14_12688_out0;
assign v$G25_3751_out0 = ! v$EQ14_12689_out0;
assign v$IR1$P_3871_out0 = v$_7607_out0;
assign v$IR1$P_3872_out0 = v$_7608_out0;
assign v$IR1$L_5356_out0 = v$_2640_out0;
assign v$IR1$L_5357_out0 = v$_2641_out0;
assign v$EDGE0_6025_out0 = v$INTERRUPT0_1967_out0;
assign v$EDGE0_6026_out0 = v$INTERRUPT0_1968_out0;
assign v$STP_6467_out0 = v$EQ6_16860_out0;
assign v$STP_6468_out0 = v$EQ6_16861_out0;
assign v$STOP$1_8134_out0 = v$EQ2_16405_out0;
assign v$STOP$1_8135_out0 = v$EQ2_16406_out0;
assign v$Q0P_12736_out0 = v$G1_15877_out0;
assign v$Q0P_12737_out0 = v$G1_15878_out0;
assign v$IR1$M_13215_out0 = v$_11286_out0;
assign v$IR1$M_13216_out0 = v$_11287_out0;
assign v$G1_13555_out0 = v$STATE_16625_out0 && v$G3_18294_out0;
assign v$G1_13558_out0 = v$STATE_16628_out0 && v$G3_18297_out0;
assign v$EQ10_13993_out0 = v$N_12322_out0 == 12'h2;
assign v$EQ10_13994_out0 = v$N_12323_out0 == 12'h2;
assign v$EQ11_14182_out0 = v$N_12322_out0 == 12'h4;
assign v$EQ11_14183_out0 = v$N_12323_out0 == 12'h4;
assign v$G28_14373_out0 = v$EQ16_11237_out0 && v$EQ15_16391_out0;
assign v$G28_14374_out0 = v$EQ16_11238_out0 && v$EQ15_16392_out0;
assign v$EQ8_14932_out0 = v$N_12322_out0 == 12'h0;
assign v$EQ8_14933_out0 = v$N_12323_out0 == 12'h0;
assign v$IR1$U_15384_out0 = v$_2130_out0;
assign v$IR1$U_15385_out0 = v$_2131_out0;
assign v$IR1$D_15458_out0 = v$_1012_out0;
assign v$IR1$D_15459_out0 = v$_1013_out0;
assign v$JLO_15598_out0 = v$EQ1_4267_out0;
assign v$JLO_15599_out0 = v$EQ1_4268_out0;
assign v$AD3_15754_out0 = v$MUX16_9038_out0;
assign v$AD3_15755_out0 = v$MUX16_9039_out0;
assign v$G22_16224_out0 = v$EQ4_17130_out0 && v$EQ13_9710_out0;
assign v$G22_16225_out0 = v$EQ4_17131_out0 && v$EQ13_9711_out0;
assign v$IR1$N_16365_out0 = v$_1999_out0;
assign v$IR1$N_16366_out0 = v$_2000_out0;
assign v$IR1$LS_17045_out0 = v$_13333_out0;
assign v$IR1$LS_17046_out0 = v$_13334_out0;
assign v$IR1$W_17168_out0 = v$_42_out0;
assign v$IR1$W_17169_out0 = v$_43_out0;
assign v$G5_17176_out0 = v$EQ3_7548_out0 && v$EQ5_1657_out0;
assign v$G5_17177_out0 = v$EQ3_7549_out0 && v$EQ5_1658_out0;
assign v$G19_17314_out0 = v$G15_13976_out0 || v$G13_17152_out0;
assign v$G19_17315_out0 = v$G15_13977_out0 || v$G13_17153_out0;
assign v$G23_17391_out0 = v$G13_15463_out0 || v$G26_13755_out0;
assign v$G23_17392_out0 = v$G13_15464_out0 || v$G26_13756_out0;
assign v$EQ7_17509_out0 = v$N_12322_out0 == 12'h1;
assign v$EQ7_17510_out0 = v$N_12323_out0 == 12'h1;
assign v$G2_17660_out0 = v$S_17002_out0 && v$EXEC2_448_out0;
assign v$G2_17661_out0 = v$S_17003_out0 && v$EXEC2_449_out0;
assign v$EQ9_18380_out0 = v$N_12322_out0 == 12'h3;
assign v$EQ9_18381_out0 = v$N_12323_out0 == 12'h3;
assign v$JEQ_18641_out0 = v$EQ5_2074_out0;
assign v$JEQ_18642_out0 = v$EQ5_2075_out0;
assign v$EQ13_19159_out0 = v$N_12322_out0 == 12'h5;
assign v$EQ13_19160_out0 = v$N_12323_out0 == 12'h5;
assign v$JEQ_1833_out0 = v$JEQ_18641_out0;
assign v$JEQ_1834_out0 = v$JEQ_18642_out0;
assign v$G32_1987_out0 = v$INTERRUPT3_3040_out0 && v$G31_10014_out0;
assign v$G32_1988_out0 = v$INTERRUPT3_3041_out0 && v$G31_10015_out0;
assign v$G3_2868_out0 = v$G2_17660_out0 && v$G4_12565_out0;
assign v$G3_2869_out0 = v$G2_17661_out0 && v$G4_12566_out0;
assign v$G28_3387_out0 = ! v$INTERRUPT3_3040_out0;
assign v$G28_3388_out0 = ! v$INTERRUPT3_3041_out0;
assign v$INTERRUPT2_4034_out0 = v$INT2_3379_out0;
assign v$INTERRUPT2_4035_out0 = v$INT2_3380_out0;
assign v$JMP_4500_out0 = v$JMP_1825_out0;
assign v$JMP_4501_out0 = v$JMP_1826_out0;
assign v$_5301_out0 = { v$Q0P_12736_out0,v$Q1P_11515_out0 };
assign v$_5302_out0 = { v$Q0P_12737_out0,v$Q1P_11516_out0 };
assign v$JLO_8424_out0 = v$JLO_15598_out0;
assign v$JLO_8425_out0 = v$JLO_15599_out0;
assign v$IR1$IS$FPU$LOAD$STORE_9261_out0 = v$G28_14373_out0;
assign v$IR1$IS$FPU$LOAD$STORE_9262_out0 = v$G28_14374_out0;
assign v$_12208_out0 = { v$IR1$N_16365_out0,v$C4_16509_out0 };
assign v$_12209_out0 = { v$IR1$N_16366_out0,v$C4_16510_out0 };
assign v$INTERRUPT0_12268_out0 = v$EDGE0_6025_out0;
assign v$INTERRUPT0_12269_out0 = v$EDGE0_6026_out0;
assign v$STP_12282_out0 = v$STP_6467_out0;
assign v$STP_12283_out0 = v$STP_6468_out0;
assign v$G16_12541_out0 = ! v$IR1$W_17168_out0;
assign v$G16_12542_out0 = ! v$IR1$W_17169_out0;
assign v$AD3_13721_out0 = v$AD3_15754_out0;
assign v$AD3_13722_out0 = v$AD3_15755_out0;
assign v$JMI_13727_out0 = v$JMI_72_out0;
assign v$JMI_13728_out0 = v$JMI_73_out0;
assign v$G24_14443_out0 = v$G25_3750_out0 && v$G4_16428_out0;
assign v$G24_14444_out0 = v$G25_3751_out0 && v$G4_16429_out0;
assign v$EQ5_14979_out0 = v$IR1$OPCODE_3102_out0 == 4'h0;
assign v$EQ5_14980_out0 = v$IR1$OPCODE_3103_out0 == 4'h0;
assign v$G10_15507_out0 = ! v$STOP$1_8134_out0;
assign v$G10_15508_out0 = ! v$STOP$1_8135_out0;
assign v$EDGE1_15855_out0 = v$G19_17314_out0;
assign v$EDGE1_15856_out0 = v$G19_17315_out0;
assign v$IS$IR1$FMUL_15879_out0 = v$G22_16224_out0;
assign v$IS$IR1$FMUL_15880_out0 = v$G22_16225_out0;
assign v$JLS_17065_out0 = v$JLS_2120_out0;
assign v$JLS_17066_out0 = v$JLS_2121_out0;
assign v$G27_17148_out0 = v$G23_17391_out0 || v$G36_8364_out0;
assign v$G27_17149_out0 = v$G23_17392_out0 || v$G36_8365_out0;
assign v$EQ3_18535_out0 = v$IR1$OPCODE_3102_out0 == 4'h0;
assign v$EQ3_18536_out0 = v$IR1$OPCODE_3103_out0 == 4'h0;
assign v$G2_19037_out0 = ! v$IR1$L_5356_out0;
assign v$G2_19038_out0 = ! v$IR1$L_5357_out0;
assign v$G8_19390_out0 = ! v$IR1$U_15384_out0;
assign v$G8_19391_out0 = ! v$IR1$U_15385_out0;
assign v$_1382_out0 = { v$_5301_out0,v$_13641_out0 };
assign v$_1383_out0 = { v$_5302_out0,v$_13642_out0 };
assign v$DIN_1883_out0 = v$_12208_out0;
assign v$DIN_1884_out0 = v$_12209_out0;
assign v$G27_4064_out0 = ! v$IR1$IS$FPU$LOAD$STORE_9261_out0;
assign v$G27_4065_out0 = ! v$IR1$IS$FPU$LOAD$STORE_9262_out0;
assign v$G17_5699_out0 = v$JLO_8424_out0 && v$G18_14086_out0;
assign v$G17_5700_out0 = v$JLO_8425_out0 && v$G18_14087_out0;
assign v$G29_5727_out0 = v$G32_1987_out0 && v$R3_15899_out0;
assign v$G29_5728_out0 = v$G32_1988_out0 && v$R3_15900_out0;
assign v$G9_6085_out0 = ! v$INTERRUPT0_12268_out0;
assign v$G9_6086_out0 = ! v$INTERRUPT0_12269_out0;
assign v$MUX17_6767_out0 = v$IS$IR1$FMUL_15879_out0 ? v$IR1$32$BITS_8191_out0 : v$IR2$FPU$32BIT_12372_out0;
assign v$MUX17_6768_out0 = v$IS$IR1$FMUL_15880_out0 ? v$IR1$32$BITS_8192_out0 : v$IR2$FPU$32BIT_12373_out0;
assign v$EDGE2_7280_out0 = v$INTERRUPT2_4034_out0;
assign v$EDGE2_7281_out0 = v$INTERRUPT2_4035_out0;
assign v$G5_7910_out0 = v$G3_2868_out0 && v$IR15_11494_out0;
assign v$G5_7911_out0 = v$G3_2869_out0 && v$IR15_11495_out0;
assign v$G20_12774_out0 = v$EQ5_14979_out0 && v$IR1$L_5356_out0;
assign v$G20_12775_out0 = v$EQ5_14980_out0 && v$IR1$L_5357_out0;
assign v$SUBEN_13429_out0 = v$G8_19390_out0;
assign v$SUBEN_13430_out0 = v$G8_19391_out0;
assign v$STALL_13723_out0 = v$G27_17148_out0;
assign v$STALL_13724_out0 = v$G27_17149_out0;
assign v$G3_14794_out0 = v$EQ3_18535_out0 && v$G2_19037_out0;
assign v$G3_14795_out0 = v$EQ3_18536_out0 && v$G2_19038_out0;
assign v$G7_15277_out0 = v$INTERRUPT0_12268_out0 && v$G1_15078_out0;
assign v$G7_15278_out0 = v$INTERRUPT0_12269_out0 && v$G1_15079_out0;
assign v$G30_16506_out0 = v$FF4_19047_out0 && v$G28_3387_out0;
assign v$G30_16507_out0 = v$FF4_19048_out0 && v$G28_3388_out0;
assign v$STP_18374_out0 = v$STP_12282_out0;
assign v$STP_18375_out0 = v$STP_12283_out0;
assign v$G15_19147_out0 = v$IR1$P_3871_out0 || v$G16_12541_out0;
assign v$G15_19148_out0 = v$IR1$P_3872_out0 || v$G16_12542_out0;
assign v$INTERRUPT2_1821_out0 = v$EDGE2_7280_out0;
assign v$INTERRUPT2_1822_out0 = v$EDGE2_7281_out0;
assign v$G27_2708_out0 = v$G30_16506_out0 && v$F3_8557_out0;
assign v$G27_2709_out0 = v$G30_16507_out0 && v$F3_8558_out0;
assign v$G8_6328_out0 = v$G7_15277_out0 && v$R0_15792_out0;
assign v$G8_6329_out0 = v$G7_15278_out0 && v$R0_15793_out0;
assign v$G43_7337_out0 = v$STALL_13723_out0 && v$IR2$VALID_4376_out0;
assign v$G43_7338_out0 = v$STALL_13724_out0 && v$IR2$VALID_4377_out0;
assign v$STP_11314_out0 = v$STP_18374_out0;
assign v$STP_11315_out0 = v$STP_18375_out0;
assign v$32BIT_11437_out0 = v$MUX17_6767_out0;
assign v$32BIT_11438_out0 = v$MUX17_6768_out0;
assign v$MUX1_12320_out0 = v$SUBEN_13429_out0 ? v$C2_12772_out0 : v$C1_18809_out0;
assign v$MUX1_12321_out0 = v$SUBEN_13430_out0 ? v$C2_12773_out0 : v$C1_18810_out0;
assign v$G10_13900_out0 = v$FF1_6306_out0 && v$G9_6085_out0;
assign v$G10_13901_out0 = v$FF1_6307_out0 && v$G9_6086_out0;
assign v$G26_18725_out0 = v$IS$IR1$FMUL_15879_out0 && v$G27_4064_out0;
assign v$G26_18726_out0 = v$IS$IR1$FMUL_15880_out0 && v$G27_4065_out0;
assign v$QP_19149_out0 = v$_1382_out0;
assign v$QP_19150_out0 = v$_1383_out0;
assign v$G10_1329_out0 = v$EQ11_14182_out0 && v$STP_11314_out0;
assign v$G10_1330_out0 = v$EQ11_14183_out0 && v$STP_11315_out0;
assign v$G33_1384_out0 = v$G29_5727_out0 || v$G27_2708_out0;
assign v$G33_1385_out0 = v$G29_5728_out0 || v$G27_2709_out0;
assign v$G11_1775_out0 = v$G10_13900_out0 && v$F0_16438_out0;
assign v$G11_1776_out0 = v$G10_13901_out0 && v$F0_16439_out0;
assign v$G8_2448_out0 = v$EQ9_18380_out0 && v$STP_11314_out0;
assign v$G8_2449_out0 = v$EQ9_18381_out0 && v$STP_11315_out0;
assign v$G7_3377_out0 = v$EQ10_13993_out0 && v$STP_11314_out0;
assign v$G7_3378_out0 = v$EQ10_13994_out0 && v$STP_11315_out0;
assign v$MUX11_4657_out0 = v$G26_18725_out0 ? v$IR1$FPU$OP_4019_out0 : v$IR2$FPU$OP_1845_out0;
assign v$MUX11_4658_out0 = v$G26_18726_out0 ? v$IR1$FPU$OP_4020_out0 : v$IR2$FPU$OP_1846_out0;
assign v$G12_5046_out0 = v$G43_7337_out0 && v$INITIAL$FETCH$OCCURRED_1691_out0;
assign v$G12_5047_out0 = v$G43_7338_out0 && v$INITIAL$FETCH$OCCURRED_1692_out0;
assign v$XOR1_5297_out0 = v$MUX1_12320_out0 ^ v$DIN_1883_out0;
assign v$XOR1_5298_out0 = v$MUX1_12321_out0 ^ v$DIN_1884_out0;
assign v$G6_5703_out0 = v$EQ7_17509_out0 && v$STP_11314_out0;
assign v$G6_5704_out0 = v$EQ7_17510_out0 && v$STP_11315_out0;
assign v$G14_6671_out0 = v$EQ13_19159_out0 && v$STP_11314_out0;
assign v$G14_6672_out0 = v$EQ13_19160_out0 && v$STP_11315_out0;
assign v$G21_7321_out0 = ! v$INTERRUPT2_1821_out0;
assign v$G21_7322_out0 = ! v$INTERRUPT2_1822_out0;
assign v$EQ5_10454_out0 = v$QP_19149_out0 == 4'hb;
assign v$EQ5_10455_out0 = v$QP_19150_out0 == 4'hb;
assign v$G25_15179_out0 = v$INTERRUPT2_1821_out0 && v$G24_12651_out0;
assign v$G25_15180_out0 = v$INTERRUPT2_1822_out0 && v$G24_12652_out0;
assign v$G9_15733_out0 = v$EQ8_14932_out0 && v$STP_11314_out0;
assign v$G9_15734_out0 = v$EQ8_14933_out0 && v$STP_11315_out0;
assign v$32BIT_16476_out0 = v$32BIT_11437_out0;
assign v$32BIT_16477_out0 = v$32BIT_11438_out0;
assign v$OP_1485_out0 = v$MUX11_4657_out0;
assign v$OP_1486_out0 = v$MUX11_4658_out0;
assign v$G37_1523_out0 = v$G12_5046_out0 && v$G48_5092_out0;
assign v$G37_1524_out0 = v$G12_5047_out0 && v$G48_5093_out0;
assign v$INTDISABLE_5214_out0 = v$G7_3377_out0;
assign v$INTDISABLE_5215_out0 = v$G7_3378_out0;
assign v$G22_5701_out0 = v$G25_15179_out0 && v$R2_4026_out0;
assign v$G22_5702_out0 = v$G25_15180_out0 && v$R2_4027_out0;
assign v$NEXTINT_7282_out0 = v$G10_1329_out0;
assign v$NEXTINT_7283_out0 = v$G10_1330_out0;
assign v$INTCLEAR_8096_out0 = v$G8_2448_out0;
assign v$INTCLEAR_8097_out0 = v$G8_2449_out0;
assign v$G23_9982_out0 = v$FF3_15648_out0 && v$G21_7321_out0;
assign v$G23_9983_out0 = v$FF3_15649_out0 && v$G21_7322_out0;
assign v$G29_11326_out0 = v$32BIT_16476_out0 && v$IR2$IS$FPU_12415_out0;
assign v$G29_11327_out0 = v$32BIT_16477_out0 && v$IR2$IS$FPU_12416_out0;
assign v$IS$32$BIT_11513_out0 = v$32BIT_16476_out0;
assign v$IS$32$BIT_11514_out0 = v$32BIT_16477_out0;
assign v$EDGE3_11552_out0 = v$G33_1384_out0;
assign v$EDGE3_11553_out0 = v$G33_1385_out0;
assign v$LDMAINPC_14212_out0 = v$G14_6671_out0;
assign v$LDMAINPC_14213_out0 = v$G14_6672_out0;
assign v$IS$32$BITS_14649_out0 = v$32BIT_16476_out0;
assign v$IS$32$BITS_14650_out0 = v$32BIT_16477_out0;
assign v$G12_15311_out0 = v$G8_6328_out0 || v$G11_1775_out0;
assign v$G12_15312_out0 = v$G8_6329_out0 || v$G11_1776_out0;
assign v$G66_17456_out0 = !(v$G69_1355_out0 && v$EQ5_10454_out0);
assign v$G66_17457_out0 = !(v$G69_1356_out0 && v$EQ5_10455_out0);
assign v$NEXTINTERRUPT_19157_out0 = v$G10_1329_out0;
assign v$NEXTINTERRUPT_19158_out0 = v$G10_1330_out0;
assign v$INTCLR_220_out0 = v$INTCLEAR_8096_out0;
assign v$INTCLR_221_out0 = v$INTCLEAR_8097_out0;
assign v$G35_1289_out0 = v$G37_1523_out0 && v$G36_17991_out0;
assign v$G35_1290_out0 = v$G37_1524_out0 && v$G36_17992_out0;
assign v$INTDISABLE_2882_out0 = v$INTDISABLE_5214_out0;
assign v$INTDISABLE_2883_out0 = v$INTDISABLE_5215_out0;
assign v$EDGE0_4146_out0 = v$G12_15311_out0;
assign v$EDGE0_4147_out0 = v$G12_15312_out0;
assign v$G34_5132_out0 = v$NEXTINTERRUPT_19157_out0 || v$FF2_1327_out0;
assign v$G34_5133_out0 = v$NEXTINTERRUPT_19158_out0 || v$FF2_1328_out0;
assign v$IS$32$BIT_11362_out0 = v$IS$32$BIT_11513_out0;
assign v$IS$32$BIT_11363_out0 = v$IS$32$BIT_11514_out0;
assign v$G20_12278_out0 = v$G23_9982_out0 && v$F2_12662_out0;
assign v$G20_12279_out0 = v$G23_9983_out0 && v$F2_12663_out0;
assign v$G15_14005_out0 = v$G6_5703_out0 || v$NEXTINT_7282_out0;
assign v$G15_14006_out0 = v$G6_5704_out0 || v$NEXTINT_7283_out0;
assign v$LDMAIN_14395_out0 = v$LDMAINPC_14212_out0;
assign v$LDMAIN_14396_out0 = v$LDMAINPC_14213_out0;
assign v$FPU$OP_14679_out0 = v$OP_1485_out0;
assign v$FPU$OP_14680_out0 = v$OP_1486_out0;
assign v$G65_14732_out0 = v$G66_17456_out0 && v$CLK4_2728_out0;
assign v$G65_14733_out0 = v$G66_17457_out0 && v$CLK4_2729_out0;
assign v$CLRINTERRUPTS_356_out0 = v$INTCLR_220_out0;
assign v$CLRINTERRUPTS_357_out0 = v$INTCLR_221_out0;
assign v$INTENABLE_3148_out0 = v$G15_14005_out0;
assign v$INTENABLE_3149_out0 = v$G15_14006_out0;
assign v$EQ5_3178_out0 = v$FPU$OP_14679_out0 == 2'h3;
assign v$EQ5_3179_out0 = v$FPU$OP_14680_out0 == 2'h3;
assign v$EQ2_4388_out0 = v$FPU$OP_14679_out0 == 2'h0;
assign v$EQ2_4389_out0 = v$FPU$OP_14680_out0 == 2'h0;
assign v$G26_10775_out0 = v$G22_5701_out0 || v$G20_12278_out0;
assign v$G26_10776_out0 = v$G22_5702_out0 || v$G20_12279_out0;
assign v$G35_10777_out0 = v$INTDISABLE_2882_out0 || v$AUTODISABLE_18814_out0;
assign v$G35_10778_out0 = v$INTDISABLE_2883_out0 || v$AUTODISABLE_18815_out0;
assign v$STOPBITERROR_12296_out0 = v$G65_14732_out0;
assign v$STOPBITERROR_12297_out0 = v$G65_14733_out0;
assign v$FPU$OP_13331_out0 = v$FPU$OP_14679_out0;
assign v$FPU$OP_13332_out0 = v$FPU$OP_14680_out0;
assign v$EQ7_14178_out0 = v$FPU$OP_14679_out0 == 2'h2;
assign v$EQ7_14179_out0 = v$FPU$OP_14680_out0 == 2'h2;
assign v$EQ3_14381_out0 = v$FPU$OP_14679_out0 == 2'h2;
assign v$EQ3_14382_out0 = v$FPU$OP_14680_out0 == 2'h2;
assign v$EQ1_15873_out0 = v$FPU$OP_14679_out0 == 2'h1;
assign v$EQ1_15874_out0 = v$FPU$OP_14680_out0 == 2'h1;
assign v$G5_16393_out0 = ! v$IS$32$BIT_11362_out0;
assign v$G5_16394_out0 = ! v$IS$32$BIT_11363_out0;
assign v$EQ8_16631_out0 = v$FPU$OP_14679_out0 == 2'h3;
assign v$EQ8_16632_out0 = v$FPU$OP_14680_out0 == 2'h3;
assign v$EQ4_17319_out0 = v$FPU$OP_14679_out0 == 2'h3;
assign v$EQ4_17320_out0 = v$FPU$OP_14680_out0 == 2'h3;
assign v$STALL_18502_out0 = v$G35_1289_out0;
assign v$STALL_18503_out0 = v$G35_1290_out0;
assign v$NEXTINTERRUPT_19041_out0 = v$G34_5132_out0;
assign v$NEXTINTERRUPT_19042_out0 = v$G34_5133_out0;
assign v$STOPERROR_306_out0 = v$STOPBITERROR_12296_out0;
assign v$STOPERROR_307_out0 = v$STOPBITERROR_12297_out0;
assign v$G30_3945_out0 = ! v$EQ8_16631_out0;
assign v$G30_3946_out0 = ! v$EQ8_16632_out0;
assign v$CLR_4601_out0 = v$CLRINTERRUPTS_356_out0;
assign v$CLR_4602_out0 = v$CLRINTERRUPTS_357_out0;
assign v$G49_5461_out0 = ! v$STALL_18502_out0;
assign v$G49_5462_out0 = ! v$STALL_18503_out0;
assign v$ADD_8527_out0 = v$EQ2_4388_out0;
assign v$ADD_8528_out0 = v$EQ2_4389_out0;
assign v$FPU$LOAD$STORE_11486_out0 = v$EQ4_17319_out0;
assign v$FPU$LOAD$STORE_11487_out0 = v$EQ4_17320_out0;
assign v$G12_12555_out0 = v$G11_13991_out0 && v$EQ5_3178_out0;
assign v$G12_12556_out0 = v$G11_13992_out0 && v$EQ5_3179_out0;
assign v$NEXTINTERRUPT_13321_out0 = v$NEXTINTERRUPT_19041_out0;
assign v$NEXTINTERRUPT_13322_out0 = v$NEXTINTERRUPT_19042_out0;
assign v$SUB_14377_out0 = v$EQ1_15873_out0;
assign v$SUB_14378_out0 = v$EQ1_15874_out0;
assign v$DISABLEINTERRUPTS_15588_out0 = v$G35_10777_out0;
assign v$DISABLEINTERRUPTS_15589_out0 = v$G35_10778_out0;
assign v$STALL_16085_out0 = v$STALL_18502_out0;
assign v$STALL_16086_out0 = v$STALL_18503_out0;
assign v$EQ1_16829_out0 = v$FPU$OP_13331_out0 == 2'h1;
assign v$EQ1_16830_out0 = v$FPU$OP_13332_out0 == 2'h1;
assign v$MUL_17628_out0 = v$EQ3_14381_out0;
assign v$MUL_17629_out0 = v$EQ3_14382_out0;
assign v$INTENABLE_18046_out0 = v$INTENABLE_3148_out0;
assign v$INTENABLE_18047_out0 = v$INTENABLE_3149_out0;
assign v$EDGE2_18729_out0 = v$G26_10775_out0;
assign v$EDGE2_18730_out0 = v$G26_10776_out0;
assign v$G31_2537_out0 = v$G29_11326_out0 && v$G30_3945_out0;
assign v$G31_2538_out0 = v$G29_11327_out0 && v$G30_3946_out0;
assign v$G2_3905_out0 = v$ADD_8527_out0 || v$SUB_14377_out0;
assign v$G2_3906_out0 = v$ADD_8528_out0 || v$SUB_14378_out0;
assign v$G4_5116_out0 = v$ERR_13343_out0 || v$STOPERROR_306_out0;
assign v$G4_5117_out0 = v$ERR_13344_out0 || v$STOPERROR_307_out0;
assign v$G6_8265_out0 = v$ADD_8527_out0 || v$SUB_14377_out0;
assign v$G6_8266_out0 = v$ADD_8528_out0 || v$SUB_14378_out0;
assign v$G28_9040_out0 = v$FPU$LOAD$STORE_11486_out0 && v$LOAD_6451_out0;
assign v$G28_9041_out0 = v$FPU$LOAD$STORE_11487_out0 && v$LOAD_6452_out0;
assign v$G27_11224_out0 = v$FPU$LOAD$STORE_11486_out0 && v$LOAD_6451_out0;
assign v$G27_11225_out0 = v$FPU$LOAD$STORE_11487_out0 && v$LOAD_6452_out0;
assign v$G27_12276_out0 = v$STP$DECODED_17154_out0 || v$G49_5461_out0;
assign v$G27_12277_out0 = v$STP$DECODED_17155_out0 || v$G49_5462_out0;
assign v$STALL_12797_out0 = v$STALL_16085_out0;
assign v$STALL_12798_out0 = v$STALL_16086_out0;
assign v$ENABLEINTERRUPTS_13141_out0 = v$INTENABLE_18046_out0;
assign v$ENABLEINTERRUPTS_13142_out0 = v$INTENABLE_18047_out0;
assign v$G21_15317_out0 = v$G20_12859_out0 && v$FPU$LOAD$STORE_11486_out0;
assign v$G21_15318_out0 = v$G20_12860_out0 && v$FPU$LOAD$STORE_11487_out0;
assign v$NEXTINTERRUPT_17397_out0 = v$NEXTINTERRUPT_13321_out0;
assign v$NEXTINTERRUPT_17398_out0 = v$NEXTINTERRUPT_13322_out0;
assign v$R_18937_out0 = v$DISABLEINTERRUPTS_15588_out0;
assign v$R_18940_out0 = v$CLR_4601_out0;
assign v$R_18948_out0 = v$DISABLEINTERRUPTS_15589_out0;
assign v$R_18951_out0 = v$CLR_4602_out0;
assign v$G8_1401_out0 = v$G27_11224_out0 && v$LOADA_5295_out0;
assign v$G8_1402_out0 = v$G27_11225_out0 && v$LOADA_5296_out0;
assign v$G3_4262_out0 = v$I0P_4512_out0 && v$NEXTINTERRUPT_17397_out0;
assign v$G3_4263_out0 = v$I0P_4513_out0 && v$NEXTINTERRUPT_17398_out0;
assign v$G1_7537_out0 = v$I2P_7810_out0 && v$NEXTINTERRUPT_17397_out0;
assign v$G1_7538_out0 = v$I2P_7811_out0 && v$NEXTINTERRUPT_17398_out0;
assign v$G2_8647_out0 = v$I3P_11324_out0 && v$NEXTINTERRUPT_17397_out0;
assign v$G2_8648_out0 = v$I3P_11325_out0 && v$NEXTINTERRUPT_17398_out0;
assign v$G3_10364_out0 = v$INITIAL$FETCH$OCCURRED_1691_out0 && v$G27_12276_out0;
assign v$G3_10365_out0 = v$INITIAL$FETCH$OCCURRED_1692_out0 && v$G27_12277_out0;
assign v$PIPELINEHALT_15423_out0 = v$STALL_12797_out0;
assign v$PIPELINEHALT_15424_out0 = v$STALL_12798_out0;
assign v$G4_16044_out0 = v$I1P_2710_out0 && v$NEXTINTERRUPT_17397_out0;
assign v$G4_16045_out0 = v$I1P_2711_out0 && v$NEXTINTERRUPT_17398_out0;
assign v$G6_16152_out0 = ! v$R_18937_out0;
assign v$G6_16155_out0 = ! v$R_18940_out0;
assign v$G6_16163_out0 = ! v$R_18948_out0;
assign v$G6_16166_out0 = ! v$R_18951_out0;
assign v$G19_16478_out0 = v$G21_15317_out0 || v$G6_8265_out0;
assign v$G19_16479_out0 = v$G21_15318_out0 || v$G6_8266_out0;
assign v$G32_16950_out0 = v$G31_2537_out0 && v$IR2$VALID_16482_out0;
assign v$G32_16951_out0 = v$G31_2538_out0 && v$IR2$VALID_16483_out0;
assign v$S_17538_out0 = v$ENABLEINTERRUPTS_13141_out0;
assign v$S_17549_out0 = v$ENABLEINTERRUPTS_13142_out0;
assign v$G9_17559_out0 = v$G28_9040_out0 && v$G10_15189_out0;
assign v$G9_17560_out0 = v$G28_9041_out0 && v$G10_15190_out0;
assign v$SetError_18196_out0 = v$G4_5116_out0;
assign v$SetError_18197_out0 = v$G4_5117_out0;
assign v$G7_1653_out0 = v$G19_16478_out0 && v$IR2$VALID_16482_out0;
assign v$G7_1654_out0 = v$G19_16479_out0 && v$IR2$VALID_16483_out0;
assign v$G9_2724_out0 = v$CLR_4601_out0 || v$G4_16044_out0;
assign v$G9_2725_out0 = v$CLR_4602_out0 || v$G4_16045_out0;
assign v$G11_3223_out0 = v$CLR_4601_out0 || v$G2_8647_out0;
assign v$G11_3224_out0 = v$CLR_4602_out0 || v$G2_8648_out0;
assign v$G10_6926_out0 = v$CLR_4601_out0 || v$G1_7537_out0;
assign v$G10_6927_out0 = v$CLR_4602_out0 || v$G1_7538_out0;
assign v$G13_8221_out0 = v$G9_17559_out0 && v$IR2$IS$FPU_12415_out0;
assign v$G13_8222_out0 = v$G9_17560_out0 && v$IR2$IS$FPU_12416_out0;
assign v$SHOULD$STORE_13280_out0 = v$G32_16950_out0;
assign v$SHOULD$STORE_13281_out0 = v$G32_16951_out0;
assign v$G8_14860_out0 = v$FF2_13616_out0 || v$S_17538_out0;
assign v$G8_14866_out0 = v$FF2_13627_out0 || v$S_17549_out0;
assign v$G8_16068_out0 = v$CLR_4601_out0 || v$G3_4262_out0;
assign v$G8_16069_out0 = v$CLR_4602_out0 || v$G3_4263_out0;
assign v$G14_16418_out0 = v$G8_1401_out0 && v$IR2$IS$FPU_12415_out0;
assign v$G14_16419_out0 = v$G8_1402_out0 && v$IR2$IS$FPU_12416_out0;
assign v$G50_16979_out0 = v$G51_14624_out0 && v$G3_10364_out0;
assign v$G50_16980_out0 = v$G51_14625_out0 && v$G3_10365_out0;
assign v$S_17547_out0 = v$SetError_18196_out0;
assign v$S_17558_out0 = v$SetError_18197_out0;
assign v$G24_249_out0 = v$G7_1653_out0 && v$G26_5343_out0;
assign v$G24_250_out0 = v$G7_1654_out0 && v$G26_5344_out0;
assign v$G33_338_out0 = v$FINISHED_8327_out0 || v$SHOULD$STORE_13280_out0;
assign v$G33_339_out0 = v$FINISHED_8328_out0 || v$SHOULD$STORE_13281_out0;
assign v$G7_14735_out0 = v$G8_14860_out0 && v$G6_16152_out0;
assign v$G7_14741_out0 = v$G8_14866_out0 && v$G6_16163_out0;
assign v$IR1$VALID_18403_out0 = v$G50_16979_out0;
assign v$IR1$VALID_18404_out0 = v$G50_16980_out0;
assign v$R_18936_out0 = v$G8_16068_out0;
assign v$R_18938_out0 = v$G10_6926_out0;
assign v$R_18939_out0 = v$G11_3223_out0;
assign v$R_18941_out0 = v$G9_2724_out0;
assign v$R_18947_out0 = v$G8_16069_out0;
assign v$R_18949_out0 = v$G10_6927_out0;
assign v$R_18950_out0 = v$G11_3224_out0;
assign v$R_18952_out0 = v$G9_2725_out0;
assign v$IR1$VALID_9829_out0 = v$IR1$VALID_18403_out0;
assign v$IR1$VALID_9830_out0 = v$IR1$VALID_18404_out0;
assign v$WENFPU_14322_out0 = v$G24_249_out0;
assign v$WENFPU_14323_out0 = v$G24_250_out0;
assign v$Q_14754_out0 = v$G7_14735_out0;
assign v$Q_14765_out0 = v$G7_14741_out0;
assign v$G6_16151_out0 = ! v$R_18936_out0;
assign v$G6_16153_out0 = ! v$R_18938_out0;
assign v$G6_16154_out0 = ! v$R_18939_out0;
assign v$G6_16156_out0 = ! v$R_18941_out0;
assign v$G6_16162_out0 = ! v$R_18947_out0;
assign v$G6_16164_out0 = ! v$R_18949_out0;
assign v$G6_16165_out0 = ! v$R_18950_out0;
assign v$G6_16167_out0 = ! v$R_18952_out0;
assign v$WENFPU_3698_out0 = v$WENFPU_14322_out0;
assign v$WENFPU_3699_out0 = v$WENFPU_14323_out0;
assign v$IR1$VALID_6037_out0 = v$IR1$VALID_9829_out0;
assign v$IR1$VALID_6038_out0 = v$IR1$VALID_9830_out0;
assign v$ENABLEINTERRUPTS_17620_out0 = v$Q_14754_out0;
assign v$ENABLEINTERRUPTS_17621_out0 = v$Q_14765_out0;
assign v$G19_352_out0 = v$EDGE0_4146_out0 && v$ENABLEINTERRUPTS_17620_out0;
assign v$G19_353_out0 = v$EDGE0_4147_out0 && v$ENABLEINTERRUPTS_17621_out0;
assign v$G22_5098_out0 = v$EDGE3_11552_out0 && v$ENABLEINTERRUPTS_17620_out0;
assign v$G22_5099_out0 = v$EDGE3_11553_out0 && v$ENABLEINTERRUPTS_17621_out0;
assign v$IR1$VALID_14622_out0 = v$IR1$VALID_6037_out0;
assign v$IR1$VALID_14623_out0 = v$IR1$VALID_6038_out0;
assign v$G21_16426_out0 = v$EDGE2_18729_out0 && v$ENABLEINTERRUPTS_17620_out0;
assign v$G21_16427_out0 = v$EDGE2_18730_out0 && v$ENABLEINTERRUPTS_17621_out0;
assign v$G20_16542_out0 = v$EDGE1_15855_out0 && v$ENABLEINTERRUPTS_17620_out0;
assign v$G20_16543_out0 = v$EDGE1_15856_out0 && v$ENABLEINTERRUPTS_17621_out0;
assign v$G13_4516_out0 = v$G21_16426_out0 || v$G22_5098_out0;
assign v$G13_4517_out0 = v$G21_16427_out0 || v$G22_5099_out0;
assign v$G24_8223_out0 = v$LASTQ_12666_out0 && v$G21_16426_out0;
assign v$G24_8224_out0 = v$LASTQ_12677_out0 && v$G21_16427_out0;
assign v$G12_12470_out0 = v$G19_352_out0 || v$G20_16542_out0;
assign v$G12_12471_out0 = v$G19_353_out0 || v$G20_16543_out0;
assign v$G26_13237_out0 = v$LASTQ_12664_out0 && v$G19_352_out0;
assign v$G26_13238_out0 = v$LASTQ_12675_out0 && v$G19_353_out0;
assign v$G25_13587_out0 = v$LASTQ_12669_out0 && v$G20_16542_out0;
assign v$G25_13588_out0 = v$LASTQ_12680_out0 && v$G20_16543_out0;
assign v$S_17537_out0 = v$G19_352_out0;
assign v$S_17539_out0 = v$G21_16426_out0;
assign v$S_17540_out0 = v$G22_5098_out0;
assign v$S_17542_out0 = v$G20_16542_out0;
assign v$S_17548_out0 = v$G19_353_out0;
assign v$S_17550_out0 = v$G21_16427_out0;
assign v$S_17551_out0 = v$G22_5099_out0;
assign v$S_17553_out0 = v$G20_16543_out0;
assign v$IR1$VALID_19035_out0 = v$IR1$VALID_14622_out0;
assign v$IR1$VALID_19036_out0 = v$IR1$VALID_14623_out0;
assign v$G23_19263_out0 = v$LASTQ_12667_out0 && v$G22_5098_out0;
assign v$G23_19264_out0 = v$LASTQ_12678_out0 && v$G22_5099_out0;
assign v$G6_279_out0 = v$G5_17176_out0 && v$IR1$VALID_19035_out0;
assign v$G6_280_out0 = v$G5_17177_out0 && v$IR1$VALID_19036_out0;
assign v$IR1$VALID_4028_out0 = v$IR1$VALID_19035_out0;
assign v$IR1$VALID_4029_out0 = v$IR1$VALID_19036_out0;
assign v$G23_7274_out0 = v$EQ8_261_out0 && v$IR1$VALID_19035_out0;
assign v$G23_7275_out0 = v$EQ8_262_out0 && v$IR1$VALID_19036_out0;
assign v$G7_10362_out0 = v$IR1$VALID_19035_out0 && v$IS$IR1$FMUL_15879_out0;
assign v$G7_10363_out0 = v$IR1$VALID_19036_out0 && v$IS$IR1$FMUL_15880_out0;
assign v$G8_14859_out0 = v$FF2_13615_out0 || v$S_17537_out0;
assign v$G8_14861_out0 = v$FF2_13617_out0 || v$S_17539_out0;
assign v$G8_14862_out0 = v$FF2_13618_out0 || v$S_17540_out0;
assign v$G8_14864_out0 = v$FF2_13620_out0 || v$S_17542_out0;
assign v$G8_14865_out0 = v$FF2_13626_out0 || v$S_17548_out0;
assign v$G8_14867_out0 = v$FF2_13628_out0 || v$S_17550_out0;
assign v$G8_14868_out0 = v$FF2_13629_out0 || v$S_17551_out0;
assign v$G8_14870_out0 = v$FF2_13631_out0 || v$S_17553_out0;
assign v$G14_15875_out0 = v$G12_12470_out0 || v$G13_4516_out0;
assign v$G14_15876_out0 = v$G12_12471_out0 || v$G13_4517_out0;
assign v$G28_15972_out0 = v$G24_8223_out0 || v$G23_19263_out0;
assign v$G28_15973_out0 = v$G24_8224_out0 || v$G23_19264_out0;
assign v$G27_19099_out0 = v$G26_13237_out0 || v$G25_13587_out0;
assign v$G27_19100_out0 = v$G26_13238_out0 || v$G25_13588_out0;
assign v$IR1$VALID_62_out0 = v$IR1$VALID_4028_out0;
assign v$IR1$VALID_63_out0 = v$IR1$VALID_4029_out0;
assign v$INCOMINGINTERRUPT_2066_out0 = v$G14_15875_out0;
assign v$INCOMINGINTERRUPT_2067_out0 = v$G14_15876_out0;
assign v$MUX9_7977_out0 = v$G6_279_out0 ? v$IR1$D_4378_out0 : v$IR2$D_15090_out0;
assign v$MUX9_7978_out0 = v$G6_280_out0 ? v$IR1$D_4379_out0 : v$IR2$D_15091_out0;
assign v$G8_13076_out0 = v$G10_10725_out0 || v$G6_279_out0;
assign v$G8_13077_out0 = v$G10_10726_out0 || v$G6_280_out0;
assign v$EXEC1$FPU_14256_out0 = v$G7_10362_out0;
assign v$EXEC1$FPU_14257_out0 = v$G7_10363_out0;
assign v$G7_14734_out0 = v$G8_14859_out0 && v$G6_16151_out0;
assign v$G7_14736_out0 = v$G8_14861_out0 && v$G6_16153_out0;
assign v$G7_14737_out0 = v$G8_14862_out0 && v$G6_16154_out0;
assign v$G7_14739_out0 = v$G8_14864_out0 && v$G6_16156_out0;
assign v$G7_14740_out0 = v$G8_14865_out0 && v$G6_16162_out0;
assign v$G7_14742_out0 = v$G8_14867_out0 && v$G6_16164_out0;
assign v$G7_14743_out0 = v$G8_14868_out0 && v$G6_16165_out0;
assign v$G7_14745_out0 = v$G8_14870_out0 && v$G6_16167_out0;
assign v$G29_16375_out0 = v$G27_19099_out0 || v$G28_15972_out0;
assign v$G29_16376_out0 = v$G27_19100_out0 || v$G28_15973_out0;
assign v$INTERRUPTOVERFLOW_2438_out0 = v$G29_16375_out0;
assign v$INTERRUPTOVERFLOW_2439_out0 = v$G29_16376_out0;
assign v$G19_3050_out0 = v$G20_12774_out0 && v$IR1$VALID_62_out0;
assign v$G19_3051_out0 = v$G20_12775_out0 && v$IR1$VALID_63_out0;
assign v$AD1_6891_out0 = v$MUX9_7977_out0;
assign v$AD1_6892_out0 = v$MUX9_7978_out0;
assign v$G13_10681_out0 = v$G8_13076_out0 || v$G23_7274_out0;
assign v$G13_10682_out0 = v$G8_13077_out0 || v$G23_7275_out0;
assign v$EXEC1_10709_out0 = v$EXEC1$FPU_14256_out0;
assign v$EXEC1_10710_out0 = v$EXEC1$FPU_14257_out0;
assign v$G17_12704_out0 = v$INCOMINGINTERRUPT_2066_out0 && v$G18_3199_out0;
assign v$G17_12705_out0 = v$INCOMINGINTERRUPT_2067_out0 && v$G18_3200_out0;
assign v$Q_14753_out0 = v$G7_14734_out0;
assign v$Q_14755_out0 = v$G7_14736_out0;
assign v$Q_14756_out0 = v$G7_14737_out0;
assign v$Q_14758_out0 = v$G7_14739_out0;
assign v$Q_14764_out0 = v$G7_14740_out0;
assign v$Q_14766_out0 = v$G7_14742_out0;
assign v$Q_14767_out0 = v$G7_14743_out0;
assign v$Q_14769_out0 = v$G7_14745_out0;
assign v$G5_15253_out0 = v$IR1$VALID_62_out0 && v$IR1$W_17168_out0;
assign v$G5_15254_out0 = v$IR1$VALID_63_out0 && v$IR1$W_17169_out0;
assign v$G4_16135_out0 = v$G3_14794_out0 && v$IR1$VALID_62_out0;
assign v$G4_16136_out0 = v$G3_14795_out0 && v$IR1$VALID_63_out0;
assign v$MUX10_3816_out0 = v$G13_10681_out0 ? v$IR1$M_13829_out0 : v$IR2$M_13567_out0;
assign v$MUX10_3817_out0 = v$G13_10682_out0 ? v$IR1$M_13830_out0 : v$IR2$M_13568_out0;
assign v$I3_5036_out0 = v$Q_14756_out0;
assign v$I3_5037_out0 = v$Q_14767_out0;
assign v$I1_5106_out0 = v$Q_14758_out0;
assign v$I1_5107_out0 = v$Q_14769_out0;
assign v$NEWINTERRUPT_5672_out0 = v$G17_12704_out0;
assign v$NEWINTERRUPT_5673_out0 = v$G17_12705_out0;
assign v$G16_6632_out0 = v$NEXTINTERRUPT_17397_out0 || v$G17_12704_out0;
assign v$G16_6633_out0 = v$NEXTINTERRUPT_17398_out0 || v$G17_12705_out0;
assign v$G6_7798_out0 = v$Q_14755_out0 || v$Q_14756_out0;
assign v$G6_7799_out0 = v$Q_14766_out0 || v$Q_14767_out0;
assign v$G7_12368_out0 = v$G5_15253_out0 || v$G6_12509_out0;
assign v$G7_12369_out0 = v$G5_15254_out0 || v$G6_12510_out0;
assign v$READ$REQUEST_15062_out0 = v$G19_3050_out0;
assign v$READ$REQUEST_15063_out0 = v$G19_3051_out0;
assign v$I2_15092_out0 = v$Q_14755_out0;
assign v$I2_15093_out0 = v$Q_14766_out0;
assign v$G11_15185_out0 = v$G4_16135_out0 && v$G10_15507_out0;
assign v$G11_15186_out0 = v$G4_16136_out0 && v$G10_15508_out0;
assign v$G23_16554_out0 = v$EXEC1_10709_out0 && v$EQ7_14178_out0;
assign v$G23_16555_out0 = v$EXEC1_10710_out0 && v$EQ7_14179_out0;
assign v$G5_16731_out0 = v$Q_14753_out0 || v$Q_14758_out0;
assign v$G5_16732_out0 = v$Q_14764_out0 || v$Q_14769_out0;
assign v$S_17541_out0 = v$INTERRUPTOVERFLOW_2438_out0;
assign v$S_17552_out0 = v$INTERRUPTOVERFLOW_2439_out0;
assign v$I0_19117_out0 = v$Q_14753_out0;
assign v$I0_19118_out0 = v$Q_14764_out0;
assign v$AD1_19284_out0 = v$AD1_6891_out0;
assign v$AD1_19285_out0 = v$AD1_6892_out0;
assign v$CAPTURE_251_out0 = v$G16_6632_out0;
assign v$CAPTURE_252_out0 = v$G16_6633_out0;
assign v$G7_1991_out0 = v$G5_16731_out0 || v$G6_7798_out0;
assign v$G7_1992_out0 = v$G5_16732_out0 || v$G6_7799_out0;
assign v$AD1_2001_out0 = v$AD1_19284_out0;
assign v$AD1_2002_out0 = v$AD1_19285_out0;
assign v$START_3879_out0 = v$G23_16554_out0;
assign v$START_3880_out0 = v$G23_16555_out0;
assign v$NEWINTERRUPT_7309_out0 = v$NEWINTERRUPT_5672_out0;
assign v$NEWINTERRUPT_7310_out0 = v$NEWINTERRUPT_5673_out0;
assign v$G4_8057_out0 = ! v$I1_5106_out0;
assign v$G4_8058_out0 = ! v$I1_5107_out0;
assign v$RAMWEN_8084_out0 = v$G11_15185_out0;
assign v$RAMWEN_8085_out0 = v$G11_15186_out0;
assign v$G2_8098_out0 = ! v$I3_5036_out0;
assign v$G2_8099_out0 = ! v$I3_5037_out0;
assign v$G3_9167_out0 = ! v$I2_15092_out0;
assign v$G3_9168_out0 = ! v$I2_15093_out0;
assign v$AD2_9422_out0 = v$MUX10_3816_out0;
assign v$AD2_9423_out0 = v$MUX10_3817_out0;
assign v$WENLDST_13078_out0 = v$G7_12368_out0;
assign v$WENLDST_13079_out0 = v$G7_12369_out0;
assign v$I3P_14197_out0 = v$I3_5036_out0;
assign v$I3P_14198_out0 = v$I3_5037_out0;
assign v$G8_14863_out0 = v$FF2_13619_out0 || v$S_17541_out0;
assign v$G8_14869_out0 = v$FF2_13630_out0 || v$S_17552_out0;
assign v$READ$REQUEST_17172_out0 = v$READ$REQUEST_15062_out0;
assign v$READ$REQUEST_17173_out0 = v$READ$REQUEST_15063_out0;
assign v$NEWINTERRUPT_4598_out0 = v$NEWINTERRUPT_7309_out0;
assign v$NEWINTERRUPT_4599_out0 = v$NEWINTERRUPT_7310_out0;
assign v$MUX1_5229_out0 = v$G16_6632_out0 ? v$G7_1991_out0 : v$FF1_13671_out0;
assign v$MUX1_5230_out0 = v$G16_6633_out0 ? v$G7_1992_out0 : v$FF1_13672_out0;
assign v$READ$REQUEST_8130_out0 = v$READ$REQUEST_17172_out0;
assign v$READ$REQUEST_8131_out0 = v$READ$REQUEST_17173_out0;
assign v$G7_11473_out0 = v$I0_19117_out0 && v$G4_8057_out0;
assign v$G7_11474_out0 = v$I0_19118_out0 && v$G4_8058_out0;
assign v$_12643_out0 = v$AD1_2001_out0[0:0];
assign v$_12643_out1 = v$AD1_2001_out0[1:1];
assign v$_12644_out0 = v$AD1_2002_out0[0:0];
assign v$_12644_out1 = v$AD1_2002_out0[1:1];
assign v$G1_14123_out0 = v$I2_15092_out0 && v$G2_8098_out0;
assign v$G1_14124_out0 = v$I2_15093_out0 && v$G2_8099_out0;
assign v$G7_14738_out0 = v$G8_14863_out0 && v$G6_16155_out0;
assign v$G7_14744_out0 = v$G8_14869_out0 && v$G6_16166_out0;
assign v$S_16063_out0 = v$START_3879_out0;
assign v$S_16066_out0 = v$START_3880_out0;
assign v$AD2_16254_out0 = v$AD2_9422_out0;
assign v$AD2_16255_out0 = v$AD2_9423_out0;
assign v$RAMWEN_16256_out0 = v$RAMWEN_8084_out0;
assign v$RAMWEN_16257_out0 = v$RAMWEN_8085_out0;
assign v$G8_18510_out0 = v$G3_9167_out0 && v$G2_8098_out0;
assign v$G8_18511_out0 = v$G3_9168_out0 && v$G2_8099_out0;
assign v$WENLDST_19239_out0 = v$WENLDST_13078_out0;
assign v$WENLDST_19240_out0 = v$WENLDST_13079_out0;
assign v$START_19327_out0 = v$START_3879_out0;
assign v$START_19328_out0 = v$START_3880_out0;
assign v$WENRAM_5184_out0 = v$RAMWEN_16256_out0;
assign v$WENRAM_5185_out0 = v$RAMWEN_16257_out0;
assign v$START_5733_out0 = v$START_19327_out0;
assign v$START_5734_out0 = v$START_19328_out0;
assign v$MUX1_6106_out0 = v$_12643_out0 ? v$REG1_5110_out0 : v$REG0_16864_out0;
assign v$MUX1_6107_out0 = v$_12644_out0 ? v$REG1_5111_out0 : v$REG0_16865_out0;
assign v$AD2_6644_out0 = v$AD2_16254_out0;
assign v$AD2_6645_out0 = v$AD2_16255_out0;
assign v$I2P_6676_out0 = v$G1_14123_out0;
assign v$I2P_6677_out0 = v$G1_14124_out0;
assign v$WENLDST_6924_out0 = v$WENLDST_19239_out0;
assign v$WENLDST_6925_out0 = v$WENLDST_19240_out0;
assign v$S_8336_out0 = v$S_16063_out0;
assign v$S_8339_out0 = v$S_16066_out0;
assign v$G12_10366_out0 = !(v$NEWINTERRUPT_4598_out0 || v$FF1_1539_out0);
assign v$G12_10367_out0 = !(v$NEWINTERRUPT_4599_out0 || v$FF1_1540_out0);
assign v$MUX2_11162_out0 = v$_12643_out0 ? v$REG3_11509_out0 : v$REG2_18120_out0;
assign v$MUX2_11163_out0 = v$_12644_out0 ? v$REG3_11510_out0 : v$REG2_18121_out0;
assign v$ISINTERRUPTED_12544_out0 = v$MUX1_5229_out0;
assign v$ISINTERRUPTED_12545_out0 = v$MUX1_5230_out0;
assign v$G6_12692_out0 = v$G7_11473_out0 && v$G8_18510_out0;
assign v$G6_12693_out0 = v$G7_11474_out0 && v$G8_18511_out0;
assign v$Q_14757_out0 = v$G7_14738_out0;
assign v$Q_14768_out0 = v$G7_14744_out0;
assign v$G9_16121_out0 = v$I1_5106_out0 && v$G8_18510_out0;
assign v$G9_16122_out0 = v$I1_5107_out0 && v$G8_18511_out0;
assign v$READ$REQUEST1_17439_out0 = v$READ$REQUEST_8130_out0;
assign v$READ$REQUEST0_19088_out0 = v$READ$REQUEST_8131_out0;
assign v$ININTERRUPT_1277_out0 = v$ISINTERRUPTED_12544_out0;
assign v$ININTERRUPT_1278_out0 = v$ISINTERRUPTED_12545_out0;
assign v$MUX3_1741_out0 = v$_12643_out1 ? v$MUX2_11162_out0 : v$MUX1_6106_out0;
assign v$MUX3_1742_out0 = v$_12644_out1 ? v$MUX2_11163_out0 : v$MUX1_6107_out0;
assign v$G11_2491_out0 = v$G9_15733_out0 && v$G12_10366_out0;
assign v$G11_2492_out0 = v$G9_15734_out0 && v$G12_10367_out0;
assign v$I0P_2632_out0 = v$G6_12692_out0;
assign v$I0P_2633_out0 = v$G6_12693_out0;
assign v$G11_3188_out0 = v$I2P_6676_out0 || v$I3P_14197_out0;
assign v$G11_3189_out0 = v$I2P_6677_out0 || v$I3P_14198_out0;
assign v$G2_4246_out0 = v$G24_14443_out0 && v$WENLDST_6924_out0;
assign v$G2_4247_out0 = v$G24_14444_out0 && v$WENLDST_6925_out0;
assign v$MUX8_4514_out0 = v$IR2$15_7754_out0 ? v$WENALU_4228_out0 : v$WENLDST_6924_out0;
assign v$MUX8_4515_out0 = v$IR2$15_7755_out0 ? v$WENALU_4229_out0 : v$WENLDST_6925_out0;
assign v$XOR1_5225_out0 = v$AD3_13721_out0 ^ v$AD2_6644_out0;
assign v$XOR1_5226_out0 = v$AD3_13722_out0 ^ v$AD2_6645_out0;
assign v$READ$REQUEST1_6717_out0 = v$READ$REQUEST1_17439_out0;
assign v$_7560_out0 = v$AD2_6644_out0[0:0];
assign v$_7560_out1 = v$AD2_6644_out0[1:1];
assign v$_7561_out0 = v$AD2_6645_out0[0:0];
assign v$_7561_out1 = v$AD2_6645_out0[1:1];
assign v$G2_7900_out0 = v$G1_13555_out0 || v$S_8336_out0;
assign v$G2_7903_out0 = v$G1_13558_out0 || v$S_8339_out0;
assign v$READ$REQUEST0_11924_out0 = v$READ$REQUEST0_19088_out0;
assign v$I1P_15425_out0 = v$G9_16121_out0;
assign v$I1P_15426_out0 = v$G9_16122_out0;
assign v$INTERRUPTOVERFLOW_15719_out0 = v$Q_14757_out0;
assign v$INTERRUPTOVERFLOW_15720_out0 = v$Q_14768_out0;
assign v$MUX15_16530_out0 = v$START_5733_out0 ? v$IS$32$BITS_14649_out0 : v$FF1_4502_out0;
assign v$MUX15_16531_out0 = v$START_5734_out0 ? v$IS$32$BITS_14650_out0 : v$FF1_4503_out0;
assign v$START_16968_out0 = v$START_5733_out0;
assign v$START_16969_out0 = v$START_5734_out0;
assign v$WENRAM_17680_out0 = v$WENRAM_5184_out0;
assign v$WENRAM_17681_out0 = v$WENRAM_5185_out0;
assign v$G3_0_out0 = v$G2_4246_out0 && v$IR1$VALID_19035_out0;
assign v$G3_1_out0 = v$G2_4247_out0 && v$IR1$VALID_19036_out0;
assign v$MUX4_1809_out0 = v$_7560_out0 ? v$R1_14351_out0 : v$R0_3503_out0;
assign v$MUX4_1810_out0 = v$_7561_out0 ? v$R1_14352_out0 : v$R0_3504_out0;
assign v$WENRAM_2535_out0 = v$WENRAM_17680_out0;
assign v$WENRAM_2536_out0 = v$WENRAM_17681_out0;
assign v$IS$32$BITS_3203_out0 = v$MUX15_16530_out0;
assign v$IS$32$BITS_3204_out0 = v$MUX15_16531_out0;
assign v$DOUT1_3375_out0 = v$MUX3_1741_out0;
assign v$DOUT1_3376_out0 = v$MUX3_1742_out0;
assign v$EQ1_3433_out0 = v$XOR1_5225_out0 == 2'h0;
assign v$EQ1_3434_out0 = v$XOR1_5226_out0 == 2'h0;
assign v$G10_3985_out0 = v$I1P_15425_out0 || v$I3P_14197_out0;
assign v$G10_3986_out0 = v$I1P_15426_out0 || v$I3P_14198_out0;
assign v$START_4398_out0 = v$START_16968_out0;
assign v$START_4399_out0 = v$START_16969_out0;
assign v$G14_5346_out0 = ! v$ININTERRUPT_1277_out0;
assign v$G14_5347_out0 = ! v$ININTERRUPT_1278_out0;
assign v$G52_8213_out0 = v$READ$REQUEST0_11924_out0 || v$FF2_14043_out0;
assign v$G44_8561_out0 = v$READ$REQUEST1_6717_out0 || v$FF1_5688_out0;
assign v$ARR1_9395_out0 = v$READ$REQUEST1_6717_out0;
assign v$ENCODED1_9898_out0 = v$G11_3188_out0;
assign v$ENCODED1_9899_out0 = v$G11_3189_out0;
assign v$G31_11288_out0 = v$NEXTINTERRUPT_19041_out0 && v$ININTERRUPT_1277_out0;
assign v$G31_11289_out0 = v$NEXTINTERRUPT_19042_out0 && v$ININTERRUPT_1278_out0;
assign v$ARR0_11485_out0 = v$READ$REQUEST0_11924_out0;
assign v$MUX5_12419_out0 = v$EQ1_19203_out0 ? v$WENFPU_3698_out0 : v$MUX8_4514_out0;
assign v$MUX5_12420_out0 = v$EQ1_19204_out0 ? v$WENFPU_3699_out0 : v$MUX8_4515_out0;
assign v$WEN_12738_out0 = v$WENRAM_17680_out0;
assign v$WEN_12739_out0 = v$WENRAM_17681_out0;
assign v$NEXTSTATE_14111_out0 = v$G2_7900_out0;
assign v$NEXTSTATE_14114_out0 = v$G2_7903_out0;
assign v$MUX5_14693_out0 = v$_7560_out0 ? v$R3_11234_out0 : v$R2_8285_out0;
assign v$MUX5_14694_out0 = v$_7561_out0 ? v$R3_11235_out0 : v$R2_8286_out0;
assign v$WEN_14820_out0 = v$WENRAM_17680_out0;
assign v$WEN_14821_out0 = v$WENRAM_17681_out0;
assign v$INTOVERFLOW_16653_out0 = v$INTERRUPTOVERFLOW_15719_out0;
assign v$INTOVERFLOW_16654_out0 = v$INTERRUPTOVERFLOW_15720_out0;
assign v$STPHALT_18735_out0 = v$G11_2491_out0;
assign v$STPHALT_18736_out0 = v$G11_2492_out0;
assign v$WENRAM1_1879_out0 = v$WENRAM_2535_out0;
assign v$RR1_2111_out0 = v$G44_8561_out0;
assign v$RD_2432_out0 = v$DOUT1_3375_out0;
assign v$RD_2433_out0 = v$DOUT1_3376_out0;
assign v$WEN_3862_out0 = v$WEN_14820_out0;
assign v$WEN_3863_out0 = v$WEN_14821_out0;
assign v$WEN_3983_out0 = v$WEN_12738_out0;
assign v$WEN_3984_out0 = v$WEN_12739_out0;
assign v$STPHALT_4478_out0 = v$STPHALT_18735_out0;
assign v$STPHALT_4479_out0 = v$STPHALT_18736_out0;
assign v$MUX6_5267_out0 = v$_7560_out1 ? v$MUX5_14693_out0 : v$MUX4_1809_out0;
assign v$MUX6_5268_out0 = v$_7561_out1 ? v$MUX5_14694_out0 : v$MUX4_1810_out0;
assign v$G29_8174_out0 = v$NEWINTERRUPT_7309_out0 || v$G31_11288_out0;
assign v$G29_8175_out0 = v$NEWINTERRUPT_7310_out0 || v$G31_11289_out0;
assign v$RR0_8403_out0 = v$G52_8213_out0;
assign v$WENRAM0_10341_out0 = v$WENRAM_2536_out0;
assign v$G33_11239_out0 = v$LDMAIN_14395_out0 || v$G14_5346_out0;
assign v$G33_11240_out0 = v$LDMAIN_14396_out0 || v$G14_5347_out0;
assign v$MUX7_11471_out0 = v$IR2$VALID$AND$NOT$FLOAD_7603_out0 ? v$MUX5_12419_out0 : v$G3_0_out0;
assign v$MUX7_11472_out0 = v$IR2$VALID$AND$NOT$FLOAD_7604_out0 ? v$MUX5_12420_out0 : v$G3_1_out0;
assign v$START_14620_out0 = v$START_4398_out0;
assign v$START_14621_out0 = v$START_4399_out0;
assign v$ENCODED0_14632_out0 = v$G10_3985_out0;
assign v$ENCODED0_14633_out0 = v$G10_3986_out0;
assign v$AD3$EQUALS$AD2_15156_out0 = v$EQ1_3433_out0;
assign v$AD3$EQUALS$AD2_15157_out0 = v$EQ1_3434_out0;
assign v$OP1_15807_out0 = v$DOUT1_3375_out0;
assign v$OP1_15808_out0 = v$DOUT1_3376_out0;
assign v$IS$32$BITS_18206_out0 = v$IS$32$BITS_3203_out0;
assign v$IS$32$BITS_18207_out0 = v$IS$32$BITS_3204_out0;
assign v$DOUT2_3714_out0 = v$MUX6_5267_out0;
assign v$DOUT2_3715_out0 = v$MUX6_5268_out0;
assign v$IS$32$BITS_4307_out0 = v$IS$32$BITS_18206_out0;
assign v$IS$32$BITS_4308_out0 = v$IS$32$BITS_18207_out0;
assign v$OP1_5658_out0 = v$OP1_15807_out0;
assign v$OP1_5659_out0 = v$OP1_15808_out0;
assign v$A_9044_out0 = v$RD_2432_out0;
assign v$A_9045_out0 = v$RD_2433_out0;
assign v$MUX15_9777_out0 = v$FINISHED_14451_out0 ? v$WENFPU_3698_out0 : v$MUX7_11471_out0;
assign v$MUX15_9778_out0 = v$FINISHED_14452_out0 ? v$WENFPU_3699_out0 : v$MUX7_11472_out0;
assign v$RDOUT_10807_out0 = v$RD_2432_out0;
assign v$RDOUT_10808_out0 = v$RD_2433_out0;
assign v$RAMWEN1_11257_out0 = v$WENRAM1_1879_out0;
assign v$WEN_12900_out0 = v$WEN_3983_out0;
assign v$WEN_12901_out0 = v$WEN_3984_out0;
assign v$_15215_out0 = { v$ENCODED0_14632_out0,v$ENCODED1_9898_out0 };
assign v$_15216_out0 = { v$ENCODED0_14633_out0,v$ENCODED1_9899_out0 };
assign v$S_16062_out0 = v$START_14620_out0;
assign v$S_16065_out0 = v$START_14621_out0;
assign v$RAMWEN0_17189_out0 = v$WENRAM0_10341_out0;
assign v$INTERRUPTNUMBER_40_out0 = v$_15215_out0;
assign v$INTERRUPTNUMBER_41_out0 = v$_15216_out0;
assign v$AWR0_1960_out0 = v$RAMWEN0_17189_out0;
assign v$WEN3_3509_out0 = v$MUX15_9777_out0;
assign v$WEN3_3510_out0 = v$MUX15_9778_out0;
assign v$DATA$IN_7364_out0 = v$RDOUT_10807_out0;
assign v$DATA$IN_7365_out0 = v$RDOUT_10808_out0;
assign v$S_8335_out0 = v$S_16062_out0;
assign v$S_8338_out0 = v$S_16065_out0;
assign v$A_11554_out0 = v$A_9044_out0;
assign v$A_11555_out0 = v$A_9045_out0;
assign v$G55_14278_out0 = v$RAMWEN0_17189_out0 || v$FF3_3598_out0;
assign v$AWR1_16492_out0 = v$RAMWEN1_11257_out0;
assign v$RM_16803_out0 = v$DOUT2_3714_out0;
assign v$RM_16804_out0 = v$DOUT2_3715_out0;
assign v$A_17040_out0 = v$OP1_5658_out0;
assign v$A_17041_out0 = v$OP1_5659_out0;
assign v$G56_18278_out0 = v$RAMWEN1_11257_out0 || v$FF4_14125_out0;
assign v$WEN_18998_out0 = v$WEN_12900_out0;
assign v$WEN_18999_out0 = v$WEN_12901_out0;
assign v$RM_19205_out0 = v$DOUT2_3714_out0;
assign v$RM_19206_out0 = v$DOUT2_3715_out0;
assign v$WR1_315_out0 = v$G56_18278_out0;
assign v$G6_730_out0 = ! v$WEN_18998_out0;
assign v$G6_731_out0 = ! v$WEN_18999_out0;
assign v$G84_1386_out0 = v$AWR1_16492_out0 || v$ARR1_9395_out0;
assign v$NINTERRUPT_1752_out0 = v$INTERRUPTNUMBER_40_out0;
assign v$NINTERRUPT_1753_out0 = v$INTERRUPTNUMBER_41_out0;
assign v$DATA$IN_1763_out0 = v$DATA$IN_7364_out0;
assign v$DATA$IN_1764_out0 = v$DATA$IN_7365_out0;
assign v$MUX1_1973_out0 = v$C_6338_out0 ? v$_12795_out0 : v$RM_16803_out0;
assign v$MUX1_1974_out0 = v$C_6339_out0 ? v$_12796_out0 : v$RM_16804_out0;
assign v$A_2743_out0 = v$A_17040_out0;
assign v$A_2744_out0 = v$A_17041_out0;
assign v$MUX13_2745_out0 = v$B$IS$RD_14695_out0 ? v$RD_2432_out0 : v$RM_19205_out0;
assign v$MUX13_2746_out0 = v$B$IS$RD_14696_out0 ? v$RD_2433_out0 : v$RM_19206_out0;
assign v$A_4354_out0 = v$A_11554_out0;
assign v$A_4355_out0 = v$A_11555_out0;
assign v$RAMDIN_7323_out0 = v$DATA$IN_7364_out0;
assign v$RAMDIN_7324_out0 = v$DATA$IN_7365_out0;
assign v$G88_7716_out0 = v$ARR0_11485_out0 || v$AWR0_1960_out0;
assign v$G2_7899_out0 = v$G1_13554_out0 || v$S_8335_out0;
assign v$G2_7902_out0 = v$G1_13557_out0 || v$S_8338_out0;
assign v$RM_10695_out0 = v$RM_19205_out0;
assign v$RM_10696_out0 = v$RM_19206_out0;
assign v$G8_13988_out0 = ! v$WEN_18998_out0;
assign v$G8_13989_out0 = ! v$WEN_18999_out0;
assign v$DATA_14697_out0 = v$DATA$IN_7364_out0;
assign v$DATA_14698_out0 = v$DATA$IN_7365_out0;
assign v$D1_14709_out0 = (v$AD3_13721_out0 == 2'b00) ? v$WEN3_3509_out0 : 1'h0;
assign v$D1_14709_out1 = (v$AD3_13721_out0 == 2'b01) ? v$WEN3_3509_out0 : 1'h0;
assign v$D1_14709_out2 = (v$AD3_13721_out0 == 2'b10) ? v$WEN3_3509_out0 : 1'h0;
assign v$D1_14709_out3 = (v$AD3_13721_out0 == 2'b11) ? v$WEN3_3509_out0 : 1'h0;
assign v$D1_14710_out0 = (v$AD3_13722_out0 == 2'b00) ? v$WEN3_3510_out0 : 1'h0;
assign v$D1_14710_out1 = (v$AD3_13722_out0 == 2'b01) ? v$WEN3_3510_out0 : 1'h0;
assign v$D1_14710_out2 = (v$AD3_13722_out0 == 2'b10) ? v$WEN3_3510_out0 : 1'h0;
assign v$D1_14710_out3 = (v$AD3_13722_out0 == 2'b11) ? v$WEN3_3510_out0 : 1'h0;
assign v$WR0_14871_out0 = v$G55_14278_out0;
assign v$A_18897_out0 = v$A_11554_out0;
assign v$A_18898_out0 = v$A_11555_out0;
assign v$IN_196_out0 = v$MUX1_1973_out0;
assign v$IN_197_out0 = v$MUX1_1974_out0;
assign v$_746_out0 = v$A_2743_out0[7:4];
assign v$_747_out0 = v$A_2744_out0[7:4];
assign v$WR0_1478_out0 = v$WR0_14871_out0;
assign v$DIN_1965_out0 = v$RAMDIN_7323_out0;
assign v$DIN_1966_out0 = v$RAMDIN_7324_out0;
assign v$_2012_out0 = { v$A$SAVED_10392_out0,v$A_4354_out0 };
assign v$_2013_out0 = { v$A$SAVED_10393_out0,v$A_4355_out0 };
assign v$A_3465_out0 = v$A_18897_out0;
assign v$A_3466_out0 = v$A_18898_out0;
assign v$_3981_out0 = v$A_2743_out0[15:12];
assign v$_3982_out0 = v$A_2744_out0[15:12];
assign v$_4322_out0 = v$A_2743_out0[3:0];
assign v$_4323_out0 = v$A_2744_out0[3:0];
assign v$DATA_4518_out0 = v$DATA_14697_out0;
assign v$DATA_4519_out0 = v$DATA_14698_out0;
assign v$_9042_out0 = v$A_2743_out0[11:8];
assign v$_9043_out0 = v$A_2744_out0[11:8];
assign v$SEL2_9803_out0 = v$NINTERRUPT_1752_out0[0:0];
assign v$SEL2_9804_out0 = v$NINTERRUPT_1753_out0[0:0];
assign v$DATA$IN0_10855_out0 = v$DATA$IN_1764_out0;
assign v$G79_13307_out0 = v$RR0_8403_out0 || v$WR0_14871_out0;
assign v$NEXTSTATE_14110_out0 = v$G2_7899_out0;
assign v$NEXTSTATE_14113_out0 = v$G2_7902_out0;
assign v$B_14677_out0 = v$MUX13_2745_out0;
assign v$B_14678_out0 = v$MUX13_2746_out0;
assign v$WR1_14940_out0 = v$WR1_315_out0;
assign v$DATA$IN1_15866_out0 = v$DATA$IN_1763_out0;
assign v$G36_17318_out0 = v$RR1_2111_out0 || v$WR1_315_out0;
assign v$SEL3_18044_out0 = v$NINTERRUPT_1752_out0[1:1];
assign v$SEL3_18045_out0 = v$NINTERRUPT_1753_out0[1:1];
assign v$RM_18797_out0 = v$RM_10695_out0;
assign v$RM_18798_out0 = v$RM_10696_out0;
assign v$SEL5_326_out0 = v$A_3465_out0[15:15];
assign v$SEL5_327_out0 = v$A_3466_out0[15:15];
assign v$MUX7_1279_out0 = v$SEL2_9803_out0 ? v$INT3_281_out0 : v$INT2_265_out0;
assign v$MUX7_1280_out0 = v$SEL2_9804_out0 ? v$INT3_282_out0 : v$INT2_266_out0;
assign v$R0_2163_out0 = v$G79_13307_out0;
assign v$PIN_3143_out0 = v$DIN_1965_out0;
assign v$PIN_3144_out0 = v$DIN_1966_out0;
assign v$B_3590_out0 = v$B_14677_out0;
assign v$B_3591_out0 = v$B_14678_out0;
assign v$_3881_out0 = v$_746_out0[1:0];
assign v$_3881_out1 = v$_746_out0[3:2];
assign v$_3882_out0 = v$_747_out0[1:0];
assign v$_3882_out1 = v$_747_out0[3:2];
assign v$IN_4524_out0 = v$IN_196_out0;
assign v$IN_4528_out0 = v$IN_197_out0;
assign v$A_9779_out0 = v$RM_18797_out0;
assign v$A_9780_out0 = v$RM_18798_out0;
assign v$DATAIN1_10016_out0 = v$DATA$IN1_15866_out0;
assign v$SEL9_10394_out0 = v$A_3465_out0[9:0];
assign v$SEL9_10395_out0 = v$A_3466_out0[9:0];
assign v$MUX13_11226_out0 = v$START_5733_out0 ? v$_2012_out0 : v$REG2_4204_out0;
assign v$MUX13_11227_out0 = v$START_5734_out0 ? v$_2013_out0 : v$REG2_4205_out0;
assign v$DATAIN0_11570_out0 = v$DATA$IN0_10855_out0;
assign v$SEL4_12427_out0 = v$DATA_4518_out0[7:0];
assign v$SEL4_12428_out0 = v$DATA_4519_out0[7:0];
assign v$SEL1_12547_out0 = v$DATA_4518_out0[11:0];
assign v$SEL1_12548_out0 = v$DATA_4519_out0[11:0];
assign v$_13839_out0 = v$_9042_out0[1:0];
assign v$_13839_out1 = v$_9042_out0[3:2];
assign v$_13840_out0 = v$_9043_out0[1:0];
assign v$_13840_out1 = v$_9043_out0[3:2];
assign v$A_14399_out0 = v$A_3465_out0;
assign v$A_14403_out0 = v$A_3466_out0;
assign v$MUX6_15024_out0 = v$SEL2_9803_out0 ? v$INT1_19145_out0 : v$INT0_16488_out0;
assign v$MUX6_15025_out0 = v$SEL2_9804_out0 ? v$INT1_19146_out0 : v$INT0_16489_out0;
assign v$_15636_out0 = v$_4322_out0[1:0];
assign v$_15636_out1 = v$_4322_out0[3:2];
assign v$_15637_out0 = v$_4323_out0[1:0];
assign v$_15637_out1 = v$_4323_out0[3:2];
assign v$THRESHOLD_16123_out0 = v$DATA_4518_out0;
assign v$THRESHOLD_16124_out0 = v$DATA_4519_out0;
assign v$SEL11_16147_out0 = v$A_3465_out0[15:15];
assign v$SEL11_16148_out0 = v$A_3466_out0[15:15];
assign v$_16430_out0 = { v$A$SAVED_15235_out0,v$A_3465_out0 };
assign v$_16431_out0 = { v$A$SAVED_15236_out0,v$A_3466_out0 };
assign v$_16841_out0 = v$_3981_out0[1:0];
assign v$_16841_out1 = v$_3981_out0[3:2];
assign v$_16842_out0 = v$_3982_out0[1:0];
assign v$_16842_out1 = v$_3982_out0[3:2];
assign v$SEL13_18204_out0 = v$A_3465_out0[15:15];
assign v$SEL13_18205_out0 = v$A_3466_out0[15:15];
assign v$R1_18512_out0 = v$G36_17318_out0;
assign v$SEL1_18848_out0 = v$DIN_1965_out0[3:0];
assign v$SEL1_18849_out0 = v$DIN_1966_out0[3:0];
assign v$MODE_50_out0 = v$SEL4_12427_out0;
assign v$MODE_51_out0 = v$SEL4_12428_out0;
assign v$_346_out0 = v$_13839_out0[0:0];
assign v$_346_out1 = v$_13839_out0[1:1];
assign v$_347_out0 = v$_13840_out0[0:0];
assign v$_347_out1 = v$_13840_out0[1:1];
assign v$SEL12_1339_out0 = v$MUX13_11226_out0[31:16];
assign v$SEL12_1340_out0 = v$MUX13_11227_out0[31:16];
assign v$_2436_out0 = { v$C8_8515_out0,v$SEL9_10394_out0 };
assign v$_2437_out0 = { v$C8_8516_out0,v$SEL9_10395_out0 };
assign v$G59_2763_out0 = v$PHALT_15747_out0 && v$R1_18512_out0;
assign v$A$32BIT_3201_out0 = v$_16430_out0;
assign v$A$32BIT_3202_out0 = v$_16431_out0;
assign v$_3332_out0 = v$_16841_out1[0:0];
assign v$_3332_out1 = v$_16841_out1[1:1];
assign v$_3333_out0 = v$_16842_out1[0:0];
assign v$_3333_out1 = v$_16842_out1[1:1];
assign v$MUX4_4023_out0 = v$G68_15429_out0 ? v$REG10_17089_out0 : v$DATAIN0_11570_out0;
assign v$_4176_out0 = v$_3881_out0[0:0];
assign v$_4176_out1 = v$_3881_out0[1:1];
assign v$_4177_out0 = v$_3882_out0[0:0];
assign v$_4177_out1 = v$_3882_out0[1:1];
assign v$_5108_out0 = v$_13839_out1[0:0];
assign v$_5108_out1 = v$_13839_out1[1:1];
assign v$_5109_out0 = v$_13840_out1[0:0];
assign v$_5109_out1 = v$_13840_out1[1:1];
assign v$_5646_out0 = v$_15636_out1[0:0];
assign v$_5646_out1 = v$_15636_out1[1:1];
assign v$_5647_out0 = v$_15637_out1[0:0];
assign v$_5647_out1 = v$_15637_out1[1:1];
assign {v$A1_6652_out1,v$A1_6652_out0 } = v$XOR1_5297_out0 + v$A_9779_out0 + v$SUBEN_13429_out0;
assign {v$A1_6653_out1,v$A1_6653_out0 } = v$XOR1_5298_out0 + v$A_9780_out0 + v$SUBEN_13430_out0;
assign v$R0_6913_out0 = v$R0_2163_out0;
assign v$SEL1_7850_out0 = v$A_14399_out0[14:10];
assign v$SEL1_7854_out0 = v$A_14403_out0[14:10];
assign v$_8229_out0 = v$PIN_3143_out0[7:0];
assign v$_8229_out1 = v$PIN_3143_out0[15:8];
assign v$_8230_out0 = v$PIN_3144_out0[7:0];
assign v$_8230_out1 = v$PIN_3144_out0[15:8];
assign v$IN_9946_out0 = v$IN_4524_out0;
assign v$IN_9950_out0 = v$IN_4528_out0;
assign v$_10697_out0 = v$_3881_out1[0:0];
assign v$_10697_out1 = v$_3881_out1[1:1];
assign v$_10698_out0 = v$_3882_out1[0:0];
assign v$_10698_out1 = v$_3882_out1[1:1];
assign v$MUX5_11398_out0 = v$G69_16415_out0 ? v$REG11_10004_out0 : v$DATAIN1_10016_out0;
assign v$_11568_out0 = v$_15636_out0[0:0];
assign v$_11568_out1 = v$_15636_out0[1:1];
assign v$_11569_out0 = v$_15637_out0[0:0];
assign v$_11569_out1 = v$_15637_out0[1:1];
assign v$R1_12459_out0 = v$R1_18512_out0;
assign v$G1_15752_out0 = ! v$SEL5_326_out0;
assign v$G1_15753_out0 = ! v$SEL5_327_out0;
assign v$_17170_out0 = v$_16841_out0[0:0];
assign v$_17170_out1 = v$_16841_out0[1:1];
assign v$_17171_out0 = v$_16842_out0[0:0];
assign v$_17171_out1 = v$_16842_out0[1:1];
assign v$A$32$BIT_17442_out0 = v$MUX13_11226_out0;
assign v$A$32$BIT_17443_out0 = v$MUX13_11227_out0;
assign v$MUX5_17586_out0 = v$SEL3_18044_out0 ? v$MUX7_1279_out0 : v$MUX6_15024_out0;
assign v$MUX5_17587_out0 = v$SEL3_18045_out0 ? v$MUX7_1280_out0 : v$MUX6_15025_out0;
assign v$B_17646_out0 = v$B_3590_out0;
assign v$B_17647_out0 = v$B_3591_out0;
assign v$B_18707_out0 = v$B_3590_out0;
assign v$B_18708_out0 = v$B_3591_out0;
assign v$A$EXP_296_out0 = v$SEL1_7850_out0;
assign v$A$EXP_300_out0 = v$SEL1_7854_out0;
assign v$_1345_out0 = v$IN_9946_out0[0:0];
assign v$_1346_out0 = v$IN_9950_out0[0:0];
assign v$A_2497_out0 = v$SEL12_1339_out0;
assign v$A_2498_out0 = v$SEL12_1340_out0;
assign v$G6_3703_out0 = v$R0_6913_out0 && v$R1_12459_out0;
assign v$_5013_out0 = v$IN_9946_out0[14:0];
assign v$_5017_out0 = v$IN_9950_out0[14:0];
assign v$SEL2_6430_out0 = v$B_17646_out0[14:0];
assign v$SEL2_6431_out0 = v$B_17647_out0[14:0];
assign v$_7735_out0 = { v$_2436_out0,v$C2_1317_out0 };
assign v$_7736_out0 = { v$_2437_out0,v$C2_1318_out0 };
assign v$8LSB_7934_out0 = v$_8229_out0;
assign v$8LSB_7935_out0 = v$_8230_out0;
assign v$COUT_8603_out0 = v$A1_6652_out1;
assign v$COUT_8604_out0 = v$A1_6653_out1;
assign v$SUM_10759_out0 = v$A1_6652_out0;
assign v$SUM_10760_out0 = v$A1_6653_out0;
assign v$_10868_out0 = v$IN_9946_out0[15:15];
assign v$_10869_out0 = v$IN_9950_out0[15:15];
assign v$EQ1_12187_out0 = v$A$32$BIT_17442_out0 == 32'h0;
assign v$EQ1_12188_out0 = v$A$32$BIT_17443_out0 == 32'h0;
assign v$G62_12543_out0 = v$G59_2763_out0 && v$PCHALT_17182_out0;
assign v$_13118_out0 = { v$B$SAVED_4066_out0,v$B_18707_out0 };
assign v$_13119_out0 = { v$B$SAVED_4067_out0,v$B_18708_out0 };
assign v$END_13282_out0 = v$_8229_out1;
assign v$END_13283_out0 = v$_8230_out1;
assign v$SEL4_13548_out0 = v$A$32BIT_3201_out0[22:0];
assign v$SEL4_13549_out0 = v$A$32BIT_3202_out0[22:0];
assign v$_13853_out0 = v$IN_9946_out0[0:0];
assign v$_13856_out0 = v$IN_9950_out0[0:0];
assign v$A_14400_out0 = v$A$32BIT_3201_out0;
assign v$A_14402_out0 = v$A$32$BIT_17442_out0;
assign v$A_14404_out0 = v$A$32BIT_3202_out0;
assign v$A_14406_out0 = v$A$32$BIT_17443_out0;
assign v$EQ3_14906_out0 = v$A$32$BIT_17442_out0 == 32'h0;
assign v$EQ3_14907_out0 = v$A$32$BIT_17443_out0 == 32'h0;
assign v$SEL6_15060_out0 = v$B_17646_out0[15:15];
assign v$SEL6_15061_out0 = v$B_17647_out0[15:15];
assign v$_15201_out0 = v$IN_9946_out0[15:1];
assign v$_15205_out0 = v$IN_9950_out0[15:1];
assign v$_15237_out0 = v$IN_9946_out0[15:1];
assign v$_15241_out0 = v$IN_9950_out0[15:1];
assign v$_17368_out0 = v$IN_9946_out0[15:1];
assign v$_17372_out0 = v$IN_9950_out0[15:1];
assign v$SEL8_18134_out0 = v$A$32$BIT_17442_out0[22:0];
assign v$SEL8_18135_out0 = v$A$32$BIT_17443_out0[22:0];
assign v$MODE_18452_out0 = v$MODE_50_out0;
assign v$MODE_18453_out0 = v$MODE_51_out0;
assign v$MUX14_1335_out0 = v$START_5733_out0 ? v$_13118_out0 : v$REG1_8170_out0;
assign v$MUX14_1336_out0 = v$START_5734_out0 ? v$_13119_out0 : v$REG1_8171_out0;
assign v$_1629_out0 = { v$C1_8287_out0,v$_5013_out0 };
assign v$_1633_out0 = { v$C1_8291_out0,v$_5017_out0 };
assign v$SEL1_3901_out0 = v$A_2497_out0[15:15];
assign v$SEL1_3902_out0 = v$A_2498_out0[15:15];
assign v$G3_4120_out0 = ! v$SEL6_15060_out0;
assign v$G3_4121_out0 = ! v$SEL6_15061_out0;
assign v$RMN_6420_out0 = v$SUM_10759_out0;
assign v$RMN_6421_out0 = v$SUM_10760_out0;
assign v$SEL1_7851_out0 = v$A_14400_out0[30:23];
assign v$SEL1_7853_out0 = v$A_14402_out0[30:23];
assign v$SEL1_7855_out0 = v$A_14404_out0[30:23];
assign v$SEL1_7857_out0 = v$A_14406_out0[30:23];
assign v$_8521_out0 = v$8LSB_7934_out0[3:0];
assign v$_8521_out1 = v$8LSB_7934_out0[7:4];
assign v$_8522_out0 = v$8LSB_7935_out0[3:0];
assign v$_8522_out1 = v$8LSB_7935_out0[7:4];
assign v$_9819_out0 = { v$_17368_out0,v$LSB_8138_out0 };
assign v$_9823_out0 = { v$_17372_out0,v$LSB_8139_out0 };
assign v$MODE_11296_out0 = v$MODE_18452_out0;
assign v$MODE_11297_out0 = v$MODE_18453_out0;
assign v$A_11864_out0 = v$A$EXP_296_out0;
assign v$A_11880_out0 = v$A$EXP_300_out0;
assign v$SEL7_13070_out0 = v$A_2497_out0[9:0];
assign v$SEL7_13071_out0 = v$A_2498_out0[9:0];
assign v$HALTVALID_13870_out0 = v$G6_3703_out0;
assign v$_13890_out0 = { v$_15201_out0,v$_13853_out0 };
assign v$_13894_out0 = { v$_15205_out0,v$_13856_out0 };
assign v$MUX6_14320_out0 = v$S$FF_11312_out0 ? v$LSB_8138_out0 : v$_10868_out0;
assign v$MUX6_14321_out0 = v$S$FF_11313_out0 ? v$LSB_8139_out0 : v$_10869_out0;
assign v$A_14401_out0 = v$A_2497_out0;
assign v$A_14405_out0 = v$A_2498_out0;
assign v$DM1_16855_out0 = v$HALTSEL_15349_out0 ? 1'h0 : v$G6_3703_out0;
assign v$DM1_16855_out1 = v$HALTSEL_15349_out0 ? v$G6_3703_out0 : 1'h0;
assign v$HALT_16989_out0 = v$G6_3703_out0;
assign v$MUX5_17662_out0 = v$S_11196_out0 ? v$_1345_out0 : v$C2_2863_out0;
assign v$MUX5_17663_out0 = v$S_11197_out0 ? v$_1346_out0 : v$C2_2864_out0;
assign v$_18382_out0 = { v$SEL4_13548_out0,v$C3_5628_out0 };
assign v$_18383_out0 = { v$SEL4_13549_out0,v$C3_5629_out0 };
assign v$A$EXP_297_out0 = v$SEL1_7851_out0;
assign v$A$EXP_299_out0 = v$SEL1_7853_out0;
assign v$A$EXP_301_out0 = v$SEL1_7855_out0;
assign v$A$EXP_303_out0 = v$SEL1_7857_out0;
assign v$_1843_out0 = { v$C6_1689_out0,v$SEL7_13070_out0 };
assign v$_1844_out0 = { v$C6_1690_out0,v$SEL7_13071_out0 };
assign v$_1855_out0 = v$_8521_out0[1:0];
assign v$_1855_out1 = v$_8521_out0[3:2];
assign v$_1856_out0 = v$_8522_out0[1:0];
assign v$_1856_out1 = v$_8522_out0[3:2];
assign v$MUX1_2798_out0 = v$G15_19147_out0 ? v$RMN_6420_out0 : v$RM_18797_out0;
assign v$MUX1_2799_out0 = v$G15_19148_out0 ? v$RMN_6421_out0 : v$RM_18798_out0;
assign v$SEL11_3883_out0 = v$MUX14_1335_out0[31:16];
assign v$SEL11_3884_out0 = v$MUX14_1336_out0[31:16];
assign v$MUX8_5638_out0 = v$IS$32$BIT_11362_out0 ? v$_18382_out0 : v$_7735_out0;
assign v$MUX8_5639_out0 = v$IS$32$BIT_11363_out0 ? v$_18383_out0 : v$_7736_out0;
assign v$HALT1_7543_out0 = v$DM1_16855_out1;
assign v$SEL4_7658_out0 = v$A_11864_out0[1:1];
assign v$SEL4_7670_out0 = v$A_11880_out0[1:1];
assign v$SEL1_7852_out0 = v$A_14401_out0[14:10];
assign v$SEL1_7856_out0 = v$A_14405_out0[14:10];
assign v$HALTVALID_8061_out0 = v$HALTVALID_13870_out0;
assign v$SEL3_8736_out0 = v$A_11864_out0[2:2];
assign v$SEL3_8748_out0 = v$A_11880_out0[2:2];
assign v$G7_10295_out0 = ! v$DM1_16855_out0;
assign v$HALT0_12252_out0 = v$DM1_16855_out0;
assign v$_12380_out0 = { v$_15237_out0,v$MUX6_14320_out0 };
assign v$_12384_out0 = { v$_15241_out0,v$MUX6_14321_out0 };
assign v$SEL5_13351_out0 = v$A_11864_out0[0:0];
assign v$SEL5_13363_out0 = v$A_11880_out0[0:0];
assign v$_13729_out0 = v$_8521_out1[1:0];
assign v$_13729_out1 = v$_8521_out1[3:2];
assign v$_13730_out0 = v$_8522_out1[1:0];
assign v$_13730_out1 = v$_8522_out1[3:2];
assign v$MUX4_16600_out0 = v$EN_17561_out0 ? v$_1629_out0 : v$IN_9946_out0;
assign v$MUX4_16604_out0 = v$EN_17565_out0 ? v$_1633_out0 : v$IN_9950_out0;
assign v$MUX10_17016_out0 = v$EQ1_16829_out0 ? v$G3_4120_out0 : v$SEL6_15060_out0;
assign v$MUX10_17017_out0 = v$EQ1_16830_out0 ? v$G3_4121_out0 : v$SEL6_15061_out0;
assign v$SEL2_17226_out0 = v$A_11864_out0[3:3];
assign v$SEL2_17238_out0 = v$A_11880_out0[3:3];
assign v$B$32$BIT_18291_out0 = v$MUX14_1335_out0;
assign v$B$32$BIT_18292_out0 = v$MUX14_1336_out0;
assign v$SEL1_18649_out0 = v$A_11864_out0[4:4];
assign v$SEL1_18651_out0 = v$A_11880_out0[4:4];
assign v$A$EXP_298_out0 = v$SEL1_7852_out0;
assign v$A$EXP_302_out0 = v$SEL1_7856_out0;
assign v$HALT0_380_out0 = v$HALT0_12252_out0;
assign v$_1649_out0 = { v$SEL2_6430_out0,v$MUX10_17016_out0 };
assign v$_1650_out0 = { v$SEL2_6431_out0,v$MUX10_17017_out0 };
assign v$A0_1891_out0 = v$SEL5_13351_out0;
assign v$A0_1903_out0 = v$SEL5_13363_out0;
assign v$EQ4_3217_out0 = v$B$32$BIT_18291_out0 == 32'h0;
assign v$EQ4_3218_out0 = v$B$32$BIT_18292_out0 == 32'h0;
assign v$_3685_out0 = v$_1855_out0[0:0];
assign v$_3685_out1 = v$_1855_out0[1:1];
assign v$_3686_out0 = v$_1856_out0[0:0];
assign v$_3686_out1 = v$_1856_out0[1:1];
assign v$A$MANTISA_3937_out0 = v$MUX8_5638_out0;
assign v$A$MANTISA_3938_out0 = v$MUX8_5639_out0;
assign v$HALT1_4317_out0 = v$HALT1_7543_out0;
assign v$SEL6_4609_out0 = v$B$32$BIT_18291_out0[22:0];
assign v$SEL6_4610_out0 = v$B$32$BIT_18292_out0[22:0];
assign v$B_5041_out0 = v$B$32$BIT_18291_out0;
assign v$B_5045_out0 = v$B$32$BIT_18292_out0;
assign v$B_6781_out0 = v$SEL11_3883_out0;
assign v$B_6782_out0 = v$SEL11_3884_out0;
assign v$MUX8_7366_out0 = v$IS$32$BITS_3203_out0 ? v$SEL8_18134_out0 : v$_1843_out0;
assign v$MUX8_7367_out0 = v$IS$32$BITS_3204_out0 ? v$SEL8_18135_out0 : v$_1844_out0;
assign v$A2_8377_out0 = v$SEL3_8736_out0;
assign v$A2_8389_out0 = v$SEL3_8748_out0;
assign v$_8404_out0 = v$_13729_out0[0:0];
assign v$_8404_out1 = v$_13729_out0[1:1];
assign v$_8405_out0 = v$_13730_out0[0:0];
assign v$_8405_out1 = v$_13730_out0[1:1];
assign v$_9743_out0 = v$_13729_out1[0:0];
assign v$_9743_out1 = v$_13729_out1[1:1];
assign v$_9744_out0 = v$_13730_out1[0:0];
assign v$_9744_out1 = v$_13730_out1[1:1];
assign v$A3_11206_out0 = v$SEL2_17226_out0;
assign v$A3_11218_out0 = v$SEL2_17238_out0;
assign v$A_11865_out0 = v$A$EXP_297_out0;
assign v$A_11869_out0 = v$A$EXP_299_out0;
assign v$A_11881_out0 = v$A$EXP_301_out0;
assign v$A_11885_out0 = v$A$EXP_303_out0;
assign v$MUX2_12603_out0 = v$G3_2800_out0 ? v$_9819_out0 : v$MUX4_16600_out0;
assign v$MUX2_12607_out0 = v$G3_2804_out0 ? v$_9823_out0 : v$MUX4_16604_out0;
assign v$_14634_out0 = v$MUX1_2798_out0[11:0];
assign v$_14634_out1 = v$MUX1_2798_out0[15:4];
assign v$_14635_out0 = v$MUX1_2799_out0[11:0];
assign v$_14635_out1 = v$MUX1_2799_out0[15:4];
assign v$_14689_out0 = v$_1855_out1[0:0];
assign v$_14689_out1 = v$_1855_out1[1:1];
assign v$_14690_out0 = v$_1856_out1[0:0];
assign v$_14690_out1 = v$_1856_out1[1:1];
assign v$A1_14949_out0 = v$SEL4_7658_out0;
assign v$A1_14961_out0 = v$SEL4_7670_out0;
assign v$A4_15624_out0 = v$SEL1_18649_out0;
assign v$A4_15626_out0 = v$SEL1_18651_out0;
assign v$G8_16329_out0 = v$G7_10295_out0 && v$DM1_16855_out1;
assign v$EQ2_16766_out0 = v$B$32$BIT_18291_out0 == 32'h0;
assign v$EQ2_16767_out0 = v$B$32$BIT_18292_out0 == 32'h0;
assign v$HALT1_3317_out0 = v$HALT1_4317_out0;
assign v$B_5040_out0 = v$B_6781_out0;
assign v$B_5044_out0 = v$B_6782_out0;
assign v$HALT0_6091_out0 = v$HALT0_380_out0;
assign v$G72_6179_out0 = ! v$HALT0_380_out0;
assign v$G5_6460_out0 = v$EQ3_14906_out0 || v$EQ4_3217_out0;
assign v$G5_6461_out0 = v$EQ3_14907_out0 || v$EQ4_3218_out0;
assign v$MUX1_6914_out0 = v$G4_4186_out0 ? v$_12380_out0 : v$MUX2_12603_out0;
assign v$MUX1_6918_out0 = v$G4_4190_out0 ? v$_12384_out0 : v$MUX2_12607_out0;
assign v$SEL2_7253_out0 = v$B_5041_out0[30:23];
assign v$SEL2_7257_out0 = v$B_5045_out0[30:23];
assign v$G78_7386_out0 = ! v$HALT1_4317_out0;
assign v$SEL5_8136_out0 = v$B_6781_out0[9:0];
assign v$SEL5_8137_out0 = v$B_6782_out0[9:0];
assign v$SEL1_10747_out0 = v$A_11865_out0[3:0];
assign v$SEL1_10748_out0 = v$A_11869_out0[3:0];
assign v$SEL1_10751_out0 = v$A_11881_out0[3:0];
assign v$SEL1_10752_out0 = v$A_11885_out0[3:0];
assign v$A_11868_out0 = v$A$EXP_298_out0;
assign v$A_11884_out0 = v$A$EXP_302_out0;
assign v$A$MANTISA_12397_out0 = v$MUX8_7366_out0;
assign v$A$MANTISA_12398_out0 = v$MUX8_7367_out0;
assign v$A$MANTISSA_13764_out0 = v$A$MANTISA_3937_out0;
assign v$A$MANTISSA_13765_out0 = v$A$MANTISA_3938_out0;
assign v$G54_13869_out0 = v$RAMWEN1_11257_out0 && v$HALT1_4317_out0;
assign v$G50_13889_out0 = ! v$HALT1_4317_out0;
assign v$SEL2_14017_out0 = v$B_6781_out0[15:15];
assign v$SEL2_14018_out0 = v$B_6782_out0[15:15];
assign v$G63_14258_out0 = v$HALT0_380_out0 || v$HALT1_4317_out0;
assign v$HALT0_14750_out0 = v$HALT0_380_out0;
assign v$RAMADDRMUX_14981_out0 = v$_14634_out0;
assign v$RAMADDRMUX_14982_out0 = v$_14635_out0;
assign v$ADDRMSB_15646_out0 = v$_14634_out1;
assign v$ADDRMSB_15647_out0 = v$_14635_out1;
assign v$G45_15949_out0 = v$READ$REQUEST1_6717_out0 && v$HALT1_4317_out0;
assign v$G3_16620_out0 = v$EQ1_12187_out0 || v$EQ2_16766_out0;
assign v$G3_16621_out0 = v$EQ1_12188_out0 || v$EQ2_16767_out0;
assign v$SEL4_17973_out0 = v$A_11865_out0[7:4];
assign v$SEL4_17974_out0 = v$A_11869_out0[7:4];
assign v$SEL4_17977_out0 = v$A_11881_out0[7:4];
assign v$SEL4_17978_out0 = v$A_11885_out0[7:4];
assign v$G53_18133_out0 = v$RAMWEN0_17189_out0 && v$HALT0_380_out0;
assign v$B_18356_out0 = v$_1649_out0;
assign v$B_18357_out0 = v$_1650_out0;
assign v$HALT1_18913_out0 = v$HALT1_4317_out0;
assign v$G51_19373_out0 = v$READ$REQUEST0_11924_out0 && v$HALT0_380_out0;
assign v$SEL12_16_out0 = v$B_18356_out0[9:0];
assign v$SEL12_17_out0 = v$B_18357_out0[9:0];
assign v$SEL3_1405_out0 = v$A$MANTISSA_13764_out0[23:12];
assign v$SEL3_1406_out0 = v$A$MANTISSA_13765_out0[23:12];
assign v$HALT_1449_out0 = v$G63_14258_out0;
assign v$MUX3_2122_out0 = v$G8_2050_out0 ? v$_13890_out0 : v$MUX1_6914_out0;
assign v$MUX3_2126_out0 = v$G8_2054_out0 ? v$_13894_out0 : v$MUX1_6918_out0;
assign v$ARBHALT0_3114_out0 = v$HALT0_6091_out0;
assign v$SEL1_3473_out0 = v$A$MANTISSA_13764_out0[11:0];
assign v$SEL1_3474_out0 = v$A$MANTISSA_13765_out0[11:0];
assign v$RAMADDRMUX_5029_out0 = v$RAMADDRMUX_14981_out0;
assign v$RAMADDRMUX_5030_out0 = v$RAMADDRMUX_14982_out0;
assign v$B_5038_out0 = v$B_18356_out0;
assign v$B_5042_out0 = v$B_18357_out0;
assign v$ARBHALT1_5693_out0 = v$HALT1_3317_out0;
assign v$G64_6675_out0 = v$G50_13889_out0 && v$R1_18512_out0;
assign v$SEL2_7252_out0 = v$B_5040_out0[14:10];
assign v$SEL2_7256_out0 = v$B_5044_out0[14:10];
assign v$G1_7651_out0 = ! v$HALT1_18913_out0;
assign v$SEL4_7661_out0 = v$A_11868_out0[1:1];
assign v$SEL4_7673_out0 = v$A_11884_out0[1:1];
assign v$G2_8434_out0 = ! v$HALT0_14750_out0;
assign v$SEL3_8739_out0 = v$A_11868_out0[2:2];
assign v$SEL3_8751_out0 = v$A_11884_out0[2:2];
assign v$A_11866_out0 = v$SEL4_17973_out0;
assign v$A_11867_out0 = v$SEL1_10747_out0;
assign v$A_11870_out0 = v$SEL4_17974_out0;
assign v$A_11871_out0 = v$SEL1_10748_out0;
assign v$A_11882_out0 = v$SEL4_17977_out0;
assign v$A_11883_out0 = v$SEL1_10751_out0;
assign v$A_11886_out0 = v$SEL4_17978_out0;
assign v$A_11887_out0 = v$SEL1_10752_out0;
assign v$SEL5_13354_out0 = v$A_11868_out0[0:0];
assign v$SEL5_13366_out0 = v$A_11884_out0[0:0];
assign v$SEL15_14189_out0 = v$B_18356_out0[15:15];
assign v$SEL15_14190_out0 = v$B_18357_out0[15:15];
assign v$G74_16338_out0 = v$REG4_11502_out0 && v$G72_6179_out0;
assign v$SEL2_17229_out0 = v$A_11868_out0[3:3];
assign v$SEL2_17241_out0 = v$A_11884_out0[3:3];
assign v$B$EXP_17297_out0 = v$SEL2_7253_out0;
assign v$B$EXP_17301_out0 = v$SEL2_7257_out0;
assign v$G1_18498_out0 = ((v$SEL1_3901_out0 && !v$SEL2_14017_out0) || (!v$SEL1_3901_out0) && v$SEL2_14017_out0);
assign v$G1_18499_out0 = ((v$SEL1_3902_out0 && !v$SEL2_14018_out0) || (!v$SEL1_3902_out0) && v$SEL2_14018_out0);
assign v$A$MANTISA_18529_out0 = v$A$MANTISA_12397_out0;
assign v$A$MANTISA_18530_out0 = v$A$MANTISA_12398_out0;
assign v$SEL1_18650_out0 = v$A_11868_out0[4:4];
assign v$SEL1_18652_out0 = v$A_11884_out0[4:4];
assign v$_18695_out0 = { v$C7_6318_out0,v$SEL5_8136_out0 };
assign v$_18696_out0 = { v$C7_6319_out0,v$SEL5_8137_out0 };
assign v$G77_18811_out0 = v$REG7_6442_out0 && v$G78_7386_out0;
assign v$_18862_out0 = { v$B$SAVED_4522_out0,v$B_18356_out0 };
assign v$_18863_out0 = { v$B$SAVED_4523_out0,v$B_18357_out0 };
assign v$RAMADDRMUX_437_out0 = v$RAMADDRMUX_5029_out0;
assign v$RAMADDRMUX_438_out0 = v$RAMADDRMUX_5030_out0;
assign v$G83_447_out0 = v$G74_16338_out0 && v$G87_5362_out0;
assign v$A0_1894_out0 = v$SEL5_13354_out0;
assign v$A0_1906_out0 = v$SEL5_13366_out0;
assign v$A_2739_out0 = v$SEL3_1405_out0;
assign v$A_2740_out0 = v$SEL1_3473_out0;
assign v$A_2741_out0 = v$SEL3_1406_out0;
assign v$A_2742_out0 = v$SEL1_3474_out0;
assign v$G3_3187_out0 = v$G1_7651_out0 && v$WR1_14940_out0;
assign v$OUT_3397_out0 = v$MUX3_2122_out0;
assign v$OUT_3401_out0 = v$MUX3_2126_out0;
assign v$G85_6462_out0 = v$G77_18811_out0 && v$G86_14102_out0;
assign v$SEL2_7250_out0 = v$B_5038_out0[14:10];
assign v$SEL2_7254_out0 = v$B_5042_out0[14:10];
assign v$SEL4_7659_out0 = v$A_11866_out0[1:1];
assign v$SEL4_7660_out0 = v$A_11867_out0[1:1];
assign v$SEL4_7662_out0 = v$A_11870_out0[1:1];
assign v$SEL4_7663_out0 = v$A_11871_out0[1:1];
assign v$SEL4_7671_out0 = v$A_11882_out0[1:1];
assign v$SEL4_7672_out0 = v$A_11883_out0[1:1];
assign v$SEL4_7674_out0 = v$A_11886_out0[1:1];
assign v$SEL4_7675_out0 = v$A_11887_out0[1:1];
assign v$HALT_7897_out0 = v$ARBHALT1_5693_out0;
assign v$HALT_7898_out0 = v$ARBHALT0_3114_out0;
assign v$A2_8380_out0 = v$SEL3_8739_out0;
assign v$A2_8392_out0 = v$SEL3_8751_out0;
assign v$SEL3_8737_out0 = v$A_11866_out0[2:2];
assign v$SEL3_8738_out0 = v$A_11867_out0[2:2];
assign v$SEL3_8740_out0 = v$A_11870_out0[2:2];
assign v$SEL3_8741_out0 = v$A_11871_out0[2:2];
assign v$SEL3_8749_out0 = v$A_11882_out0[2:2];
assign v$SEL3_8750_out0 = v$A_11883_out0[2:2];
assign v$SEL3_8752_out0 = v$A_11886_out0[2:2];
assign v$SEL3_8753_out0 = v$A_11887_out0[2:2];
assign v$A3_11209_out0 = v$SEL2_17229_out0;
assign v$A3_11221_out0 = v$SEL2_17241_out0;
assign v$MUX7_13312_out0 = v$IS$32$BITS_3203_out0 ? v$SEL6_4609_out0 : v$_18695_out0;
assign v$MUX7_13313_out0 = v$IS$32$BITS_3204_out0 ? v$SEL6_4610_out0 : v$_18696_out0;
assign v$SIGN_13329_out0 = v$G1_18498_out0;
assign v$SIGN_13330_out0 = v$G1_18499_out0;
assign v$SEL5_13352_out0 = v$A_11866_out0[0:0];
assign v$SEL5_13353_out0 = v$A_11867_out0[0:0];
assign v$SEL5_13355_out0 = v$A_11870_out0[0:0];
assign v$SEL5_13356_out0 = v$A_11871_out0[0:0];
assign v$SEL5_13364_out0 = v$A_11882_out0[0:0];
assign v$SEL5_13365_out0 = v$A_11883_out0[0:0];
assign v$SEL5_13367_out0 = v$A_11886_out0[0:0];
assign v$SEL5_13368_out0 = v$A_11887_out0[0:0];
assign v$G4_13766_out0 = v$G2_8434_out0 && v$WR0_1478_out0;
assign v$G6_14205_out0 = ((v$SEL11_16147_out0 && !v$SEL15_14189_out0) || (!v$SEL11_16147_out0) && v$SEL15_14189_out0);
assign v$G6_14206_out0 = ((v$SEL11_16148_out0 && !v$SEL15_14190_out0) || (!v$SEL11_16148_out0) && v$SEL15_14190_out0);
assign v$A1_14952_out0 = v$SEL4_7661_out0;
assign v$A1_14964_out0 = v$SEL4_7673_out0;
assign v$B_15041_out0 = v$B$EXP_17297_out0;
assign v$B_15057_out0 = v$B$EXP_17301_out0;
assign v$A$MANTISA_15148_out0 = v$A$MANTISA_18529_out0;
assign v$A$MANTISA_15149_out0 = v$A$MANTISA_18530_out0;
assign v$A4_15625_out0 = v$SEL1_18650_out0;
assign v$A4_15627_out0 = v$SEL1_18652_out0;
assign v$_16853_out0 = { v$C10_9279_out0,v$SEL12_16_out0 };
assign v$_16854_out0 = { v$C10_9280_out0,v$SEL12_17_out0 };
assign v$SEL2_17227_out0 = v$A_11866_out0[3:3];
assign v$SEL2_17228_out0 = v$A_11867_out0[3:3];
assign v$SEL2_17230_out0 = v$A_11870_out0[3:3];
assign v$SEL2_17231_out0 = v$A_11871_out0[3:3];
assign v$SEL2_17239_out0 = v$A_11882_out0[3:3];
assign v$SEL2_17240_out0 = v$A_11883_out0[3:3];
assign v$SEL2_17242_out0 = v$A_11886_out0[3:3];
assign v$SEL2_17243_out0 = v$A_11887_out0[3:3];
assign v$B$EXP_17296_out0 = v$SEL2_7252_out0;
assign v$B$EXP_17300_out0 = v$SEL2_7256_out0;
assign v$G57_18569_out0 = v$G62_12543_out0 || v$G64_6675_out0;
assign v$B$32BIT_19081_out0 = v$_18862_out0;
assign v$B$32BIT_19082_out0 = v$_18863_out0;
assign v$SIGN_1529_out0 = v$SIGN_13329_out0;
assign v$SIGN_1530_out0 = v$SIGN_13329_out0;
assign v$SIGN_1531_out0 = v$SIGN_13330_out0;
assign v$SIGN_1532_out0 = v$SIGN_13330_out0;
assign v$A0_1892_out0 = v$SEL5_13352_out0;
assign v$A0_1893_out0 = v$SEL5_13353_out0;
assign v$A0_1895_out0 = v$SEL5_13355_out0;
assign v$A0_1896_out0 = v$SEL5_13356_out0;
assign v$A0_1904_out0 = v$SEL5_13364_out0;
assign v$A0_1905_out0 = v$SEL5_13365_out0;
assign v$A0_1907_out0 = v$SEL5_13367_out0;
assign v$A0_1908_out0 = v$SEL5_13368_out0;
assign v$G5_2865_out0 = v$G4_13766_out0 || v$G3_3187_out0;
assign v$HALT_3106_out0 = v$HALT_7897_out0;
assign v$HALT_3107_out0 = v$HALT_7898_out0;
assign v$B$MANTISA_3213_out0 = v$MUX7_13312_out0;
assign v$B$MANTISA_3214_out0 = v$MUX7_13313_out0;
assign v$IN_4525_out0 = v$OUT_3397_out0;
assign v$IN_4529_out0 = v$OUT_3401_out0;
assign v$IS$SUB_4611_out0 = v$G6_14205_out0;
assign v$IS$SUB_4612_out0 = v$G6_14206_out0;
assign v$B_5039_out0 = v$B$32BIT_19081_out0;
assign v$B_5043_out0 = v$B$32BIT_19082_out0;
assign v$SEL8_7593_out0 = v$B$32BIT_19081_out0[22:0];
assign v$SEL8_7594_out0 = v$B$32BIT_19082_out0[22:0];
assign v$G90_8368_out0 = v$PHALT0$PREV_7940_out0 || v$G83_447_out0;
assign v$A2_8378_out0 = v$SEL3_8737_out0;
assign v$A2_8379_out0 = v$SEL3_8738_out0;
assign v$A2_8381_out0 = v$SEL3_8740_out0;
assign v$A2_8382_out0 = v$SEL3_8741_out0;
assign v$A2_8390_out0 = v$SEL3_8749_out0;
assign v$A2_8391_out0 = v$SEL3_8750_out0;
assign v$A2_8393_out0 = v$SEL3_8752_out0;
assign v$A2_8394_out0 = v$SEL3_8753_out0;
assign v$SEL1_8397_out0 = v$A_2739_out0[7:0];
assign v$SEL1_8398_out0 = v$A_2740_out0[7:0];
assign v$SEL1_8399_out0 = v$A_2741_out0[7:0];
assign v$SEL1_8400_out0 = v$A_2742_out0[7:0];
assign v$SEL3_9376_out0 = v$B_15041_out0[7:4];
assign v$SEL3_9380_out0 = v$B_15057_out0[7:4];
assign v$A3_11207_out0 = v$SEL2_17227_out0;
assign v$A3_11208_out0 = v$SEL2_17228_out0;
assign v$A3_11210_out0 = v$SEL2_17230_out0;
assign v$A3_11211_out0 = v$SEL2_17231_out0;
assign v$A3_11219_out0 = v$SEL2_17239_out0;
assign v$A3_11220_out0 = v$SEL2_17240_out0;
assign v$A3_11222_out0 = v$SEL2_17242_out0;
assign v$A3_11223_out0 = v$SEL2_17243_out0;
assign v$SEL3_12468_out0 = v$A$MANTISA_15148_out0[22:0];
assign v$SEL3_12469_out0 = v$A$MANTISA_15149_out0[22:0];
assign v$A1_14950_out0 = v$SEL4_7659_out0;
assign v$A1_14951_out0 = v$SEL4_7660_out0;
assign v$A1_14953_out0 = v$SEL4_7662_out0;
assign v$A1_14954_out0 = v$SEL4_7663_out0;
assign v$A1_14962_out0 = v$SEL4_7671_out0;
assign v$A1_14963_out0 = v$SEL4_7672_out0;
assign v$A1_14965_out0 = v$SEL4_7674_out0;
assign v$A1_14966_out0 = v$SEL4_7675_out0;
assign v$B_15040_out0 = v$B$EXP_17296_out0;
assign v$B_15056_out0 = v$B$EXP_17300_out0;
assign v$RAM$ADDR_15811_out0 = v$RAMADDRMUX_437_out0;
assign v$RAM$ADDR_15812_out0 = v$RAMADDRMUX_438_out0;
assign v$_15937_out0 = { v$_16853_out0,v$C1_16526_out0 };
assign v$_15938_out0 = { v$_16854_out0,v$C1_16527_out0 };
assign v$SEL1_16347_out0 = v$A$MANTISA_15148_out0[22:0];
assign v$SEL1_16348_out0 = v$A$MANTISA_15149_out0[22:0];
assign v$B$EXP_17294_out0 = v$SEL2_7250_out0;
assign v$B$EXP_17298_out0 = v$SEL2_7254_out0;
assign v$SEL2_18085_out0 = v$B_15041_out0[3:0];
assign v$SEL2_18089_out0 = v$B_15057_out0[3:0];
assign v$G89_18384_out0 = v$G85_6462_out0 || v$PHALT1$PREV_7682_out0;
assign v$SELIN_18816_out0 = v$G57_18569_out0;
assign v$SEL3_19229_out0 = v$A_2739_out0[11:8];
assign v$SEL3_19230_out0 = v$A_2740_out0[11:8];
assign v$SEL3_19231_out0 = v$A_2741_out0[11:8];
assign v$SEL3_19232_out0 = v$A_2742_out0[11:8];
assign v$B$MANTISA_4226_out0 = v$B$MANTISA_3213_out0;
assign v$B$MANTISA_4227_out0 = v$B$MANTISA_3214_out0;
assign v$SEL7_4333_out0 = v$B_15040_out0[3:3];
assign v$SEL7_4345_out0 = v$B_15056_out0[3:3];
assign v$SEL6_6093_out0 = v$B_15040_out0[4:4];
assign v$SEL6_6095_out0 = v$B_15056_out0[4:4];
assign v$RAM$ADDR_6656_out0 = v$RAM$ADDR_15811_out0;
assign v$RAM$ADDR_6657_out0 = v$RAM$ADDR_15812_out0;
assign v$SEL2_7251_out0 = v$B_5039_out0[30:23];
assign v$SEL2_7255_out0 = v$B_5043_out0[30:23];
assign v$RAMADDRESS_7270_out0 = v$RAM$ADDR_15811_out0;
assign v$RAMADDRESS_7271_out0 = v$RAM$ADDR_15812_out0;
assign v$V0_7741_out0 = v$G90_8368_out0;
assign v$_7943_out0 = { v$SEL8_7593_out0,v$C6_1725_out0 };
assign v$_7944_out0 = { v$SEL8_7594_out0,v$C6_1726_out0 };
assign v$IN_9947_out0 = v$IN_4525_out0;
assign v$IN_9951_out0 = v$IN_4529_out0;
assign v$SEL9_11345_out0 = v$B_15040_out0[1:1];
assign v$SEL9_11357_out0 = v$B_15056_out0[1:1];
assign v$A_11856_out0 = v$SEL3_19229_out0;
assign v$A_11857_out0 = v$SEL1_8397_out0;
assign v$A_11860_out0 = v$SEL3_19230_out0;
assign v$A_11861_out0 = v$SEL1_8398_out0;
assign v$A_11872_out0 = v$SEL3_19231_out0;
assign v$A_11873_out0 = v$SEL1_8399_out0;
assign v$A_11876_out0 = v$SEL3_19232_out0;
assign v$A_11877_out0 = v$SEL1_8400_out0;
assign v$SEL10_13198_out0 = v$B_15040_out0[0:0];
assign v$SEL10_13210_out0 = v$B_15056_out0[0:0];
assign v$SEL8_13493_out0 = v$B_15040_out0[2:2];
assign v$SEL8_13505_out0 = v$B_15056_out0[2:2];
assign v$B_15036_out0 = v$B$EXP_17294_out0;
assign v$B_15042_out0 = v$SEL3_9376_out0;
assign v$B_15043_out0 = v$SEL2_18085_out0;
assign v$B_15052_out0 = v$B$EXP_17298_out0;
assign v$B_15058_out0 = v$SEL3_9380_out0;
assign v$B_15059_out0 = v$SEL2_18089_out0;
assign v$IS$SUB_16036_out0 = v$IS$SUB_4611_out0;
assign v$IS$SUB_16037_out0 = v$IS$SUB_4612_out0;
assign v$MUX2_16447_out0 = v$SELIN_18816_out0 ? v$MUX5_11398_out0 : v$MUX4_4023_out0;
assign v$ADDRESS_16504_out0 = v$RAM$ADDR_15811_out0;
assign v$ADDRESS_16505_out0 = v$RAM$ADDR_15812_out0;
assign v$V1_17321_out0 = v$G89_18384_out0;
assign v$HALT_18283_out0 = v$HALT_3106_out0;
assign v$HALT_18284_out0 = v$HALT_3107_out0;
assign v$MEMHALT_18405_out0 = v$HALT_3106_out0;
assign v$MEMHALT_18406_out0 = v$HALT_3107_out0;
assign v$MUX5_1767_out0 = v$IS$32$BIT_11362_out0 ? v$_7943_out0 : v$_15937_out0;
assign v$MUX5_1768_out0 = v$IS$32$BIT_11363_out0 ? v$_7944_out0 : v$_15938_out0;
assign v$B0_3845_out0 = v$SEL10_13198_out0;
assign v$B0_3857_out0 = v$SEL10_13210_out0;
assign v$SEL7_4330_out0 = v$B_15036_out0[3:3];
assign v$SEL7_4334_out0 = v$B_15042_out0[3:3];
assign v$SEL7_4335_out0 = v$B_15043_out0[3:3];
assign v$SEL7_4342_out0 = v$B_15052_out0[3:3];
assign v$SEL7_4346_out0 = v$B_15058_out0[3:3];
assign v$SEL7_4347_out0 = v$B_15059_out0[3:3];
assign v$_5014_out0 = v$IN_9947_out0[13:0];
assign v$_5018_out0 = v$IN_9951_out0[13:0];
assign v$B$MANTISA_5124_out0 = v$B$MANTISA_4226_out0;
assign v$B$MANTISA_5125_out0 = v$B$MANTISA_4227_out0;
assign v$SEL6_6092_out0 = v$B_15036_out0[4:4];
assign v$SEL6_6094_out0 = v$B_15052_out0[4:4];
assign v$ADDRESS_6098_out0 = v$ADDRESS_16504_out0;
assign v$ADDRESS_6099_out0 = v$ADDRESS_16505_out0;
assign v$RAM$ADDR1_6700_out0 = v$RAM$ADDR_6656_out0;
assign v$SEL4_7652_out0 = v$A_11856_out0[1:1];
assign v$SEL4_7655_out0 = v$A_11860_out0[1:1];
assign v$SEL4_7664_out0 = v$A_11872_out0[1:1];
assign v$SEL4_7667_out0 = v$A_11876_out0[1:1];
assign v$SEL3_8730_out0 = v$A_11856_out0[2:2];
assign v$SEL3_8733_out0 = v$A_11860_out0[2:2];
assign v$SEL3_8742_out0 = v$A_11872_out0[2:2];
assign v$SEL3_8745_out0 = v$A_11876_out0[2:2];
assign v$VALID1_9151_out0 = v$V1_17321_out0;
assign v$SEL1_10745_out0 = v$A_11857_out0[3:0];
assign v$SEL1_10746_out0 = v$A_11861_out0[3:0];
assign v$SEL1_10749_out0 = v$A_11873_out0[3:0];
assign v$SEL1_10750_out0 = v$A_11877_out0[3:0];
assign v$SEL9_11342_out0 = v$B_15036_out0[1:1];
assign v$SEL9_11346_out0 = v$B_15042_out0[1:1];
assign v$SEL9_11347_out0 = v$B_15043_out0[1:1];
assign v$SEL9_11354_out0 = v$B_15052_out0[1:1];
assign v$SEL9_11358_out0 = v$B_15058_out0[1:1];
assign v$SEL9_11359_out0 = v$B_15059_out0[1:1];
assign v$_12334_out0 = v$IN_9947_out0[15:15];
assign v$_12335_out0 = v$IN_9951_out0[15:15];
assign v$RAM$ADDR0_13120_out0 = v$RAM$ADDR_6657_out0;
assign v$SEL10_13195_out0 = v$B_15036_out0[0:0];
assign v$SEL10_13199_out0 = v$B_15042_out0[0:0];
assign v$SEL10_13200_out0 = v$B_15043_out0[0:0];
assign v$SEL10_13207_out0 = v$B_15052_out0[0:0];
assign v$SEL10_13211_out0 = v$B_15058_out0[0:0];
assign v$SEL10_13212_out0 = v$B_15059_out0[0:0];
assign v$RAMADDRESS_13291_out0 = v$RAMADDRESS_7270_out0;
assign v$RAMADDRESS_13292_out0 = v$RAMADDRESS_7271_out0;
assign v$SEL5_13345_out0 = v$A_11856_out0[0:0];
assign v$SEL5_13348_out0 = v$A_11860_out0[0:0];
assign v$SEL5_13357_out0 = v$A_11872_out0[0:0];
assign v$SEL5_13360_out0 = v$A_11876_out0[0:0];
assign v$HALT_13471_out0 = v$HALT_18283_out0;
assign v$HALT_13472_out0 = v$HALT_18284_out0;
assign v$SEL8_13490_out0 = v$B_15036_out0[2:2];
assign v$SEL8_13494_out0 = v$B_15042_out0[2:2];
assign v$SEL8_13495_out0 = v$B_15043_out0[2:2];
assign v$SEL8_13502_out0 = v$B_15052_out0[2:2];
assign v$SEL8_13506_out0 = v$B_15058_out0[2:2];
assign v$SEL8_13507_out0 = v$B_15059_out0[2:2];
assign v$IS$SUB_13643_out0 = v$IS$SUB_16036_out0;
assign v$IS$SUB_13644_out0 = v$IS$SUB_16037_out0;
assign v$VALID0_13990_out0 = v$V0_7741_out0;
assign v$_14777_out0 = v$IN_9947_out0[1:0];
assign v$_14778_out0 = v$IN_9951_out0[1:0];
assign v$B1_14831_out0 = v$SEL9_11345_out0;
assign v$B1_14843_out0 = v$SEL9_11357_out0;
assign v$_15202_out0 = v$IN_9947_out0[15:2];
assign v$_15206_out0 = v$IN_9951_out0[15:2];
assign v$_15238_out0 = v$IN_9947_out0[15:2];
assign v$_15242_out0 = v$IN_9951_out0[15:2];
assign v$SEL2_17220_out0 = v$A_11856_out0[3:3];
assign v$SEL2_17223_out0 = v$A_11860_out0[3:3];
assign v$SEL2_17232_out0 = v$A_11872_out0[3:3];
assign v$SEL2_17235_out0 = v$A_11876_out0[3:3];
assign v$B2_17253_out0 = v$SEL8_13493_out0;
assign v$B2_17265_out0 = v$SEL8_13505_out0;
assign v$B$EXP_17295_out0 = v$SEL2_7251_out0;
assign v$B$EXP_17299_out0 = v$SEL2_7255_out0;
assign v$_17369_out0 = v$IN_9947_out0[15:2];
assign v$_17373_out0 = v$IN_9951_out0[15:2];
assign v$B4_17534_out0 = v$SEL6_6093_out0;
assign v$B4_17536_out0 = v$SEL6_6095_out0;
assign v$_17652_out0 = v$IN_9947_out0[1:0];
assign v$_17653_out0 = v$IN_9951_out0[1:0];
assign v$SEL4_17971_out0 = v$A_11857_out0[7:4];
assign v$SEL4_17972_out0 = v$A_11861_out0[7:4];
assign v$SEL4_17975_out0 = v$A_11873_out0[7:4];
assign v$SEL4_17976_out0 = v$A_11877_out0[7:4];
assign v$B3_18469_out0 = v$SEL7_4333_out0;
assign v$B3_18481_out0 = v$SEL7_4345_out0;
assign v$G28_19161_out0 = v$MEMHALT_18405_out0 || v$PIPELINEHALT_15423_out0;
assign v$G28_19162_out0 = v$MEMHALT_18406_out0 || v$PIPELINEHALT_15424_out0;
assign v$_1630_out0 = { v$C1_8288_out0,v$_5014_out0 };
assign v$_1634_out0 = { v$C1_8292_out0,v$_5018_out0 };
assign v$G37_1672_out0 = !((v$B4_17534_out0 && !v$A4_15625_out0) || (!v$B4_17534_out0) && v$A4_15625_out0);
assign v$G37_1674_out0 = !((v$B4_17536_out0 && !v$A4_15627_out0) || (!v$B4_17536_out0) && v$A4_15627_out0);
assign v$A0_1885_out0 = v$SEL5_13345_out0;
assign v$A0_1888_out0 = v$SEL5_13348_out0;
assign v$A0_1897_out0 = v$SEL5_13357_out0;
assign v$A0_1900_out0 = v$SEL5_13360_out0;
assign v$RAMAddress_2469_out0 = v$RAMADDRESS_13291_out0;
assign v$RAMAddress_2470_out0 = v$RAMADDRESS_13292_out0;
assign v$SEL4_2485_out0 = v$B$MANTISA_5124_out0[22:0];
assign v$SEL4_2486_out0 = v$B$MANTISA_5125_out0[22:0];
assign v$EQ1_3162_out0 = v$ADDRESS_6098_out0 == 12'hff8;
assign v$EQ1_3163_out0 = v$ADDRESS_6099_out0 == 12'hff8;
assign v$G21_3731_out0 = ! v$B1_14831_out0;
assign v$G21_3743_out0 = ! v$B1_14843_out0;
assign v$EQ5_3752_out0 = v$ADDRESS_6098_out0 == 12'hff7;
assign v$EQ5_3753_out0 = v$ADDRESS_6099_out0 == 12'hff7;
assign v$B0_3842_out0 = v$SEL10_13195_out0;
assign v$B0_3846_out0 = v$SEL10_13199_out0;
assign v$B0_3847_out0 = v$SEL10_13200_out0;
assign v$B0_3854_out0 = v$SEL10_13207_out0;
assign v$B0_3858_out0 = v$SEL10_13211_out0;
assign v$B0_3859_out0 = v$SEL10_13212_out0;
assign v$G8_3916_out0 = !((v$A3_11209_out0 && !v$B3_18469_out0) || (!v$A3_11209_out0) && v$B3_18469_out0);
assign v$G8_3928_out0 = !((v$A3_11221_out0 && !v$B3_18481_out0) || (!v$A3_11221_out0) && v$B3_18481_out0);
assign v$MUX3_3953_out0 = v$IS$SUB_13643_out0 ? v$C8_14199_out0 : v$C1_16843_out0;
assign v$MUX3_3954_out0 = v$IS$SUB_13644_out0 ? v$C8_14200_out0 : v$C1_16844_out0;
assign v$G36_6193_out0 = !((v$B3_18469_out0 && !v$A3_11209_out0) || (!v$B3_18469_out0) && v$A3_11209_out0);
assign v$G36_6205_out0 = !((v$B3_18481_out0 && !v$A3_11221_out0) || (!v$B3_18481_out0) && v$A3_11221_out0);
assign v$EXTHALT_6705_out0 = v$G28_19161_out0;
assign v$EXTHALT_6706_out0 = v$G28_19162_out0;
assign v$G6_6792_out0 = ! v$B3_18469_out0;
assign v$G6_6804_out0 = ! v$B3_18481_out0;
assign v$G3_7805_out0 = !((v$A4_15625_out0 && !v$B4_17534_out0) || (!v$A4_15625_out0) && v$B4_17534_out0);
assign v$G3_7807_out0 = !((v$A4_15627_out0 && !v$B4_17536_out0) || (!v$A4_15627_out0) && v$B4_17536_out0);
assign v$MUX5_8281_out0 = v$S_10894_out0 ? v$_14777_out0 : v$C1_3229_out0;
assign v$MUX5_8282_out0 = v$S_10895_out0 ? v$_14778_out0 : v$C1_3230_out0;
assign v$A2_8371_out0 = v$SEL3_8730_out0;
assign v$A2_8374_out0 = v$SEL3_8733_out0;
assign v$A2_8383_out0 = v$SEL3_8742_out0;
assign v$A2_8386_out0 = v$SEL3_8745_out0;
assign v$G17_8496_out0 = !((v$A0_1894_out0 && !v$B0_3845_out0) || (!v$A0_1894_out0) && v$B0_3845_out0);
assign v$G17_8508_out0 = !((v$A0_1906_out0 && !v$B0_3857_out0) || (!v$A0_1906_out0) && v$B0_3857_out0);
assign v$V0_9720_out0 = v$VALID0_13990_out0;
assign v$_9820_out0 = { v$_17369_out0,v$S$REG_3653_out0 };
assign v$_9824_out0 = { v$_17373_out0,v$S$REG_3654_out0 };
assign v$A3_11200_out0 = v$SEL2_17220_out0;
assign v$A3_11203_out0 = v$SEL2_17223_out0;
assign v$A3_11212_out0 = v$SEL2_17232_out0;
assign v$A3_11215_out0 = v$SEL2_17235_out0;
assign v$SEL2_11519_out0 = v$B$MANTISA_5124_out0[22:0];
assign v$SEL2_11520_out0 = v$B$MANTISA_5125_out0[22:0];
assign v$A_11858_out0 = v$SEL4_17971_out0;
assign v$A_11859_out0 = v$SEL1_10745_out0;
assign v$A_11862_out0 = v$SEL4_17972_out0;
assign v$A_11863_out0 = v$SEL1_10746_out0;
assign v$A_11874_out0 = v$SEL4_17975_out0;
assign v$A_11875_out0 = v$SEL1_10749_out0;
assign v$A_11878_out0 = v$SEL4_17976_out0;
assign v$A_11879_out0 = v$SEL1_10750_out0;
assign v$EQ3_12280_out0 = v$ADDRESS_6098_out0 == 12'hffa;
assign v$EQ3_12281_out0 = v$ADDRESS_6099_out0 == 12'hffa;
assign v$G23_12749_out0 = ! v$B0_3845_out0;
assign v$G23_12761_out0 = ! v$B0_3857_out0;
assign v$RAMADDR1_13239_out0 = v$RAM$ADDR1_6700_out0;
assign v$G33_13684_out0 = !((v$A0_1894_out0 && !v$B0_3845_out0) || (!v$A0_1894_out0) && v$B0_3845_out0);
assign v$G33_13696_out0 = !((v$A0_1906_out0 && !v$B0_3857_out0) || (!v$A0_1906_out0) && v$B0_3857_out0);
assign v$G1_13768_out0 = ! v$B4_17534_out0;
assign v$G1_13770_out0 = ! v$B4_17536_out0;
assign v$_13803_out0 = { v$_12334_out0,v$_12334_out0 };
assign v$_13804_out0 = { v$_12335_out0,v$_12335_out0 };
assign v$_13891_out0 = { v$_15202_out0,v$_17652_out0 };
assign v$_13895_out0 = { v$_15206_out0,v$_17653_out0 };
assign v$G15_14231_out0 = !((v$A2_8380_out0 && !v$B2_17253_out0) || (!v$A2_8380_out0) && v$B2_17253_out0);
assign v$G15_14243_out0 = !((v$A2_8392_out0 && !v$B2_17265_out0) || (!v$A2_8392_out0) && v$B2_17265_out0);
assign v$B1_14828_out0 = v$SEL9_11342_out0;
assign v$B1_14832_out0 = v$SEL9_11346_out0;
assign v$B1_14833_out0 = v$SEL9_11347_out0;
assign v$B1_14840_out0 = v$SEL9_11354_out0;
assign v$B1_14844_out0 = v$SEL9_11358_out0;
assign v$B1_14845_out0 = v$SEL9_11359_out0;
assign v$A1_14943_out0 = v$SEL4_7652_out0;
assign v$A1_14946_out0 = v$SEL4_7655_out0;
assign v$A1_14955_out0 = v$SEL4_7664_out0;
assign v$A1_14958_out0 = v$SEL4_7667_out0;
assign v$B_15037_out0 = v$B$EXP_17295_out0;
assign v$B_15053_out0 = v$B$EXP_17299_out0;
assign v$G35_15131_out0 = !((v$A2_8380_out0 && !v$B2_17253_out0) || (!v$A2_8380_out0) && v$B2_17253_out0);
assign v$G35_15143_out0 = !((v$A2_8392_out0 && !v$B2_17265_out0) || (!v$A2_8392_out0) && v$B2_17265_out0);
assign v$CIN_15670_out0 = v$IS$SUB_13643_out0;
assign v$CIN_15673_out0 = v$IS$SUB_13644_out0;
assign v$EQ12_15715_out0 = v$ADDRESS_6098_out0 == 12'hff6;
assign v$EQ12_15716_out0 = v$ADDRESS_6099_out0 == 12'hff6;
assign v$S_16064_out0 = v$HALT_13471_out0;
assign v$S_16067_out0 = v$HALT_13472_out0;
assign v$B$MANTISA_16181_out0 = v$MUX5_1767_out0;
assign v$B$MANTISA_16182_out0 = v$MUX5_1768_out0;
assign v$G12_17103_out0 = ! v$B2_17253_out0;
assign v$G12_17115_out0 = ! v$B2_17265_out0;
assign v$EQ4_17198_out0 = v$ADDRESS_6098_out0 == 12'hffb;
assign v$EQ4_17199_out0 = v$ADDRESS_6099_out0 == 12'hffb;
assign v$B2_17250_out0 = v$SEL8_13490_out0;
assign v$B2_17254_out0 = v$SEL8_13494_out0;
assign v$B2_17255_out0 = v$SEL8_13495_out0;
assign v$B2_17262_out0 = v$SEL8_13502_out0;
assign v$B2_17266_out0 = v$SEL8_13506_out0;
assign v$B2_17267_out0 = v$SEL8_13507_out0;
assign v$G16_17482_out0 = !((v$A1_14952_out0 && !v$B1_14831_out0) || (!v$A1_14952_out0) && v$B1_14831_out0);
assign v$G16_17494_out0 = !((v$A1_14964_out0 && !v$B1_14843_out0) || (!v$A1_14964_out0) && v$B1_14843_out0);
assign v$EQ2_17513_out0 = v$ADDRESS_6098_out0 == 12'hff9;
assign v$EQ2_17514_out0 = v$ADDRESS_6099_out0 == 12'hff9;
assign v$B4_17533_out0 = v$SEL6_6092_out0;
assign v$B4_17535_out0 = v$SEL6_6094_out0;
assign v$RAMADDR0_17579_out0 = v$RAM$ADDR0_13120_out0;
assign v$G34_17940_out0 = !((v$A1_14952_out0 && !v$B1_14831_out0) || (!v$A1_14952_out0) && v$B1_14831_out0);
assign v$G34_17952_out0 = !((v$A1_14964_out0 && !v$B1_14843_out0) || (!v$A1_14964_out0) && v$B1_14843_out0);
assign v$V1_18443_out0 = v$VALID1_9151_out0;
assign v$B3_18466_out0 = v$SEL7_4330_out0;
assign v$B3_18470_out0 = v$SEL7_4334_out0;
assign v$B3_18471_out0 = v$SEL7_4335_out0;
assign v$B3_18478_out0 = v$SEL7_4342_out0;
assign v$B3_18482_out0 = v$SEL7_4346_out0;
assign v$B3_18483_out0 = v$SEL7_4347_out0;
assign v$G65_18812_out0 = v$HALT_13471_out0 || v$G64_6638_out0;
assign v$G65_18813_out0 = v$HALT_13472_out0 || v$G64_6639_out0;
assign v$G13_200_out0 = v$EQ12_15715_out0 && v$WEN_3862_out0;
assign v$G13_201_out0 = v$EQ12_15716_out0 && v$WEN_3863_out0;
assign v$MUX6_1472_out0 = v$FF1_16930_out0 ? v$S$REG_3653_out0 : v$_13803_out0;
assign v$MUX6_1473_out0 = v$FF1_16931_out0 ? v$S$REG_3654_out0 : v$_13804_out0;
assign v$A4XNORB4_1536_out0 = v$G3_7805_out0;
assign v$A4XNORB4_1538_out0 = v$G3_7807_out0;
assign v$A0XNORB0_1592_out0 = v$G17_8496_out0;
assign v$A0XNORB0_1604_out0 = v$G17_8508_out0;
assign v$G37_1671_out0 = !((v$B4_17533_out0 && !v$A4_15624_out0) || (!v$B4_17533_out0) && v$A4_15624_out0);
assign v$G37_1673_out0 = !((v$B4_17535_out0 && !v$A4_15626_out0) || (!v$B4_17535_out0) && v$A4_15626_out0);
assign v$B$MANTISSA_2870_out0 = v$B$MANTISA_16181_out0;
assign v$B$MANTISSA_2871_out0 = v$B$MANTISA_16182_out0;
assign v$ADD_3164_out0 = v$RAMAddress_2469_out0;
assign v$ADD_3165_out0 = v$RAMAddress_2470_out0;
assign v$G21_3728_out0 = ! v$B1_14828_out0;
assign v$G21_3732_out0 = ! v$B1_14832_out0;
assign v$G21_3733_out0 = ! v$B1_14833_out0;
assign v$G21_3740_out0 = ! v$B1_14840_out0;
assign v$G21_3744_out0 = ! v$B1_14844_out0;
assign v$G21_3745_out0 = ! v$B1_14845_out0;
assign v$G8_3913_out0 = !((v$A3_11206_out0 && !v$B3_18466_out0) || (!v$A3_11206_out0) && v$B3_18466_out0);
assign v$G8_3917_out0 = !((v$A3_11210_out0 && !v$B3_18470_out0) || (!v$A3_11210_out0) && v$B3_18470_out0);
assign v$G8_3918_out0 = !((v$A3_11211_out0 && !v$B3_18471_out0) || (!v$A3_11211_out0) && v$B3_18471_out0);
assign v$G8_3925_out0 = !((v$A3_11218_out0 && !v$B3_18478_out0) || (!v$A3_11218_out0) && v$B3_18478_out0);
assign v$G8_3929_out0 = !((v$A3_11222_out0 && !v$B3_18482_out0) || (!v$A3_11222_out0) && v$B3_18482_out0);
assign v$G8_3930_out0 = !((v$A3_11223_out0 && !v$B3_18483_out0) || (!v$A3_11223_out0) && v$B3_18483_out0);
assign v$A2XNORB2_4668_out0 = v$G15_14231_out0;
assign v$A2XNORB2_4680_out0 = v$G15_14243_out0;
assign v$G30_5138_out0 = !(v$EXTHALT_6705_out0 || v$STPHALT_4478_out0);
assign v$G30_5139_out0 = !(v$EXTHALT_6706_out0 || v$STPHALT_4479_out0);
assign v$G36_6190_out0 = !((v$B3_18466_out0 && !v$A3_11206_out0) || (!v$B3_18466_out0) && v$A3_11206_out0);
assign v$G36_6194_out0 = !((v$B3_18470_out0 && !v$A3_11210_out0) || (!v$B3_18470_out0) && v$A3_11210_out0);
assign v$G36_6195_out0 = !((v$B3_18471_out0 && !v$A3_11211_out0) || (!v$B3_18471_out0) && v$A3_11211_out0);
assign v$G36_6202_out0 = !((v$B3_18478_out0 && !v$A3_11218_out0) || (!v$B3_18478_out0) && v$A3_11218_out0);
assign v$G36_6206_out0 = !((v$B3_18482_out0 && !v$A3_11222_out0) || (!v$B3_18482_out0) && v$A3_11222_out0);
assign v$G36_6207_out0 = !((v$B3_18483_out0 && !v$A3_11223_out0) || (!v$B3_18483_out0) && v$A3_11223_out0);
assign v$G6_6789_out0 = ! v$B3_18466_out0;
assign v$G6_6793_out0 = ! v$B3_18470_out0;
assign v$G6_6794_out0 = ! v$B3_18471_out0;
assign v$G6_6801_out0 = ! v$B3_18478_out0;
assign v$G6_6805_out0 = ! v$B3_18482_out0;
assign v$G6_6806_out0 = ! v$B3_18483_out0;
assign v$MUX6_7182_out0 = v$G70_14638_out0 ? v$REG12_3553_out0 : v$RAMADDR1_13239_out0;
assign v$G5_7224_out0 = v$A3_11209_out0 && v$G6_6792_out0;
assign v$G5_7236_out0 = v$A3_11221_out0 && v$G6_6804_out0;
assign v$G38_7618_out0 = v$G33_13684_out0 && v$G34_17940_out0;
assign v$G38_7630_out0 = v$G33_13696_out0 && v$G34_17952_out0;
assign v$SEL4_7653_out0 = v$A_11858_out0[1:1];
assign v$SEL4_7654_out0 = v$A_11859_out0[1:1];
assign v$SEL4_7656_out0 = v$A_11862_out0[1:1];
assign v$SEL4_7657_out0 = v$A_11863_out0[1:1];
assign v$SEL4_7665_out0 = v$A_11874_out0[1:1];
assign v$SEL4_7666_out0 = v$A_11875_out0[1:1];
assign v$SEL4_7668_out0 = v$A_11878_out0[1:1];
assign v$SEL4_7669_out0 = v$A_11879_out0[1:1];
assign v$G3_7804_out0 = !((v$A4_15624_out0 && !v$B4_17533_out0) || (!v$A4_15624_out0) && v$B4_17533_out0);
assign v$G3_7806_out0 = !((v$A4_15626_out0 && !v$B4_17535_out0) || (!v$A4_15626_out0) && v$B4_17535_out0);
assign v$G3_7838_out0 = v$EQ2_17513_out0 && v$WEN_3862_out0;
assign v$G3_7839_out0 = v$EQ2_17514_out0 && v$WEN_3863_out0;
assign v$S_8337_out0 = v$S_16064_out0;
assign v$S_8340_out0 = v$S_16067_out0;
assign v$G17_8493_out0 = !((v$A0_1891_out0 && !v$B0_3842_out0) || (!v$A0_1891_out0) && v$B0_3842_out0);
assign v$G17_8497_out0 = !((v$A0_1895_out0 && !v$B0_3846_out0) || (!v$A0_1895_out0) && v$B0_3846_out0);
assign v$G17_8498_out0 = !((v$A0_1896_out0 && !v$B0_3847_out0) || (!v$A0_1896_out0) && v$B0_3847_out0);
assign v$G17_8505_out0 = !((v$A0_1903_out0 && !v$B0_3854_out0) || (!v$A0_1903_out0) && v$B0_3854_out0);
assign v$G17_8509_out0 = !((v$A0_1907_out0 && !v$B0_3858_out0) || (!v$A0_1907_out0) && v$B0_3858_out0);
assign v$G17_8510_out0 = !((v$A0_1908_out0 && !v$B0_3859_out0) || (!v$A0_1908_out0) && v$B0_3859_out0);
assign v$SEL3_8731_out0 = v$A_11858_out0[2:2];
assign v$SEL3_8732_out0 = v$A_11859_out0[2:2];
assign v$SEL3_8734_out0 = v$A_11862_out0[2:2];
assign v$SEL3_8735_out0 = v$A_11863_out0[2:2];
assign v$SEL3_8743_out0 = v$A_11874_out0[2:2];
assign v$SEL3_8744_out0 = v$A_11875_out0[2:2];
assign v$SEL3_8746_out0 = v$A_11878_out0[2:2];
assign v$SEL3_8747_out0 = v$A_11879_out0[2:2];
assign v$G66_9020_out0 = ! v$G65_18812_out0;
assign v$G66_9021_out0 = ! v$G65_18813_out0;
assign v$SEL3_9375_out0 = v$B_15037_out0[7:4];
assign v$SEL3_9379_out0 = v$B_15053_out0[7:4];
assign v$MUX3_9451_out0 = v$G66_9263_out0 ? v$REG9_16701_out0 : v$RAMADDR0_17579_out0;
assign v$G20_10312_out0 = v$A1_14952_out0 && v$G21_3731_out0;
assign v$G20_10324_out0 = v$A1_14964_out0 && v$G21_3743_out0;
assign v$G2_10852_out0 = v$A4_15625_out0 && v$G1_13768_out0;
assign v$G2_10854_out0 = v$A4_15627_out0 && v$G1_13770_out0;
assign v$G25_11448_out0 = v$A0_1894_out0 && v$G23_12749_out0;
assign v$G25_11460_out0 = v$A0_1906_out0 && v$G23_12761_out0;
assign v$G23_12746_out0 = ! v$B0_3842_out0;
assign v$G23_12750_out0 = ! v$B0_3846_out0;
assign v$G23_12751_out0 = ! v$B0_3847_out0;
assign v$G23_12758_out0 = ! v$B0_3854_out0;
assign v$G23_12762_out0 = ! v$B0_3858_out0;
assign v$G23_12763_out0 = ! v$B0_3859_out0;
assign v$G5_13317_out0 = v$EQ5_3752_out0 && v$WEN_3862_out0;
assign v$G5_13318_out0 = v$EQ5_3753_out0 && v$WEN_3863_out0;
assign v$SEL5_13346_out0 = v$A_11858_out0[0:0];
assign v$SEL5_13347_out0 = v$A_11859_out0[0:0];
assign v$SEL5_13349_out0 = v$A_11862_out0[0:0];
assign v$SEL5_13350_out0 = v$A_11863_out0[0:0];
assign v$SEL5_13358_out0 = v$A_11874_out0[0:0];
assign v$SEL5_13359_out0 = v$A_11875_out0[0:0];
assign v$SEL5_13361_out0 = v$A_11878_out0[0:0];
assign v$SEL5_13362_out0 = v$A_11879_out0[0:0];
assign v$G33_13681_out0 = !((v$A0_1891_out0 && !v$B0_3842_out0) || (!v$A0_1891_out0) && v$B0_3842_out0);
assign v$G33_13685_out0 = !((v$A0_1895_out0 && !v$B0_3846_out0) || (!v$A0_1895_out0) && v$B0_3846_out0);
assign v$G33_13686_out0 = !((v$A0_1896_out0 && !v$B0_3847_out0) || (!v$A0_1896_out0) && v$B0_3847_out0);
assign v$G33_13693_out0 = !((v$A0_1903_out0 && !v$B0_3854_out0) || (!v$A0_1903_out0) && v$B0_3854_out0);
assign v$G33_13697_out0 = !((v$A0_1907_out0 && !v$B0_3858_out0) || (!v$A0_1907_out0) && v$B0_3858_out0);
assign v$G33_13698_out0 = !((v$A0_1908_out0 && !v$B0_3859_out0) || (!v$A0_1908_out0) && v$B0_3859_out0);
assign v$G1_13767_out0 = ! v$B4_17533_out0;
assign v$G1_13769_out0 = ! v$B4_17535_out0;
assign v$G15_14228_out0 = !((v$A2_8377_out0 && !v$B2_17250_out0) || (!v$A2_8377_out0) && v$B2_17250_out0);
assign v$G15_14232_out0 = !((v$A2_8381_out0 && !v$B2_17254_out0) || (!v$A2_8381_out0) && v$B2_17254_out0);
assign v$G15_14233_out0 = !((v$A2_8382_out0 && !v$B2_17255_out0) || (!v$A2_8382_out0) && v$B2_17255_out0);
assign v$G15_14240_out0 = !((v$A2_8389_out0 && !v$B2_17262_out0) || (!v$A2_8389_out0) && v$B2_17262_out0);
assign v$G15_14244_out0 = !((v$A2_8393_out0 && !v$B2_17266_out0) || (!v$A2_8393_out0) && v$B2_17266_out0);
assign v$G15_14245_out0 = !((v$A2_8394_out0 && !v$B2_17267_out0) || (!v$A2_8394_out0) && v$B2_17267_out0);
assign v$G2_14274_out0 = v$EQ3_12280_out0 && v$WEN_3862_out0;
assign v$G2_14275_out0 = v$EQ3_12281_out0 && v$WEN_3863_out0;
assign v$VALID_15094_out0 = v$V1_18443_out0;
assign v$VALID_15095_out0 = v$V0_9720_out0;
assign v$G35_15128_out0 = !((v$A2_8377_out0 && !v$B2_17250_out0) || (!v$A2_8377_out0) && v$B2_17250_out0);
assign v$G35_15132_out0 = !((v$A2_8381_out0 && !v$B2_17254_out0) || (!v$A2_8381_out0) && v$B2_17254_out0);
assign v$G35_15133_out0 = !((v$A2_8382_out0 && !v$B2_17255_out0) || (!v$A2_8382_out0) && v$B2_17255_out0);
assign v$G35_15140_out0 = !((v$A2_8389_out0 && !v$B2_17262_out0) || (!v$A2_8389_out0) && v$B2_17262_out0);
assign v$G35_15144_out0 = !((v$A2_8393_out0 && !v$B2_17266_out0) || (!v$A2_8393_out0) && v$B2_17266_out0);
assign v$G35_15145_out0 = !((v$A2_8394_out0 && !v$B2_17267_out0) || (!v$A2_8394_out0) && v$B2_17267_out0);
assign v$A3XNORB3_15332_out0 = v$G8_3916_out0;
assign v$A3XNORB3_15344_out0 = v$G8_3928_out0;
assign v$G4_15735_out0 = v$EQ1_3162_out0 && v$WEN_3862_out0;
assign v$G4_15736_out0 = v$EQ1_3163_out0 && v$WEN_3863_out0;
assign v$G11_16239_out0 = v$A2_8380_out0 && v$G12_17103_out0;
assign v$G11_16251_out0 = v$A2_8392_out0 && v$G12_17115_out0;
assign v$MUX4_16601_out0 = v$EN_17562_out0 ? v$_1630_out0 : v$IN_9947_out0;
assign v$MUX4_16605_out0 = v$EN_17566_out0 ? v$_1634_out0 : v$IN_9951_out0;
assign v$A1XNORB1_16668_out0 = v$G16_17482_out0;
assign v$A1XNORB1_16680_out0 = v$G16_17494_out0;
assign v$G12_17100_out0 = ! v$B2_17250_out0;
assign v$G12_17104_out0 = ! v$B2_17254_out0;
assign v$G12_17105_out0 = ! v$B2_17255_out0;
assign v$G12_17112_out0 = ! v$B2_17262_out0;
assign v$G12_17116_out0 = ! v$B2_17266_out0;
assign v$G12_17117_out0 = ! v$B2_17267_out0;
assign v$G1_17122_out0 = v$EQ4_17198_out0 && v$WEN_3862_out0;
assign v$G1_17123_out0 = v$EQ4_17199_out0 && v$WEN_3863_out0;
assign v$SEL2_17221_out0 = v$A_11858_out0[3:3];
assign v$SEL2_17222_out0 = v$A_11859_out0[3:3];
assign v$SEL2_17224_out0 = v$A_11862_out0[3:3];
assign v$SEL2_17225_out0 = v$A_11863_out0[3:3];
assign v$SEL2_17233_out0 = v$A_11874_out0[3:3];
assign v$SEL2_17234_out0 = v$A_11875_out0[3:3];
assign v$SEL2_17236_out0 = v$A_11878_out0[3:3];
assign v$SEL2_17237_out0 = v$A_11879_out0[3:3];
assign v$G16_17479_out0 = !((v$A1_14949_out0 && !v$B1_14828_out0) || (!v$A1_14949_out0) && v$B1_14828_out0);
assign v$G16_17483_out0 = !((v$A1_14953_out0 && !v$B1_14832_out0) || (!v$A1_14953_out0) && v$B1_14832_out0);
assign v$G16_17484_out0 = !((v$A1_14954_out0 && !v$B1_14833_out0) || (!v$A1_14954_out0) && v$B1_14833_out0);
assign v$G16_17491_out0 = !((v$A1_14961_out0 && !v$B1_14840_out0) || (!v$A1_14961_out0) && v$B1_14840_out0);
assign v$G16_17495_out0 = !((v$A1_14965_out0 && !v$B1_14844_out0) || (!v$A1_14965_out0) && v$B1_14844_out0);
assign v$G16_17496_out0 = !((v$A1_14966_out0 && !v$B1_14845_out0) || (!v$A1_14966_out0) && v$B1_14845_out0);
assign v$G34_17937_out0 = !((v$A1_14949_out0 && !v$B1_14828_out0) || (!v$A1_14949_out0) && v$B1_14828_out0);
assign v$G34_17941_out0 = !((v$A1_14953_out0 && !v$B1_14832_out0) || (!v$A1_14953_out0) && v$B1_14832_out0);
assign v$G34_17942_out0 = !((v$A1_14954_out0 && !v$B1_14833_out0) || (!v$A1_14954_out0) && v$B1_14833_out0);
assign v$G34_17949_out0 = !((v$A1_14961_out0 && !v$B1_14840_out0) || (!v$A1_14961_out0) && v$B1_14840_out0);
assign v$G34_17953_out0 = !((v$A1_14965_out0 && !v$B1_14844_out0) || (!v$A1_14965_out0) && v$B1_14844_out0);
assign v$G34_17954_out0 = !((v$A1_14966_out0 && !v$B1_14845_out0) || (!v$A1_14966_out0) && v$B1_14845_out0);
assign v$CIN_17984_out0 = v$CIN_15670_out0;
assign v$CIN_17987_out0 = v$CIN_15673_out0;
assign v$G39_18002_out0 = v$G36_6193_out0 && v$G37_1672_out0;
assign v$G39_18004_out0 = v$G36_6205_out0 && v$G37_1674_out0;
assign v$SEL2_18084_out0 = v$B_15037_out0[3:0];
assign v$SEL2_18088_out0 = v$B_15053_out0[3:0];
assign v$I3REGISTERWRITE_1419_out0 = v$G1_17122_out0;
assign v$I3REGISTERWRITE_1420_out0 = v$G1_17123_out0;
assign v$SEL4_1527_out0 = v$B$MANTISSA_2870_out0[23:12];
assign v$SEL4_1528_out0 = v$B$MANTISSA_2871_out0[23:12];
assign v$A4XNORB4_1535_out0 = v$G3_7804_out0;
assign v$A4XNORB4_1537_out0 = v$G3_7806_out0;
assign v$A0XNORB0_1589_out0 = v$G17_8493_out0;
assign v$A0XNORB0_1593_out0 = v$G17_8497_out0;
assign v$A0XNORB0_1594_out0 = v$G17_8498_out0;
assign v$A0XNORB0_1601_out0 = v$G17_8505_out0;
assign v$A0XNORB0_1605_out0 = v$G17_8509_out0;
assign v$A0XNORB0_1606_out0 = v$G17_8510_out0;
assign v$COUNTEREN_1782_out0 = v$G13_200_out0;
assign v$COUNTEREN_1783_out0 = v$G13_201_out0;
assign v$A0_1886_out0 = v$SEL5_13346_out0;
assign v$A0_1887_out0 = v$SEL5_13347_out0;
assign v$A0_1889_out0 = v$SEL5_13349_out0;
assign v$A0_1890_out0 = v$SEL5_13350_out0;
assign v$A0_1898_out0 = v$SEL5_13358_out0;
assign v$A0_1899_out0 = v$SEL5_13359_out0;
assign v$A0_1901_out0 = v$SEL5_13361_out0;
assign v$A0_1902_out0 = v$SEL5_13362_out0;
assign v$MUX1_2011_out0 = v$SELIN_18816_out0 ? v$MUX6_7182_out0 : v$MUX3_9451_out0;
assign v$G7_2443_out0 = v$A4XNORB4_1536_out0 && v$G5_7224_out0;
assign v$G7_2445_out0 = v$A4XNORB4_1538_out0 && v$G5_7236_out0;
assign v$I1REGISTERWRITE_3139_out0 = v$G3_7838_out0;
assign v$I1REGISTERWRITE_3140_out0 = v$G3_7839_out0;
assign v$I0REGISTERWRITE_3578_out0 = v$G4_15735_out0;
assign v$I0REGISTERWRITE_3579_out0 = v$G4_15736_out0;
assign v$ModeRegAdd_4164_out0 = v$ADD_3164_out0 == 12'hffc;
assign v$ModeRegAdd_4165_out0 = v$ADD_3165_out0 == 12'hffc;
assign v$G13_4573_out0 = v$A3XNORB3_15332_out0 && v$G11_16239_out0;
assign v$G13_4585_out0 = v$A3XNORB3_15344_out0 && v$G11_16251_out0;
assign v$A2XNORB2_4665_out0 = v$G15_14228_out0;
assign v$A2XNORB2_4669_out0 = v$G15_14232_out0;
assign v$A2XNORB2_4670_out0 = v$G15_14233_out0;
assign v$A2XNORB2_4677_out0 = v$G15_14240_out0;
assign v$A2XNORB2_4681_out0 = v$G15_14244_out0;
assign v$A2XNORB2_4682_out0 = v$G15_14245_out0;
assign v$MODEEN_6041_out0 = v$G5_13317_out0;
assign v$MODEEN_6042_out0 = v$G5_13318_out0;
assign v$G5_7221_out0 = v$A3_11206_out0 && v$G6_6789_out0;
assign v$G5_7225_out0 = v$A3_11210_out0 && v$G6_6793_out0;
assign v$G5_7226_out0 = v$A3_11211_out0 && v$G6_6794_out0;
assign v$G5_7233_out0 = v$A3_11218_out0 && v$G6_6801_out0;
assign v$G5_7237_out0 = v$A3_11222_out0 && v$G6_6805_out0;
assign v$G5_7238_out0 = v$A3_11223_out0 && v$G6_6806_out0;
assign v$G38_7615_out0 = v$G33_13681_out0 && v$G34_17937_out0;
assign v$G38_7619_out0 = v$G33_13685_out0 && v$G34_17941_out0;
assign v$G38_7620_out0 = v$G33_13686_out0 && v$G34_17942_out0;
assign v$G38_7627_out0 = v$G33_13693_out0 && v$G34_17949_out0;
assign v$G38_7631_out0 = v$G33_13697_out0 && v$G34_17953_out0;
assign v$G38_7632_out0 = v$G33_13698_out0 && v$G34_17954_out0;
assign v$A4$COMP$B4_7726_out0 = v$G2_10852_out0;
assign v$A4$COMP$B4_7728_out0 = v$G2_10854_out0;
assign v$StatRegAdd_8059_out0 = v$ADD_3164_out0 == 12'hffd;
assign v$StatRegAdd_8060_out0 = v$ADD_3165_out0 == 12'hffd;
assign v$A2_8372_out0 = v$SEL3_8731_out0;
assign v$A2_8373_out0 = v$SEL3_8732_out0;
assign v$A2_8375_out0 = v$SEL3_8734_out0;
assign v$A2_8376_out0 = v$SEL3_8735_out0;
assign v$A2_8384_out0 = v$SEL3_8743_out0;
assign v$A2_8385_out0 = v$SEL3_8744_out0;
assign v$A2_8387_out0 = v$SEL3_8746_out0;
assign v$A2_8388_out0 = v$SEL3_8747_out0;
assign v$EN_9408_out0 = v$G30_5138_out0;
assign v$EN_9409_out0 = v$G30_5139_out0;
assign v$G20_10309_out0 = v$A1_14949_out0 && v$G21_3728_out0;
assign v$G20_10313_out0 = v$A1_14953_out0 && v$G21_3732_out0;
assign v$G20_10314_out0 = v$A1_14954_out0 && v$G21_3733_out0;
assign v$G20_10321_out0 = v$A1_14961_out0 && v$G21_3740_out0;
assign v$G20_10325_out0 = v$A1_14965_out0 && v$G21_3744_out0;
assign v$G20_10326_out0 = v$A1_14966_out0 && v$G21_3745_out0;
assign v$G2_10851_out0 = v$A4_15624_out0 && v$G1_13767_out0;
assign v$G2_10853_out0 = v$A4_15626_out0 && v$G1_13769_out0;
assign v$A3_11201_out0 = v$SEL2_17221_out0;
assign v$A3_11202_out0 = v$SEL2_17222_out0;
assign v$A3_11204_out0 = v$SEL2_17224_out0;
assign v$A3_11205_out0 = v$SEL2_17225_out0;
assign v$A3_11213_out0 = v$SEL2_17233_out0;
assign v$A3_11214_out0 = v$SEL2_17234_out0;
assign v$A3_11216_out0 = v$SEL2_17236_out0;
assign v$A3_11217_out0 = v$SEL2_17237_out0;
assign v$G25_11445_out0 = v$A0_1891_out0 && v$G23_12746_out0;
assign v$G25_11449_out0 = v$A0_1895_out0 && v$G23_12750_out0;
assign v$G25_11450_out0 = v$A0_1896_out0 && v$G23_12751_out0;
assign v$G25_11457_out0 = v$A0_1903_out0 && v$G23_12758_out0;
assign v$G25_11461_out0 = v$A0_1907_out0 && v$G23_12762_out0;
assign v$G25_11462_out0 = v$A0_1908_out0 && v$G23_12763_out0;
assign v$_12381_out0 = { v$_15238_out0,v$MUX6_1472_out0 };
assign v$_12385_out0 = { v$_15242_out0,v$MUX6_1473_out0 };
assign v$I2REGISTERWRITE_12504_out0 = v$G2_14274_out0;
assign v$I2REGISTERWRITE_12505_out0 = v$G2_14275_out0;
assign v$MUX2_12604_out0 = v$G3_2801_out0 ? v$_9820_out0 : v$MUX4_16601_out0;
assign v$MUX2_12608_out0 = v$G3_2805_out0 ? v$_9824_out0 : v$MUX4_16605_out0;
assign v$RXRegAdd_13546_out0 = v$ADD_3164_out0 == 12'hffe;
assign v$RXRegAdd_13547_out0 = v$ADD_3165_out0 == 12'hffe;
assign v$G28_13600_out0 = v$A1XNORB1_16668_out0 && v$G25_11448_out0;
assign v$G28_13612_out0 = v$A1XNORB1_16680_out0 && v$G25_11460_out0;
assign v$G22_13921_out0 = v$A2XNORB2_4668_out0 && v$G20_10312_out0;
assign v$G22_13933_out0 = v$A2XNORB2_4680_out0 && v$G20_10324_out0;
assign v$G40_13954_out0 = v$G35_15131_out0 && v$G39_18002_out0;
assign v$G40_13955_out0 = v$G35_15132_out0 && v$G36_6194_out0;
assign v$G40_13956_out0 = v$G35_15133_out0 && v$G36_6195_out0;
assign v$G40_13966_out0 = v$G35_15143_out0 && v$G39_18004_out0;
assign v$G40_13967_out0 = v$G35_15144_out0 && v$G36_6206_out0;
assign v$G40_13968_out0 = v$G35_15145_out0 && v$G36_6207_out0;
assign v$SEL2_14330_out0 = v$B$MANTISSA_2870_out0[11:0];
assign v$SEL2_14331_out0 = v$B$MANTISSA_2871_out0[11:0];
assign v$A1_14944_out0 = v$SEL4_7653_out0;
assign v$A1_14945_out0 = v$SEL4_7654_out0;
assign v$A1_14947_out0 = v$SEL4_7656_out0;
assign v$A1_14948_out0 = v$SEL4_7657_out0;
assign v$A1_14956_out0 = v$SEL4_7665_out0;
assign v$A1_14957_out0 = v$SEL4_7666_out0;
assign v$A1_14959_out0 = v$SEL4_7668_out0;
assign v$A1_14960_out0 = v$SEL4_7669_out0;
assign v$B_15038_out0 = v$SEL3_9375_out0;
assign v$B_15039_out0 = v$SEL2_18084_out0;
assign v$B_15054_out0 = v$SEL3_9379_out0;
assign v$B_15055_out0 = v$SEL2_18088_out0;
assign v$StatRegAdd1_15154_out0 = v$ADD_3164_out0 == 12'hffd;
assign v$StatRegAdd1_15155_out0 = v$ADD_3165_out0 == 12'hffd;
assign v$A3XNORB3_15329_out0 = v$G8_3913_out0;
assign v$A3XNORB3_15333_out0 = v$G8_3917_out0;
assign v$A3XNORB3_15334_out0 = v$G8_3918_out0;
assign v$A3XNORB3_15341_out0 = v$G8_3925_out0;
assign v$A3XNORB3_15345_out0 = v$G8_3929_out0;
assign v$A3XNORB3_15346_out0 = v$G8_3930_out0;
assign v$TXRegAdd_16193_out0 = v$ADD_3164_out0 == 12'hfff;
assign v$TXRegAdd_16194_out0 = v$ADD_3165_out0 == 12'hfff;
assign v$G11_16236_out0 = v$A2_8377_out0 && v$G12_17100_out0;
assign v$G11_16240_out0 = v$A2_8381_out0 && v$G12_17104_out0;
assign v$G11_16241_out0 = v$A2_8382_out0 && v$G12_17105_out0;
assign v$G11_16248_out0 = v$A2_8389_out0 && v$G12_17112_out0;
assign v$G11_16252_out0 = v$A2_8393_out0 && v$G12_17116_out0;
assign v$G11_16253_out0 = v$A2_8394_out0 && v$G12_17117_out0;
assign v$A1XNORB1_16665_out0 = v$G16_17479_out0;
assign v$A1XNORB1_16669_out0 = v$G16_17483_out0;
assign v$A1XNORB1_16670_out0 = v$G16_17484_out0;
assign v$A1XNORB1_16677_out0 = v$G16_17491_out0;
assign v$A1XNORB1_16681_out0 = v$G16_17495_out0;
assign v$A1XNORB1_16682_out0 = v$G16_17496_out0;
assign v$CIN_16718_out0 = v$CIN_17984_out0;
assign v$CIN_16721_out0 = v$CIN_17987_out0;
assign v$G39_18001_out0 = v$G36_6190_out0 && v$G37_1671_out0;
assign v$G39_18003_out0 = v$G36_6202_out0 && v$G37_1673_out0;
assign v$VALID_19282_out0 = v$VALID_15094_out0;
assign v$VALID_19283_out0 = v$VALID_15095_out0;
assign v$G7_2442_out0 = v$A4XNORB4_1535_out0 && v$G5_7221_out0;
assign v$G7_2444_out0 = v$A4XNORB4_1537_out0 && v$G5_7233_out0;
assign v$SEL7_4331_out0 = v$B_15038_out0[3:3];
assign v$SEL7_4332_out0 = v$B_15039_out0[3:3];
assign v$SEL7_4343_out0 = v$B_15054_out0[3:3];
assign v$SEL7_4344_out0 = v$B_15055_out0[3:3];
assign v$G13_4570_out0 = v$A3XNORB3_15329_out0 && v$G11_16236_out0;
assign v$G13_4574_out0 = v$A3XNORB3_15333_out0 && v$G11_16240_out0;
assign v$G13_4575_out0 = v$A3XNORB3_15334_out0 && v$G11_16241_out0;
assign v$G13_4582_out0 = v$A3XNORB3_15341_out0 && v$G11_16248_out0;
assign v$G13_4586_out0 = v$A3XNORB3_15345_out0 && v$G11_16252_out0;
assign v$G13_4587_out0 = v$A3XNORB3_15346_out0 && v$G11_16253_out0;
assign v$G27_4998_out0 = v$A2XNORB2_4668_out0 && v$G28_13600_out0;
assign v$G27_5010_out0 = v$A2XNORB2_4680_out0 && v$G28_13612_out0;
assign v$A3$COMP$B3_5169_out0 = v$G7_2443_out0;
assign v$A3$COMP$B3_5170_out0 = v$G5_7225_out0;
assign v$A3$COMP$B3_5171_out0 = v$G5_7226_out0;
assign v$A3$COMP$B3_5181_out0 = v$G7_2445_out0;
assign v$A3$COMP$B3_5182_out0 = v$G5_7237_out0;
assign v$A3$COMP$B3_5183_out0 = v$G5_7238_out0;
assign v$G18_5197_out0 = v$A3XNORB3_15332_out0 && v$G22_13921_out0;
assign v$G18_5209_out0 = v$A3XNORB3_15344_out0 && v$G22_13933_out0;
assign v$MUX1_6915_out0 = v$G4_4187_out0 ? v$_12381_out0 : v$MUX2_12604_out0;
assign v$MUX1_6919_out0 = v$G4_4191_out0 ? v$_12385_out0 : v$MUX2_12608_out0;
assign v$A4$COMP$B4_7725_out0 = v$G2_10851_out0;
assign v$A4$COMP$B4_7727_out0 = v$G2_10853_out0;
assign v$G3_7926_out0 = v$TXRegAdd_16193_out0 && v$WEN_18998_out0;
assign v$G3_7927_out0 = v$TXRegAdd_16194_out0 && v$WEN_18999_out0;
assign v$G7_8043_out0 = v$StatRegAdd1_15154_out0 && v$G8_13988_out0;
assign v$G7_8044_out0 = v$StatRegAdd1_15155_out0 && v$G8_13989_out0;
assign v$I0EN_8356_out0 = v$I0REGISTERWRITE_3578_out0;
assign v$I0EN_8357_out0 = v$I0REGISTERWRITE_3579_out0;
assign v$G5_8754_out0 = v$RXRegAdd_13546_out0 && v$G6_730_out0;
assign v$G5_8755_out0 = v$RXRegAdd_13547_out0 && v$G6_731_out0;
assign v$CINA_8815_out0 = v$CIN_16718_out0;
assign v$CINA_8938_out0 = v$CIN_16721_out0;
assign v$SEL9_11343_out0 = v$B_15038_out0[1:1];
assign v$SEL9_11344_out0 = v$B_15039_out0[1:1];
assign v$SEL9_11355_out0 = v$B_15054_out0[1:1];
assign v$SEL9_11356_out0 = v$B_15055_out0[1:1];
assign v$G41_11383_out0 = v$G38_7618_out0 && v$G40_13954_out0;
assign v$G41_11384_out0 = v$G38_7619_out0 && v$G40_13955_out0;
assign v$G41_11385_out0 = v$G38_7620_out0 && v$G40_13956_out0;
assign v$G41_11395_out0 = v$G38_7630_out0 && v$G40_13966_out0;
assign v$G41_11396_out0 = v$G38_7631_out0 && v$G40_13967_out0;
assign v$G41_11397_out0 = v$G38_7632_out0 && v$G40_13968_out0;
assign v$B_12696_out0 = v$SEL4_1527_out0;
assign v$B_12697_out0 = v$SEL2_14330_out0;
assign v$B_12698_out0 = v$SEL4_1528_out0;
assign v$B_12699_out0 = v$SEL2_14331_out0;
assign v$SEL10_13196_out0 = v$B_15038_out0[0:0];
assign v$SEL10_13197_out0 = v$B_15039_out0[0:0];
assign v$SEL10_13208_out0 = v$B_15054_out0[0:0];
assign v$SEL10_13209_out0 = v$B_15055_out0[0:0];
assign v$G14_13228_out0 = v$A4XNORB4_1536_out0 && v$G13_4573_out0;
assign v$G14_13230_out0 = v$A4XNORB4_1538_out0 && v$G13_4585_out0;
assign v$SEL8_13491_out0 = v$B_15038_out0[2:2];
assign v$SEL8_13492_out0 = v$B_15039_out0[2:2];
assign v$SEL8_13503_out0 = v$B_15054_out0[2:2];
assign v$SEL8_13504_out0 = v$B_15055_out0[2:2];
assign v$G28_13597_out0 = v$A1XNORB1_16665_out0 && v$G25_11445_out0;
assign v$G28_13601_out0 = v$A1XNORB1_16669_out0 && v$G25_11449_out0;
assign v$G28_13602_out0 = v$A1XNORB1_16670_out0 && v$G25_11450_out0;
assign v$G28_13609_out0 = v$A1XNORB1_16677_out0 && v$G25_11457_out0;
assign v$G28_13613_out0 = v$A1XNORB1_16681_out0 && v$G25_11461_out0;
assign v$G28_13614_out0 = v$A1XNORB1_16682_out0 && v$G25_11462_out0;
assign v$G22_13918_out0 = v$A2XNORB2_4665_out0 && v$G20_10309_out0;
assign v$G22_13922_out0 = v$A2XNORB2_4669_out0 && v$G20_10313_out0;
assign v$G22_13923_out0 = v$A2XNORB2_4670_out0 && v$G20_10314_out0;
assign v$G22_13930_out0 = v$A2XNORB2_4677_out0 && v$G20_10321_out0;
assign v$G22_13934_out0 = v$A2XNORB2_4681_out0 && v$G20_10325_out0;
assign v$G22_13935_out0 = v$A2XNORB2_4682_out0 && v$G20_10326_out0;
assign v$G40_13951_out0 = v$G35_15128_out0 && v$G39_18001_out0;
assign v$G40_13963_out0 = v$G35_15140_out0 && v$G39_18003_out0;
assign v$COUNTEREN_14035_out0 = v$COUNTEREN_1782_out0;
assign v$COUNTEREN_14036_out0 = v$COUNTEREN_1783_out0;
assign v$RAMADDR_14184_out0 = v$MUX1_2011_out0;
assign v$ENMODE_15175_out0 = v$MODEEN_6041_out0;
assign v$ENMODE_15176_out0 = v$MODEEN_6042_out0;
assign v$G9_16183_out0 = v$ModeRegAdd_4164_out0 && v$WEN_18998_out0;
assign v$G9_16184_out0 = v$ModeRegAdd_4165_out0 && v$WEN_18999_out0;
assign v$I2EN_16345_out0 = v$I2REGISTERWRITE_12504_out0;
assign v$I2EN_16346_out0 = v$I2REGISTERWRITE_12505_out0;
assign v$G1_17020_out0 = v$StatRegAdd_8059_out0 && v$WEN_18998_out0;
assign v$G1_17021_out0 = v$StatRegAdd_8060_out0 && v$WEN_18999_out0;
assign v$I3EN_18387_out0 = v$I3REGISTERWRITE_1419_out0;
assign v$I3EN_18388_out0 = v$I3REGISTERWRITE_1420_out0;
assign v$VALID_18531_out0 = v$VALID_19282_out0;
assign v$VALID_18532_out0 = v$VALID_19283_out0;
assign v$I1EN_19009_out0 = v$I1REGISTERWRITE_3139_out0;
assign v$I1EN_19010_out0 = v$I1REGISTERWRITE_3140_out0;
assign v$MUX3_2123_out0 = v$G8_2051_out0 ? v$_13891_out0 : v$MUX1_6915_out0;
assign v$MUX3_2127_out0 = v$G8_2055_out0 ? v$_13895_out0 : v$MUX1_6919_out0;
assign v$A2$COMP$B2_2144_out0 = v$G14_13228_out0;
assign v$A2$COMP$B2_2145_out0 = v$G13_4574_out0;
assign v$A2$COMP$B2_2146_out0 = v$G13_4575_out0;
assign v$A2$COMP$B2_2156_out0 = v$G14_13230_out0;
assign v$A2$COMP$B2_2157_out0 = v$G13_4586_out0;
assign v$A2$COMP$B2_2158_out0 = v$G13_4587_out0;
assign v$B0_3843_out0 = v$SEL10_13196_out0;
assign v$B0_3844_out0 = v$SEL10_13197_out0;
assign v$B0_3855_out0 = v$SEL10_13208_out0;
assign v$B0_3856_out0 = v$SEL10_13209_out0;
assign v$VALID_3893_out0 = v$VALID_18531_out0;
assign v$VALID_3894_out0 = v$VALID_18532_out0;
assign v$ModeWrite_4621_out0 = v$G9_16183_out0;
assign v$ModeWrite_4622_out0 = v$G9_16184_out0;
assign v$G27_4995_out0 = v$A2XNORB2_4665_out0 && v$G28_13597_out0;
assign v$G27_4999_out0 = v$A2XNORB2_4669_out0 && v$G28_13601_out0;
assign v$G27_5000_out0 = v$A2XNORB2_4670_out0 && v$G28_13602_out0;
assign v$G27_5007_out0 = v$A2XNORB2_4677_out0 && v$G28_13609_out0;
assign v$G27_5011_out0 = v$A2XNORB2_4681_out0 && v$G28_13613_out0;
assign v$G27_5012_out0 = v$A2XNORB2_4682_out0 && v$G28_13614_out0;
assign v$A3$COMP$B3_5166_out0 = v$G7_2442_out0;
assign v$A3$COMP$B3_5178_out0 = v$G7_2444_out0;
assign v$G18_5194_out0 = v$A3XNORB3_15329_out0 && v$G22_13918_out0;
assign v$G18_5198_out0 = v$A3XNORB3_15333_out0 && v$G22_13922_out0;
assign v$G18_5199_out0 = v$A3XNORB3_15334_out0 && v$G22_13923_out0;
assign v$G18_5206_out0 = v$A3XNORB3_15341_out0 && v$G22_13930_out0;
assign v$G18_5210_out0 = v$A3XNORB3_15345_out0 && v$G22_13934_out0;
assign v$G18_5211_out0 = v$A3XNORB3_15346_out0 && v$G22_13935_out0;
assign v$THRESHOLD$WRITE_7550_out0 = v$COUNTEREN_14035_out0;
assign v$THRESHOLD$WRITE_7551_out0 = v$COUNTEREN_14036_out0;
assign v$ENMODE_8055_out0 = v$ENMODE_15175_out0;
assign v$ENMODE_8056_out0 = v$ENMODE_15176_out0;
assign v$RAMADDR_9116_out0 = v$RAMADDR_14184_out0;
assign v$SEL4_9954_out0 = v$B_12696_out0[11:8];
assign v$SEL4_9955_out0 = v$B_12697_out0[11:8];
assign v$SEL4_9956_out0 = v$B_12698_out0[11:8];
assign v$SEL4_9957_out0 = v$B_12699_out0[11:8];
assign v$STRead_10348_out0 = v$G7_8043_out0;
assign v$STRead_10349_out0 = v$G7_8044_out0;
assign v$STClr_10669_out0 = v$G1_17020_out0;
assign v$STClr_10670_out0 = v$G1_17021_out0;
assign v$G19_10700_out0 = v$A4XNORB4_1536_out0 && v$G18_5197_out0;
assign v$G19_10702_out0 = v$A4XNORB4_1538_out0 && v$G18_5209_out0;
assign v$G41_11380_out0 = v$G38_7615_out0 && v$G40_13951_out0;
assign v$G41_11392_out0 = v$G38_7627_out0 && v$G40_13963_out0;
assign v$G14_13227_out0 = v$A4XNORB4_1535_out0 && v$G13_4570_out0;
assign v$G14_13229_out0 = v$A4XNORB4_1537_out0 && v$G13_4582_out0;
assign v$B1_14829_out0 = v$SEL9_11343_out0;
assign v$B1_14830_out0 = v$SEL9_11344_out0;
assign v$B1_14841_out0 = v$SEL9_11355_out0;
assign v$B1_14842_out0 = v$SEL9_11356_out0;
assign v$G24_16288_out0 = v$A3XNORB3_15332_out0 && v$G27_4998_out0;
assign v$G24_16300_out0 = v$A3XNORB3_15344_out0 && v$G27_5010_out0;
assign v$RXRead_16983_out0 = v$G5_8754_out0;
assign v$RXRead_16984_out0 = v$G5_8755_out0;
assign v$B2_17251_out0 = v$SEL8_13491_out0;
assign v$B2_17252_out0 = v$SEL8_13492_out0;
assign v$B2_17263_out0 = v$SEL8_13503_out0;
assign v$B2_17264_out0 = v$SEL8_13504_out0;
assign v$TXWrite_18136_out0 = v$G3_7926_out0;
assign v$TXWrite_18137_out0 = v$G3_7927_out0;
assign v$SEL2_18152_out0 = v$B_12696_out0[7:0];
assign v$SEL2_18153_out0 = v$B_12697_out0[7:0];
assign v$SEL2_18154_out0 = v$B_12698_out0[7:0];
assign v$SEL2_18155_out0 = v$B_12699_out0[7:0];
assign v$B3_18467_out0 = v$SEL7_4331_out0;
assign v$B3_18468_out0 = v$SEL7_4332_out0;
assign v$B3_18479_out0 = v$SEL7_4343_out0;
assign v$B3_18480_out0 = v$SEL7_4344_out0;
assign v$SAME_19345_out0 = v$G41_11383_out0;
assign v$SAME_19347_out0 = v$G41_11384_out0;
assign v$SAME_19348_out0 = v$G41_11385_out0;
assign v$SAME_19361_out0 = v$G41_11395_out0;
assign v$SAME_19363_out0 = v$G41_11396_out0;
assign v$SAME_19364_out0 = v$G41_11397_out0;
assign v$R_1641_out0 = v$VALID_3893_out0;
assign v$R_1644_out0 = v$VALID_3894_out0;
assign v$STATUSREAD_1795_out0 = v$STRead_10348_out0;
assign v$STATUSREAD_1796_out0 = v$STRead_10349_out0;
assign v$A2$COMP$B2_2141_out0 = v$G14_13227_out0;
assign v$A2$COMP$B2_2153_out0 = v$G14_13229_out0;
assign v$OUT_3398_out0 = v$MUX3_2123_out0;
assign v$OUT_3402_out0 = v$MUX3_2127_out0;
assign v$G21_3729_out0 = ! v$B1_14829_out0;
assign v$G21_3730_out0 = ! v$B1_14830_out0;
assign v$G21_3741_out0 = ! v$B1_14841_out0;
assign v$G21_3742_out0 = ! v$B1_14842_out0;
assign v$G8_3914_out0 = !((v$A3_11207_out0 && !v$B3_18467_out0) || (!v$A3_11207_out0) && v$B3_18467_out0);
assign v$G8_3915_out0 = !((v$A3_11208_out0 && !v$B3_18468_out0) || (!v$A3_11208_out0) && v$B3_18468_out0);
assign v$G8_3926_out0 = !((v$A3_11219_out0 && !v$B3_18479_out0) || (!v$A3_11219_out0) && v$B3_18479_out0);
assign v$G8_3927_out0 = !((v$A3_11220_out0 && !v$B3_18480_out0) || (!v$A3_11220_out0) && v$B3_18480_out0);
assign v$G36_6191_out0 = !((v$B3_18467_out0 && !v$A3_11207_out0) || (!v$B3_18467_out0) && v$A3_11207_out0);
assign v$G36_6192_out0 = !((v$B3_18468_out0 && !v$A3_11208_out0) || (!v$B3_18468_out0) && v$A3_11208_out0);
assign v$G36_6203_out0 = !((v$B3_18479_out0 && !v$A3_11219_out0) || (!v$B3_18479_out0) && v$A3_11219_out0);
assign v$G36_6204_out0 = !((v$B3_18480_out0 && !v$A3_11220_out0) || (!v$B3_18480_out0) && v$A3_11220_out0);
assign v$STATUSCLR_6234_out0 = v$STClr_10669_out0;
assign v$STATUSCLR_6235_out0 = v$STClr_10670_out0;
assign v$G6_6790_out0 = ! v$B3_18467_out0;
assign v$G6_6791_out0 = ! v$B3_18468_out0;
assign v$G6_6802_out0 = ! v$B3_18479_out0;
assign v$G6_6803_out0 = ! v$B3_18480_out0;
assign v$G17_8494_out0 = !((v$A0_1892_out0 && !v$B0_3843_out0) || (!v$A0_1892_out0) && v$B0_3843_out0);
assign v$G17_8495_out0 = !((v$A0_1893_out0 && !v$B0_3844_out0) || (!v$A0_1893_out0) && v$B0_3844_out0);
assign v$G17_8506_out0 = !((v$A0_1904_out0 && !v$B0_3855_out0) || (!v$A0_1904_out0) && v$B0_3855_out0);
assign v$G17_8507_out0 = !((v$A0_1905_out0 && !v$B0_3856_out0) || (!v$A0_1905_out0) && v$B0_3856_out0);
assign v$LOWER$SAME_10636_out0 = v$SAME_19348_out0;
assign v$LOWER$SAME_10640_out0 = v$SAME_19364_out0;
assign v$G19_10699_out0 = v$A4XNORB4_1535_out0 && v$G18_5194_out0;
assign v$G19_10701_out0 = v$A4XNORB4_1537_out0 && v$G18_5206_out0;
assign v$TXWRITE_11608_out0 = v$TXWrite_18136_out0;
assign v$TXWRITE_11609_out0 = v$TXWrite_18137_out0;
assign v$G26_11897_out0 = v$A4XNORB4_1536_out0 && v$G24_16288_out0;
assign v$G26_11899_out0 = v$A4XNORB4_1538_out0 && v$G24_16300_out0;
assign v$G23_12747_out0 = ! v$B0_3843_out0;
assign v$G23_12748_out0 = ! v$B0_3844_out0;
assign v$G23_12759_out0 = ! v$B0_3855_out0;
assign v$G23_12760_out0 = ! v$B0_3856_out0;
assign v$A1$COMP$B1_13089_out0 = v$G19_10700_out0;
assign v$A1$COMP$B1_13090_out0 = v$G18_5198_out0;
assign v$A1$COMP$B1_13091_out0 = v$G18_5199_out0;
assign v$A1$COMP$B1_13101_out0 = v$G19_10702_out0;
assign v$A1$COMP$B1_13102_out0 = v$G18_5210_out0;
assign v$A1$COMP$B1_13103_out0 = v$G18_5211_out0;
assign v$G33_13682_out0 = !((v$A0_1892_out0 && !v$B0_3843_out0) || (!v$A0_1892_out0) && v$B0_3843_out0);
assign v$G33_13683_out0 = !((v$A0_1893_out0 && !v$B0_3844_out0) || (!v$A0_1893_out0) && v$B0_3844_out0);
assign v$G33_13694_out0 = !((v$A0_1904_out0 && !v$B0_3855_out0) || (!v$A0_1904_out0) && v$B0_3855_out0);
assign v$G33_13695_out0 = !((v$A0_1905_out0 && !v$B0_3856_out0) || (!v$A0_1905_out0) && v$B0_3856_out0);
assign v$G5_14126_out0 = v$EQUAL_16432_out0 || v$THRESHOLD$WRITE_7550_out0;
assign v$G5_14127_out0 = v$EQUAL_16433_out0 || v$THRESHOLD$WRITE_7551_out0;
assign v$G15_14229_out0 = !((v$A2_8378_out0 && !v$B2_17251_out0) || (!v$A2_8378_out0) && v$B2_17251_out0);
assign v$G15_14230_out0 = !((v$A2_8379_out0 && !v$B2_17252_out0) || (!v$A2_8379_out0) && v$B2_17252_out0);
assign v$G15_14241_out0 = !((v$A2_8390_out0 && !v$B2_17263_out0) || (!v$A2_8390_out0) && v$B2_17263_out0);
assign v$G15_14242_out0 = !((v$A2_8391_out0 && !v$B2_17264_out0) || (!v$A2_8391_out0) && v$B2_17264_out0);
assign v$B_15028_out0 = v$SEL4_9954_out0;
assign v$B_15029_out0 = v$SEL2_18152_out0;
assign v$B_15032_out0 = v$SEL4_9955_out0;
assign v$B_15033_out0 = v$SEL2_18153_out0;
assign v$B_15044_out0 = v$SEL4_9956_out0;
assign v$B_15045_out0 = v$SEL2_18154_out0;
assign v$B_15048_out0 = v$SEL4_9957_out0;
assign v$B_15049_out0 = v$SEL2_18155_out0;
assign v$G35_15129_out0 = !((v$A2_8378_out0 && !v$B2_17251_out0) || (!v$A2_8378_out0) && v$B2_17251_out0);
assign v$G35_15130_out0 = !((v$A2_8379_out0 && !v$B2_17252_out0) || (!v$A2_8379_out0) && v$B2_17252_out0);
assign v$G35_15141_out0 = !((v$A2_8390_out0 && !v$B2_17263_out0) || (!v$A2_8390_out0) && v$B2_17263_out0);
assign v$G35_15142_out0 = !((v$A2_8391_out0 && !v$B2_17264_out0) || (!v$A2_8391_out0) && v$B2_17264_out0);
assign v$MODEWRITE_15321_out0 = v$ModeWrite_4621_out0;
assign v$MODEWRITE_15322_out0 = v$ModeWrite_4622_out0;
assign v$HIGHER$SAME_15641_out0 = v$SAME_19347_out0;
assign v$HIGHER$SAME_15645_out0 = v$SAME_19363_out0;
assign v$G24_16285_out0 = v$A3XNORB3_15329_out0 && v$G27_4995_out0;
assign v$G24_16289_out0 = v$A3XNORB3_15333_out0 && v$G27_4999_out0;
assign v$G24_16290_out0 = v$A3XNORB3_15334_out0 && v$G27_5000_out0;
assign v$G24_16297_out0 = v$A3XNORB3_15341_out0 && v$G27_5007_out0;
assign v$G24_16301_out0 = v$A3XNORB3_15345_out0 && v$G27_5011_out0;
assign v$G24_16302_out0 = v$A3XNORB3_15346_out0 && v$G27_5012_out0;
assign v$RXREAD_16458_out0 = v$RXRead_16983_out0;
assign v$RXREAD_16459_out0 = v$RXRead_16984_out0;
assign v$EN_16500_out0 = v$ENMODE_8055_out0;
assign v$EN_16501_out0 = v$ENMODE_8056_out0;
assign v$G12_17101_out0 = ! v$B2_17251_out0;
assign v$G12_17102_out0 = ! v$B2_17252_out0;
assign v$G12_17113_out0 = ! v$B2_17263_out0;
assign v$G12_17114_out0 = ! v$B2_17264_out0;
assign v$G16_17480_out0 = !((v$A1_14950_out0 && !v$B1_14829_out0) || (!v$A1_14950_out0) && v$B1_14829_out0);
assign v$G16_17481_out0 = !((v$A1_14951_out0 && !v$B1_14830_out0) || (!v$A1_14951_out0) && v$B1_14830_out0);
assign v$G16_17492_out0 = !((v$A1_14962_out0 && !v$B1_14841_out0) || (!v$A1_14962_out0) && v$B1_14841_out0);
assign v$G16_17493_out0 = !((v$A1_14963_out0 && !v$B1_14842_out0) || (!v$A1_14963_out0) && v$B1_14842_out0);
assign v$G34_17938_out0 = !((v$A1_14950_out0 && !v$B1_14829_out0) || (!v$A1_14950_out0) && v$B1_14829_out0);
assign v$G34_17939_out0 = !((v$A1_14951_out0 && !v$B1_14830_out0) || (!v$A1_14951_out0) && v$B1_14830_out0);
assign v$G34_17950_out0 = !((v$A1_14962_out0 && !v$B1_14841_out0) || (!v$A1_14962_out0) && v$B1_14841_out0);
assign v$G34_17951_out0 = !((v$A1_14963_out0 && !v$B1_14842_out0) || (!v$A1_14963_out0) && v$B1_14842_out0);
assign v$SAME_18970_out0 = v$SAME_19345_out0;
assign v$SAME_18974_out0 = v$SAME_19361_out0;
assign v$RAMADDR_19265_out0 = v$RAMADDR_9116_out0;
assign v$SAME_19341_out0 = v$G41_11380_out0;
assign v$SAME_19357_out0 = v$G41_11392_out0;
assign v$A0XNORB0_1590_out0 = v$G17_8494_out0;
assign v$A0XNORB0_1591_out0 = v$G17_8495_out0;
assign v$A0XNORB0_1602_out0 = v$G17_8506_out0;
assign v$A0XNORB0_1603_out0 = v$G17_8507_out0;
assign v$R_1745_out0 = v$R_1641_out0;
assign v$R_1748_out0 = v$R_1644_out0;
assign v$WREN_2730_out0 = v$TXWRITE_11608_out0;
assign v$WREN_2731_out0 = v$TXWRITE_11609_out0;
assign v$SEL7_4324_out0 = v$B_15028_out0[3:3];
assign v$SEL7_4327_out0 = v$B_15032_out0[3:3];
assign v$SEL7_4336_out0 = v$B_15044_out0[3:3];
assign v$SEL7_4339_out0 = v$B_15048_out0[3:3];
assign v$G1_4372_out0 = v$STATUSREAD_1795_out0 || v$RXREAD_16458_out0;
assign v$G1_4373_out0 = v$STATUSREAD_1796_out0 || v$RXREAD_16459_out0;
assign v$IN_4526_out0 = v$OUT_3398_out0;
assign v$IN_4530_out0 = v$OUT_3402_out0;
assign v$A2XNORB2_4666_out0 = v$G15_14229_out0;
assign v$A2XNORB2_4667_out0 = v$G15_14230_out0;
assign v$A2XNORB2_4678_out0 = v$G15_14241_out0;
assign v$A2XNORB2_4679_out0 = v$G15_14242_out0;
assign v$RXreset_6240_out0 = v$RXREAD_16458_out0;
assign v$RXreset_6241_out0 = v$RXREAD_16459_out0;
assign v$G5_7222_out0 = v$A3_11207_out0 && v$G6_6790_out0;
assign v$G5_7223_out0 = v$A3_11208_out0 && v$G6_6791_out0;
assign v$G5_7234_out0 = v$A3_11219_out0 && v$G6_6802_out0;
assign v$G5_7235_out0 = v$A3_11220_out0 && v$G6_6803_out0;
assign v$_7595_out0 = v$RAMADDR_19265_out0[3:0];
assign v$_7595_out1 = v$RAMADDR_19265_out0[11:8];
assign v$G38_7616_out0 = v$G33_13682_out0 && v$G34_17938_out0;
assign v$G38_7617_out0 = v$G33_13683_out0 && v$G34_17939_out0;
assign v$G38_7628_out0 = v$G33_13694_out0 && v$G34_17950_out0;
assign v$G38_7629_out0 = v$G33_13695_out0 && v$G34_17951_out0;
assign v$A0$COMP$B0_8312_out0 = v$G26_11897_out0;
assign v$A0$COMP$B0_8313_out0 = v$G24_16289_out0;
assign v$A0$COMP$B0_8314_out0 = v$G24_16290_out0;
assign v$A0$COMP$B0_8324_out0 = v$G26_11899_out0;
assign v$A0$COMP$B0_8325_out0 = v$G24_16301_out0;
assign v$A0$COMP$B0_8326_out0 = v$G24_16302_out0;
assign v$SEL3_9373_out0 = v$B_15029_out0[7:4];
assign v$SEL3_9374_out0 = v$B_15033_out0[7:4];
assign v$SEL3_9377_out0 = v$B_15045_out0[7:4];
assign v$SEL3_9378_out0 = v$B_15049_out0[7:4];
assign v$G1_9762_out0 = v$LOWER$SAME_10636_out0 && v$HIGHER$SAME_15641_out0;
assign v$G1_9766_out0 = v$LOWER$SAME_10640_out0 && v$HIGHER$SAME_15645_out0;
assign v$G20_10310_out0 = v$A1_14950_out0 && v$G21_3729_out0;
assign v$G20_10311_out0 = v$A1_14951_out0 && v$G21_3730_out0;
assign v$G20_10322_out0 = v$A1_14962_out0 && v$G21_3741_out0;
assign v$G20_10323_out0 = v$A1_14963_out0 && v$G21_3742_out0;
assign v$SEL9_11336_out0 = v$B_15028_out0[1:1];
assign v$SEL9_11339_out0 = v$B_15032_out0[1:1];
assign v$SEL9_11348_out0 = v$B_15044_out0[1:1];
assign v$SEL9_11351_out0 = v$B_15048_out0[1:1];
assign v$G25_11446_out0 = v$A0_1892_out0 && v$G23_12747_out0;
assign v$G25_11447_out0 = v$A0_1893_out0 && v$G23_12748_out0;
assign v$G25_11458_out0 = v$A0_1904_out0 && v$G23_12759_out0;
assign v$G25_11459_out0 = v$A0_1905_out0 && v$G23_12760_out0;
assign v$G26_11896_out0 = v$A4XNORB4_1535_out0 && v$G24_16285_out0;
assign v$G26_11898_out0 = v$A4XNORB4_1537_out0 && v$G24_16297_out0;
assign v$A1$COMP$B1_13086_out0 = v$G19_10699_out0;
assign v$A1$COMP$B1_13098_out0 = v$G19_10701_out0;
assign v$SEL10_13189_out0 = v$B_15028_out0[0:0];
assign v$SEL10_13192_out0 = v$B_15032_out0[0:0];
assign v$SEL10_13201_out0 = v$B_15044_out0[0:0];
assign v$SEL10_13204_out0 = v$B_15048_out0[0:0];
assign v$Clear_13319_out0 = v$STATUSCLR_6234_out0;
assign v$Clear_13320_out0 = v$STATUSCLR_6235_out0;
assign v$SEL8_13484_out0 = v$B_15028_out0[2:2];
assign v$SEL8_13487_out0 = v$B_15032_out0[2:2];
assign v$SEL8_13496_out0 = v$B_15044_out0[2:2];
assign v$SEL8_13499_out0 = v$B_15048_out0[2:2];
assign v$G40_13952_out0 = v$G35_15129_out0 && v$G36_6191_out0;
assign v$G40_13953_out0 = v$G35_15130_out0 && v$G36_6192_out0;
assign v$G40_13964_out0 = v$G35_15141_out0 && v$G36_6203_out0;
assign v$G40_13965_out0 = v$G35_15142_out0 && v$G36_6204_out0;
assign v$TXSet_14941_out0 = v$TXWRITE_11608_out0;
assign v$TXSet_14942_out0 = v$TXWRITE_11609_out0;
assign v$A3XNORB3_15330_out0 = v$G8_3914_out0;
assign v$A3XNORB3_15331_out0 = v$G8_3915_out0;
assign v$A3XNORB3_15342_out0 = v$G8_3926_out0;
assign v$A3XNORB3_15343_out0 = v$G8_3927_out0;
assign v$G11_16237_out0 = v$A2_8378_out0 && v$G12_17101_out0;
assign v$G11_16238_out0 = v$A2_8379_out0 && v$G12_17102_out0;
assign v$G11_16249_out0 = v$A2_8390_out0 && v$G12_17113_out0;
assign v$G11_16250_out0 = v$A2_8391_out0 && v$G12_17114_out0;
assign v$A1XNORB1_16666_out0 = v$G16_17480_out0;
assign v$A1XNORB1_16667_out0 = v$G16_17481_out0;
assign v$A1XNORB1_16678_out0 = v$G16_17492_out0;
assign v$A1XNORB1_16679_out0 = v$G16_17493_out0;
assign v$SEL2_18082_out0 = v$B_15029_out0[3:0];
assign v$SEL2_18083_out0 = v$B_15033_out0[3:0];
assign v$SEL2_18086_out0 = v$B_15045_out0[3:0];
assign v$SEL2_18087_out0 = v$B_15049_out0[3:0];
assign v$MUX1_18934_out0 = v$G5_14126_out0 ? v$C3_12770_out0 : v$A1_14282_out0;
assign v$MUX1_18935_out0 = v$G5_14127_out0 ? v$C3_12771_out0 : v$A1_14283_out0;
assign v$SAME_18968_out0 = v$SAME_19341_out0;
assign v$SAME_18972_out0 = v$SAME_19357_out0;
assign v$G32_420_out0 = v$A1$COMP$B1_13089_out0 || v$A0$COMP$B0_8312_out0;
assign v$G32_421_out0 = v$A1$COMP$B1_13090_out0 || v$A0$COMP$B0_8313_out0;
assign v$G32_422_out0 = v$A1$COMP$B1_13091_out0 || v$A0$COMP$B0_8314_out0;
assign v$G32_432_out0 = v$A1$COMP$B1_13101_out0 || v$A0$COMP$B0_8324_out0;
assign v$G32_433_out0 = v$A1$COMP$B1_13102_out0 || v$A0$COMP$B0_8325_out0;
assign v$G32_434_out0 = v$A1$COMP$B1_13103_out0 || v$A0$COMP$B0_8326_out0;
assign v$SEL8_2132_out0 = v$_7595_out1[7:7];
assign v$SEL3_3340_out0 = v$_7595_out1[2:2];
assign v$B0_3836_out0 = v$SEL10_13189_out0;
assign v$B0_3839_out0 = v$SEL10_13192_out0;
assign v$B0_3848_out0 = v$SEL10_13201_out0;
assign v$B0_3851_out0 = v$SEL10_13204_out0;
assign v$G13_4571_out0 = v$A3XNORB3_15330_out0 && v$G11_16237_out0;
assign v$G13_4572_out0 = v$A3XNORB3_15331_out0 && v$G11_16238_out0;
assign v$G13_4583_out0 = v$A3XNORB3_15342_out0 && v$G11_16249_out0;
assign v$G13_4584_out0 = v$A3XNORB3_15343_out0 && v$G11_16250_out0;
assign v$A3$COMP$B3_5167_out0 = v$G5_7222_out0;
assign v$A3$COMP$B3_5168_out0 = v$G5_7223_out0;
assign v$A3$COMP$B3_5179_out0 = v$G5_7234_out0;
assign v$A3$COMP$B3_5180_out0 = v$G5_7235_out0;
assign v$SEL1_7288_out0 = v$_7595_out1[0:0];
assign v$A0$COMP$B0_8309_out0 = v$G26_11896_out0;
assign v$A0$COMP$B0_8321_out0 = v$G26_11898_out0;
assign v$IN_9948_out0 = v$IN_4526_out0;
assign v$IN_9952_out0 = v$IN_4530_out0;
assign v$G41_11381_out0 = v$G38_7616_out0 && v$G40_13952_out0;
assign v$G41_11382_out0 = v$G38_7617_out0 && v$G40_13953_out0;
assign v$G41_11393_out0 = v$G38_7628_out0 && v$G40_13964_out0;
assign v$G41_11394_out0 = v$G38_7629_out0 && v$G40_13965_out0;
assign v$WREN_11505_out0 = v$WREN_2730_out0;
assign v$WREN_11506_out0 = v$WREN_2731_out0;
assign v$SEL5_12186_out0 = v$_7595_out1[4:4];
assign v$TXSet_13235_out0 = v$TXSet_14941_out0;
assign v$TXSet_13236_out0 = v$TXSet_14942_out0;
assign v$G28_13598_out0 = v$A1XNORB1_16666_out0 && v$G25_11446_out0;
assign v$G28_13599_out0 = v$A1XNORB1_16667_out0 && v$G25_11447_out0;
assign v$G28_13610_out0 = v$A1XNORB1_16678_out0 && v$G25_11458_out0;
assign v$G28_13611_out0 = v$A1XNORB1_16679_out0 && v$G25_11459_out0;
assign v$G22_13919_out0 = v$A2XNORB2_4666_out0 && v$G20_10310_out0;
assign v$G22_13920_out0 = v$A2XNORB2_4667_out0 && v$G20_10311_out0;
assign v$G22_13931_out0 = v$A2XNORB2_4678_out0 && v$G20_10322_out0;
assign v$G22_13932_out0 = v$A2XNORB2_4679_out0 && v$G20_10323_out0;
assign v$B1_14822_out0 = v$SEL9_11336_out0;
assign v$B1_14825_out0 = v$SEL9_11339_out0;
assign v$B1_14834_out0 = v$SEL9_11348_out0;
assign v$B1_14837_out0 = v$SEL9_11351_out0;
assign v$SEL6_14846_out0 = v$_7595_out1[5:5];
assign v$B_15030_out0 = v$SEL3_9373_out0;
assign v$B_15031_out0 = v$SEL2_18082_out0;
assign v$B_15034_out0 = v$SEL3_9374_out0;
assign v$B_15035_out0 = v$SEL2_18083_out0;
assign v$B_15046_out0 = v$SEL3_9377_out0;
assign v$B_15047_out0 = v$SEL2_18086_out0;
assign v$B_15050_out0 = v$SEL3_9378_out0;
assign v$B_15051_out0 = v$SEL2_18087_out0;
assign v$Clear_15245_out0 = v$Clear_13319_out0;
assign v$Clear_15246_out0 = v$Clear_13320_out0;
assign v$USELESS_16072_out0 = v$_7595_out0;
assign v$SEL2_16440_out0 = v$_7595_out1[1:1];
assign v$SEL4_17042_out0 = v$_7595_out1[3:3];
assign v$B2_17244_out0 = v$SEL8_13484_out0;
assign v$B2_17247_out0 = v$SEL8_13487_out0;
assign v$B2_17256_out0 = v$SEL8_13496_out0;
assign v$B2_17259_out0 = v$SEL8_13499_out0;
assign v$SEL7_17604_out0 = v$_7595_out1[6:6];
assign v$G3_18295_out0 = ! v$R_1745_out0;
assign v$G3_18298_out0 = ! v$R_1748_out0;
assign v$B3_18460_out0 = v$SEL7_4324_out0;
assign v$B3_18463_out0 = v$SEL7_4327_out0;
assign v$B3_18472_out0 = v$SEL7_4336_out0;
assign v$B3_18475_out0 = v$SEL7_4339_out0;
assign v$G18_18705_out0 = v$WREN_2730_out0 || v$G19_8570_out0;
assign v$G18_18706_out0 = v$WREN_2731_out0 || v$G19_8571_out0;
assign v$R_18943_out0 = v$RXreset_6240_out0;
assign v$R_18954_out0 = v$RXreset_6241_out0;
assign v$SAME_19346_out0 = v$G1_9762_out0;
assign v$SAME_19362_out0 = v$G1_9766_out0;
assign v$G32_417_out0 = v$A1$COMP$B1_13086_out0 || v$A0$COMP$B0_8309_out0;
assign v$G32_429_out0 = v$A1$COMP$B1_13098_out0 || v$A0$COMP$B0_8321_out0;
assign v$_1709_out0 = v$IN_9948_out0[15:15];
assign v$_1710_out0 = v$IN_9952_out0[15:15];
assign v$A2$COMP$B2_2142_out0 = v$G13_4571_out0;
assign v$A2$COMP$B2_2143_out0 = v$G13_4572_out0;
assign v$A2$COMP$B2_2154_out0 = v$G13_4583_out0;
assign v$A2$COMP$B2_2155_out0 = v$G13_4584_out0;
assign v$G21_3722_out0 = ! v$B1_14822_out0;
assign v$G21_3725_out0 = ! v$B1_14825_out0;
assign v$G21_3734_out0 = ! v$B1_14834_out0;
assign v$G21_3737_out0 = ! v$B1_14837_out0;
assign v$G8_3907_out0 = !((v$A3_11200_out0 && !v$B3_18460_out0) || (!v$A3_11200_out0) && v$B3_18460_out0);
assign v$G8_3910_out0 = !((v$A3_11203_out0 && !v$B3_18463_out0) || (!v$A3_11203_out0) && v$B3_18463_out0);
assign v$G8_3919_out0 = !((v$A3_11212_out0 && !v$B3_18472_out0) || (!v$A3_11212_out0) && v$B3_18472_out0);
assign v$G8_3922_out0 = !((v$A3_11215_out0 && !v$B3_18475_out0) || (!v$A3_11215_out0) && v$B3_18475_out0);
assign v$SEL7_4325_out0 = v$B_15030_out0[3:3];
assign v$SEL7_4326_out0 = v$B_15031_out0[3:3];
assign v$SEL7_4328_out0 = v$B_15034_out0[3:3];
assign v$SEL7_4329_out0 = v$B_15035_out0[3:3];
assign v$SEL7_4337_out0 = v$B_15046_out0[3:3];
assign v$SEL7_4338_out0 = v$B_15047_out0[3:3];
assign v$SEL7_4340_out0 = v$B_15050_out0[3:3];
assign v$SEL7_4341_out0 = v$B_15051_out0[3:3];
assign v$G27_4996_out0 = v$A2XNORB2_4666_out0 && v$G28_13598_out0;
assign v$G27_4997_out0 = v$A2XNORB2_4667_out0 && v$G28_13599_out0;
assign v$G27_5008_out0 = v$A2XNORB2_4678_out0 && v$G28_13610_out0;
assign v$G27_5009_out0 = v$A2XNORB2_4679_out0 && v$G28_13611_out0;
assign v$_5015_out0 = v$IN_9948_out0[11:0];
assign v$_5019_out0 = v$IN_9952_out0[11:0];
assign v$G18_5195_out0 = v$A3XNORB3_15330_out0 && v$G22_13919_out0;
assign v$G18_5196_out0 = v$A3XNORB3_15331_out0 && v$G22_13920_out0;
assign v$G18_5207_out0 = v$A3XNORB3_15342_out0 && v$G22_13931_out0;
assign v$G18_5208_out0 = v$A3XNORB3_15343_out0 && v$G22_13932_out0;
assign v$G3_5216_out0 = v$SEL5_12186_out0 && v$SEL6_14846_out0;
assign v$G36_6184_out0 = !((v$B3_18460_out0 && !v$A3_11200_out0) || (!v$B3_18460_out0) && v$A3_11200_out0);
assign v$G36_6187_out0 = !((v$B3_18463_out0 && !v$A3_11203_out0) || (!v$B3_18463_out0) && v$A3_11203_out0);
assign v$G36_6196_out0 = !((v$B3_18472_out0 && !v$A3_11212_out0) || (!v$B3_18472_out0) && v$A3_11212_out0);
assign v$G36_6199_out0 = !((v$B3_18475_out0 && !v$A3_11215_out0) || (!v$B3_18475_out0) && v$A3_11215_out0);
assign v$G4_6660_out0 = v$SEL7_17604_out0 && v$SEL8_2132_out0;
assign v$G6_6783_out0 = ! v$B3_18460_out0;
assign v$G6_6786_out0 = ! v$B3_18463_out0;
assign v$G6_6795_out0 = ! v$B3_18472_out0;
assign v$G6_6798_out0 = ! v$B3_18475_out0;
assign v$_7691_out0 = v$IN_9948_out0[3:0];
assign v$_7692_out0 = v$IN_9952_out0[3:0];
assign v$ShiftEN_8039_out0 = v$G18_18705_out0;
assign v$ShiftEN_8040_out0 = v$G18_18706_out0;
assign v$G17_8487_out0 = !((v$A0_1885_out0 && !v$B0_3836_out0) || (!v$A0_1885_out0) && v$B0_3836_out0);
assign v$G17_8490_out0 = !((v$A0_1888_out0 && !v$B0_3839_out0) || (!v$A0_1888_out0) && v$B0_3839_out0);
assign v$G17_8499_out0 = !((v$A0_1897_out0 && !v$B0_3848_out0) || (!v$A0_1897_out0) && v$B0_3848_out0);
assign v$G17_8502_out0 = !((v$A0_1900_out0 && !v$B0_3851_out0) || (!v$A0_1900_out0) && v$B0_3851_out0);
assign v$G9_9018_out0 = v$TXSet_13235_out0 && v$TXLast_11914_out0;
assign v$G9_9019_out0 = v$TXSet_13236_out0 && v$TXLast_11915_out0;
assign v$G17_9229_out0 = ! v$WREN_11505_out0;
assign v$G17_9230_out0 = ! v$WREN_11506_out0;
assign v$SEL9_11337_out0 = v$B_15030_out0[1:1];
assign v$SEL9_11338_out0 = v$B_15031_out0[1:1];
assign v$SEL9_11340_out0 = v$B_15034_out0[1:1];
assign v$SEL9_11341_out0 = v$B_15035_out0[1:1];
assign v$SEL9_11349_out0 = v$B_15046_out0[1:1];
assign v$SEL9_11350_out0 = v$B_15047_out0[1:1];
assign v$SEL9_11352_out0 = v$B_15050_out0[1:1];
assign v$SEL9_11353_out0 = v$B_15051_out0[1:1];
assign v$G2_12265_out0 = v$SEL3_3340_out0 && v$SEL4_17042_out0;
assign v$G23_12740_out0 = ! v$B0_3836_out0;
assign v$G23_12743_out0 = ! v$B0_3839_out0;
assign v$G23_12752_out0 = ! v$B0_3848_out0;
assign v$G23_12755_out0 = ! v$B0_3851_out0;
assign v$SEL10_13190_out0 = v$B_15030_out0[0:0];
assign v$SEL10_13191_out0 = v$B_15031_out0[0:0];
assign v$SEL10_13193_out0 = v$B_15034_out0[0:0];
assign v$SEL10_13194_out0 = v$B_15035_out0[0:0];
assign v$SEL10_13202_out0 = v$B_15046_out0[0:0];
assign v$SEL10_13203_out0 = v$B_15047_out0[0:0];
assign v$SEL10_13205_out0 = v$B_15050_out0[0:0];
assign v$SEL10_13206_out0 = v$B_15051_out0[0:0];
assign v$SEL8_13485_out0 = v$B_15030_out0[2:2];
assign v$SEL8_13486_out0 = v$B_15031_out0[2:2];
assign v$SEL8_13488_out0 = v$B_15034_out0[2:2];
assign v$SEL8_13489_out0 = v$B_15035_out0[2:2];
assign v$SEL8_13497_out0 = v$B_15046_out0[2:2];
assign v$SEL8_13498_out0 = v$B_15047_out0[2:2];
assign v$SEL8_13500_out0 = v$B_15050_out0[2:2];
assign v$SEL8_13501_out0 = v$B_15051_out0[2:2];
assign v$G1_13556_out0 = v$STATE_16626_out0 && v$G3_18295_out0;
assign v$G1_13559_out0 = v$STATE_16629_out0 && v$G3_18298_out0;
assign v$G33_13675_out0 = !((v$A0_1885_out0 && !v$B0_3836_out0) || (!v$A0_1885_out0) && v$B0_3836_out0);
assign v$G33_13678_out0 = !((v$A0_1888_out0 && !v$B0_3839_out0) || (!v$A0_1888_out0) && v$B0_3839_out0);
assign v$G33_13687_out0 = !((v$A0_1897_out0 && !v$B0_3848_out0) || (!v$A0_1897_out0) && v$B0_3848_out0);
assign v$G33_13690_out0 = !((v$A0_1900_out0 && !v$B0_3851_out0) || (!v$A0_1900_out0) && v$B0_3851_out0);
assign v$_13854_out0 = v$IN_9948_out0[3:0];
assign v$_13857_out0 = v$IN_9952_out0[3:0];
assign v$G15_14222_out0 = !((v$A2_8371_out0 && !v$B2_17244_out0) || (!v$A2_8371_out0) && v$B2_17244_out0);
assign v$G15_14225_out0 = !((v$A2_8374_out0 && !v$B2_17247_out0) || (!v$A2_8374_out0) && v$B2_17247_out0);
assign v$G15_14234_out0 = !((v$A2_8383_out0 && !v$B2_17256_out0) || (!v$A2_8383_out0) && v$B2_17256_out0);
assign v$G15_14237_out0 = !((v$A2_8386_out0 && !v$B2_17259_out0) || (!v$A2_8386_out0) && v$B2_17259_out0);
assign v$G1_15015_out0 = v$SEL1_7288_out0 && v$SEL2_16440_out0;
assign v$G35_15122_out0 = !((v$A2_8371_out0 && !v$B2_17244_out0) || (!v$A2_8371_out0) && v$B2_17244_out0);
assign v$G35_15125_out0 = !((v$A2_8374_out0 && !v$B2_17247_out0) || (!v$A2_8374_out0) && v$B2_17247_out0);
assign v$G35_15134_out0 = !((v$A2_8383_out0 && !v$B2_17256_out0) || (!v$A2_8383_out0) && v$B2_17256_out0);
assign v$G35_15137_out0 = !((v$A2_8386_out0 && !v$B2_17259_out0) || (!v$A2_8386_out0) && v$B2_17259_out0);
assign v$_15203_out0 = v$IN_9948_out0[15:4];
assign v$_15207_out0 = v$IN_9952_out0[15:4];
assign v$_15239_out0 = v$IN_9948_out0[15:4];
assign v$_15243_out0 = v$IN_9952_out0[15:4];
assign v$G31_16106_out0 = v$A2$COMP$B2_2144_out0 || v$G32_420_out0;
assign v$G31_16107_out0 = v$A2$COMP$B2_2145_out0 || v$G32_421_out0;
assign v$G31_16108_out0 = v$A2$COMP$B2_2146_out0 || v$G32_422_out0;
assign v$G31_16118_out0 = v$A2$COMP$B2_2156_out0 || v$G32_432_out0;
assign v$G31_16119_out0 = v$A2$COMP$B2_2157_out0 || v$G32_433_out0;
assign v$G31_16120_out0 = v$A2$COMP$B2_2158_out0 || v$G32_434_out0;
assign v$G6_16158_out0 = ! v$R_18943_out0;
assign v$G6_16169_out0 = ! v$R_18954_out0;
assign v$G12_17094_out0 = ! v$B2_17244_out0;
assign v$G12_17097_out0 = ! v$B2_17247_out0;
assign v$G12_17106_out0 = ! v$B2_17256_out0;
assign v$G12_17109_out0 = ! v$B2_17259_out0;
assign v$_17370_out0 = v$IN_9948_out0[15:4];
assign v$_17374_out0 = v$IN_9952_out0[15:4];
assign v$G16_17473_out0 = !((v$A1_14943_out0 && !v$B1_14822_out0) || (!v$A1_14943_out0) && v$B1_14822_out0);
assign v$G16_17476_out0 = !((v$A1_14946_out0 && !v$B1_14825_out0) || (!v$A1_14946_out0) && v$B1_14825_out0);
assign v$G16_17485_out0 = !((v$A1_14955_out0 && !v$B1_14834_out0) || (!v$A1_14955_out0) && v$B1_14834_out0);
assign v$G16_17488_out0 = !((v$A1_14958_out0 && !v$B1_14837_out0) || (!v$A1_14958_out0) && v$B1_14837_out0);
assign v$S_17543_out0 = v$TXSet_13235_out0;
assign v$S_17554_out0 = v$TXSet_13236_out0;
assign v$G34_17931_out0 = !((v$A1_14943_out0 && !v$B1_14822_out0) || (!v$A1_14943_out0) && v$B1_14822_out0);
assign v$G34_17934_out0 = !((v$A1_14946_out0 && !v$B1_14825_out0) || (!v$A1_14946_out0) && v$B1_14825_out0);
assign v$G34_17943_out0 = !((v$A1_14955_out0 && !v$B1_14834_out0) || (!v$A1_14955_out0) && v$B1_14834_out0);
assign v$G34_17946_out0 = !((v$A1_14958_out0 && !v$B1_14837_out0) || (!v$A1_14958_out0) && v$B1_14837_out0);
assign v$R_18944_out0 = v$Clear_15245_out0;
assign v$R_18945_out0 = v$Clear_15245_out0;
assign v$R_18946_out0 = v$Clear_15245_out0;
assign v$R_18955_out0 = v$Clear_15246_out0;
assign v$R_18956_out0 = v$Clear_15246_out0;
assign v$R_18957_out0 = v$Clear_15246_out0;
assign v$SAME_18971_out0 = v$SAME_19346_out0;
assign v$SAME_18975_out0 = v$SAME_19362_out0;
assign v$SAME_19343_out0 = v$G41_11381_out0;
assign v$SAME_19344_out0 = v$G41_11382_out0;
assign v$SAME_19359_out0 = v$G41_11393_out0;
assign v$SAME_19360_out0 = v$G41_11394_out0;
assign v$MUX1_435_out0 = v$G17_9229_out0 ? v$FF2_3160_out0 : v$_3685_out0;
assign v$MUX1_436_out0 = v$G17_9230_out0 ? v$FF2_3161_out0 : v$_3686_out0;
assign v$G5_1268_out0 = v$FF2_13622_out0 && v$G6_16158_out0;
assign v$G5_1273_out0 = v$FF2_13633_out0 && v$G6_16169_out0;
assign v$A0XNORB0_1583_out0 = v$G17_8487_out0;
assign v$A0XNORB0_1586_out0 = v$G17_8490_out0;
assign v$A0XNORB0_1595_out0 = v$G17_8499_out0;
assign v$A0XNORB0_1598_out0 = v$G17_8502_out0;
assign v$_1631_out0 = { v$C1_8289_out0,v$_5015_out0 };
assign v$_1635_out0 = { v$C1_8293_out0,v$_5019_out0 };
assign v$MUX8_1651_out0 = v$G17_9229_out0 ? v$C1_13423_out0 : v$_9743_out1;
assign v$MUX8_1652_out0 = v$G17_9230_out0 ? v$C1_13424_out0 : v$_9744_out1;
assign v$G30_1939_out0 = v$A3$COMP$B3_5169_out0 || v$G31_16106_out0;
assign v$G30_1940_out0 = v$A3$COMP$B3_5170_out0 || v$G31_16107_out0;
assign v$G30_1941_out0 = v$A3$COMP$B3_5171_out0 || v$G31_16108_out0;
assign v$G30_1951_out0 = v$A3$COMP$B3_5181_out0 || v$G31_16118_out0;
assign v$G30_1952_out0 = v$A3$COMP$B3_5182_out0 || v$G31_16119_out0;
assign v$G30_1953_out0 = v$A3$COMP$B3_5183_out0 || v$G31_16120_out0;
assign v$B0_3837_out0 = v$SEL10_13190_out0;
assign v$B0_3838_out0 = v$SEL10_13191_out0;
assign v$B0_3840_out0 = v$SEL10_13193_out0;
assign v$B0_3841_out0 = v$SEL10_13194_out0;
assign v$B0_3849_out0 = v$SEL10_13202_out0;
assign v$B0_3850_out0 = v$SEL10_13203_out0;
assign v$B0_3852_out0 = v$SEL10_13205_out0;
assign v$B0_3853_out0 = v$SEL10_13206_out0;
assign v$A2XNORB2_4659_out0 = v$G15_14222_out0;
assign v$A2XNORB2_4662_out0 = v$G15_14225_out0;
assign v$A2XNORB2_4671_out0 = v$G15_14234_out0;
assign v$A2XNORB2_4674_out0 = v$G15_14237_out0;
assign v$G5_6084_out0 = v$G1_15015_out0 && v$G2_12265_out0;
assign v$G5_7215_out0 = v$A3_11200_out0 && v$G6_6783_out0;
assign v$G5_7218_out0 = v$A3_11203_out0 && v$G6_6786_out0;
assign v$G5_7227_out0 = v$A3_11212_out0 && v$G6_6795_out0;
assign v$G5_7230_out0 = v$A3_11215_out0 && v$G6_6798_out0;
assign v$G38_7609_out0 = v$G33_13675_out0 && v$G34_17931_out0;
assign v$G38_7612_out0 = v$G33_13678_out0 && v$G34_17934_out0;
assign v$G38_7621_out0 = v$G33_13687_out0 && v$G34_17943_out0;
assign v$G38_7624_out0 = v$G33_13690_out0 && v$G34_17946_out0;
assign v$G2_7901_out0 = v$G1_13556_out0 || v$S_8337_out0;
assign v$G2_7904_out0 = v$G1_13559_out0 || v$S_8340_out0;
assign v$MUX6_9458_out0 = v$G17_9229_out0 ? v$FF7_18731_out0 : v$_8404_out1;
assign v$MUX6_9459_out0 = v$G17_9230_out0 ? v$FF7_18732_out0 : v$_8405_out1;
assign v$_9821_out0 = { v$_17370_out0,v$LSBS_15901_out0 };
assign v$_9825_out0 = { v$_17374_out0,v$LSBS_15902_out0 };
assign v$MUX7_9855_out0 = v$G17_9229_out0 ? v$FF8_8346_out0 : v$_9743_out0;
assign v$MUX7_9856_out0 = v$G17_9230_out0 ? v$FF8_8347_out0 : v$_9744_out0;
assign v$G20_10303_out0 = v$A1_14943_out0 && v$G21_3722_out0;
assign v$G20_10306_out0 = v$A1_14946_out0 && v$G21_3725_out0;
assign v$G20_10315_out0 = v$A1_14955_out0 && v$G21_3734_out0;
assign v$G20_10318_out0 = v$A1_14958_out0 && v$G21_3737_out0;
assign v$_10333_out0 = { v$_1709_out0,v$_1709_out0 };
assign v$_10334_out0 = { v$_1710_out0,v$_1710_out0 };
assign v$LOWER$SAME_10635_out0 = v$SAME_19344_out0;
assign v$LOWER$SAME_10639_out0 = v$SAME_19360_out0;
assign v$G25_11439_out0 = v$A0_1885_out0 && v$G23_12740_out0;
assign v$G25_11442_out0 = v$A0_1888_out0 && v$G23_12743_out0;
assign v$G25_11451_out0 = v$A0_1897_out0 && v$G23_12752_out0;
assign v$G25_11454_out0 = v$A0_1900_out0 && v$G23_12755_out0;
assign v$MUX4_12210_out0 = v$IS$32$BITS_3203_out0 ? v$SAME_18971_out0 : v$SAME_18970_out0;
assign v$MUX4_12211_out0 = v$IS$32$BITS_3204_out0 ? v$SAME_18975_out0 : v$SAME_18974_out0;
assign v$G4_12405_out0 = v$G5_1267_out0 || v$S_17543_out0;
assign v$G4_12410_out0 = v$G5_1272_out0 || v$S_17554_out0;
assign v$A1$COMP$B1_13087_out0 = v$G18_5195_out0;
assign v$A1$COMP$B1_13088_out0 = v$G18_5196_out0;
assign v$A1$COMP$B1_13099_out0 = v$G18_5207_out0;
assign v$A1$COMP$B1_13100_out0 = v$G18_5208_out0;
assign v$MUX2_13871_out0 = v$G17_9229_out0 ? v$FF3_271_out0 : v$_3685_out1;
assign v$MUX2_13872_out0 = v$G17_9230_out0 ? v$FF3_272_out0 : v$_3686_out1;
assign v$_13892_out0 = { v$_15203_out0,v$_13854_out0 };
assign v$_13896_out0 = { v$_15207_out0,v$_13857_out0 };
assign v$G40_13945_out0 = v$G35_15122_out0 && v$G36_6184_out0;
assign v$G40_13948_out0 = v$G35_15125_out0 && v$G36_6187_out0;
assign v$G40_13957_out0 = v$G35_15134_out0 && v$G36_6196_out0;
assign v$G40_13960_out0 = v$G35_15137_out0 && v$G36_6199_out0;
assign v$B1_14823_out0 = v$SEL9_11337_out0;
assign v$B1_14824_out0 = v$SEL9_11338_out0;
assign v$B1_14826_out0 = v$SEL9_11340_out0;
assign v$B1_14827_out0 = v$SEL9_11341_out0;
assign v$B1_14835_out0 = v$SEL9_11349_out0;
assign v$B1_14836_out0 = v$SEL9_11350_out0;
assign v$B1_14838_out0 = v$SEL9_11352_out0;
assign v$B1_14839_out0 = v$SEL9_11353_out0;
assign v$MUX5_15088_out0 = v$S_10809_out0 ? v$_7691_out0 : v$C1_13395_out0;
assign v$MUX5_15089_out0 = v$S_10810_out0 ? v$_7692_out0 : v$C1_13396_out0;
assign v$A3XNORB3_15323_out0 = v$G8_3907_out0;
assign v$A3XNORB3_15326_out0 = v$G8_3910_out0;
assign v$A3XNORB3_15335_out0 = v$G8_3919_out0;
assign v$A3XNORB3_15338_out0 = v$G8_3922_out0;
assign v$HIGHER$SAME_15640_out0 = v$SAME_19343_out0;
assign v$HIGHER$SAME_15644_out0 = v$SAME_19359_out0;
assign v$G31_16103_out0 = v$A2$COMP$B2_2141_out0 || v$G32_417_out0;
assign v$G31_16115_out0 = v$A2$COMP$B2_2153_out0 || v$G32_429_out0;
assign v$G6_16159_out0 = ! v$R_18944_out0;
assign v$G6_16160_out0 = ! v$R_18945_out0;
assign v$G6_16161_out0 = ! v$R_18946_out0;
assign v$G6_16170_out0 = ! v$R_18955_out0;
assign v$G6_16171_out0 = ! v$R_18956_out0;
assign v$G6_16172_out0 = ! v$R_18957_out0;
assign v$MUX4_16228_out0 = v$G17_9229_out0 ? v$FF5_16956_out0 : v$_14689_out1;
assign v$MUX4_16229_out0 = v$G17_9230_out0 ? v$FF5_16957_out0 : v$_14690_out1;
assign v$G11_16230_out0 = v$A2_8371_out0 && v$G12_17094_out0;
assign v$G11_16233_out0 = v$A2_8374_out0 && v$G12_17097_out0;
assign v$G11_16242_out0 = v$A2_8383_out0 && v$G12_17106_out0;
assign v$G11_16245_out0 = v$A2_8386_out0 && v$G12_17109_out0;
assign v$G24_16286_out0 = v$A3XNORB3_15330_out0 && v$G27_4996_out0;
assign v$G24_16287_out0 = v$A3XNORB3_15331_out0 && v$G27_4997_out0;
assign v$G24_16298_out0 = v$A3XNORB3_15342_out0 && v$G27_5008_out0;
assign v$G24_16299_out0 = v$A3XNORB3_15343_out0 && v$G27_5009_out0;
assign v$A1XNORB1_16659_out0 = v$G16_17473_out0;
assign v$A1XNORB1_16662_out0 = v$G16_17476_out0;
assign v$A1XNORB1_16671_out0 = v$G16_17485_out0;
assign v$A1XNORB1_16674_out0 = v$G16_17488_out0;
assign v$B2_17245_out0 = v$SEL8_13485_out0;
assign v$B2_17246_out0 = v$SEL8_13486_out0;
assign v$B2_17248_out0 = v$SEL8_13488_out0;
assign v$B2_17249_out0 = v$SEL8_13489_out0;
assign v$B2_17257_out0 = v$SEL8_13497_out0;
assign v$B2_17258_out0 = v$SEL8_13498_out0;
assign v$B2_17260_out0 = v$SEL8_13500_out0;
assign v$B2_17261_out0 = v$SEL8_13501_out0;
assign v$S_17545_out0 = v$G9_9018_out0;
assign v$S_17556_out0 = v$G9_9019_out0;
assign v$G6_18041_out0 = v$G3_5216_out0 && v$G4_6660_out0;
assign v$MUX3_18332_out0 = v$G17_9229_out0 ? v$FF4_2541_out0 : v$_14689_out0;
assign v$MUX3_18333_out0 = v$G17_9230_out0 ? v$FF4_2542_out0 : v$_14690_out0;
assign v$B3_18461_out0 = v$SEL7_4325_out0;
assign v$B3_18462_out0 = v$SEL7_4326_out0;
assign v$B3_18464_out0 = v$SEL7_4328_out0;
assign v$B3_18465_out0 = v$SEL7_4329_out0;
assign v$B3_18473_out0 = v$SEL7_4337_out0;
assign v$B3_18474_out0 = v$SEL7_4338_out0;
assign v$B3_18476_out0 = v$SEL7_4340_out0;
assign v$B3_18477_out0 = v$SEL7_4341_out0;
assign v$MUX5_19171_out0 = v$G17_9229_out0 ? v$FF6_15909_out0 : v$_8404_out0;
assign v$MUX5_19172_out0 = v$G17_9230_out0 ? v$FF6_15910_out0 : v$_8405_out0;
assign v$G5_1269_out0 = v$FF2_13623_out0 && v$G6_16159_out0;
assign v$G5_1270_out0 = v$FF2_13624_out0 && v$G6_16160_out0;
assign v$G5_1271_out0 = v$FF2_13625_out0 && v$G6_16161_out0;
assign v$G5_1274_out0 = v$FF2_13634_out0 && v$G6_16170_out0;
assign v$G5_1275_out0 = v$FF2_13635_out0 && v$G6_16171_out0;
assign v$G5_1276_out0 = v$FF2_13636_out0 && v$G6_16172_out0;
assign v$G30_1936_out0 = v$A3$COMP$B3_5166_out0 || v$G31_16103_out0;
assign v$G30_1948_out0 = v$A3$COMP$B3_5178_out0 || v$G31_16115_out0;
assign v$G21_3723_out0 = ! v$B1_14823_out0;
assign v$G21_3724_out0 = ! v$B1_14824_out0;
assign v$G21_3726_out0 = ! v$B1_14826_out0;
assign v$G21_3727_out0 = ! v$B1_14827_out0;
assign v$G21_3735_out0 = ! v$B1_14835_out0;
assign v$G21_3736_out0 = ! v$B1_14836_out0;
assign v$G21_3738_out0 = ! v$B1_14838_out0;
assign v$G21_3739_out0 = ! v$B1_14839_out0;
assign v$G8_3908_out0 = !((v$A3_11201_out0 && !v$B3_18461_out0) || (!v$A3_11201_out0) && v$B3_18461_out0);
assign v$G8_3909_out0 = !((v$A3_11202_out0 && !v$B3_18462_out0) || (!v$A3_11202_out0) && v$B3_18462_out0);
assign v$G8_3911_out0 = !((v$A3_11204_out0 && !v$B3_18464_out0) || (!v$A3_11204_out0) && v$B3_18464_out0);
assign v$G8_3912_out0 = !((v$A3_11205_out0 && !v$B3_18465_out0) || (!v$A3_11205_out0) && v$B3_18465_out0);
assign v$G8_3920_out0 = !((v$A3_11213_out0 && !v$B3_18473_out0) || (!v$A3_11213_out0) && v$B3_18473_out0);
assign v$G8_3921_out0 = !((v$A3_11214_out0 && !v$B3_18474_out0) || (!v$A3_11214_out0) && v$B3_18474_out0);
assign v$G8_3923_out0 = !((v$A3_11216_out0 && !v$B3_18476_out0) || (!v$A3_11216_out0) && v$B3_18476_out0);
assign v$G8_3924_out0 = !((v$A3_11217_out0 && !v$B3_18477_out0) || (!v$A3_11217_out0) && v$B3_18477_out0);
assign v$OUT_4090_out0 = v$G30_1940_out0;
assign v$OUT_4091_out0 = v$G30_1941_out0;
assign v$OUT_4106_out0 = v$G30_1952_out0;
assign v$OUT_4107_out0 = v$G30_1953_out0;
assign v$G13_4564_out0 = v$A3XNORB3_15323_out0 && v$G11_16230_out0;
assign v$G13_4567_out0 = v$A3XNORB3_15326_out0 && v$G11_16233_out0;
assign v$G13_4576_out0 = v$A3XNORB3_15335_out0 && v$G11_16242_out0;
assign v$G13_4579_out0 = v$A3XNORB3_15338_out0 && v$G11_16245_out0;
assign v$A3$COMP$B3_5160_out0 = v$G5_7215_out0;
assign v$A3$COMP$B3_5163_out0 = v$G5_7218_out0;
assign v$A3$COMP$B3_5172_out0 = v$G5_7227_out0;
assign v$A3$COMP$B3_5175_out0 = v$G5_7230_out0;
assign v$G36_6185_out0 = !((v$B3_18461_out0 && !v$A3_11201_out0) || (!v$B3_18461_out0) && v$A3_11201_out0);
assign v$G36_6186_out0 = !((v$B3_18462_out0 && !v$A3_11202_out0) || (!v$B3_18462_out0) && v$A3_11202_out0);
assign v$G36_6188_out0 = !((v$B3_18464_out0 && !v$A3_11204_out0) || (!v$B3_18464_out0) && v$A3_11204_out0);
assign v$G36_6189_out0 = !((v$B3_18465_out0 && !v$A3_11205_out0) || (!v$B3_18465_out0) && v$A3_11205_out0);
assign v$G36_6197_out0 = !((v$B3_18473_out0 && !v$A3_11213_out0) || (!v$B3_18473_out0) && v$A3_11213_out0);
assign v$G36_6198_out0 = !((v$B3_18474_out0 && !v$A3_11214_out0) || (!v$B3_18474_out0) && v$A3_11214_out0);
assign v$G36_6200_out0 = !((v$B3_18476_out0 && !v$A3_11216_out0) || (!v$B3_18476_out0) && v$A3_11216_out0);
assign v$G36_6201_out0 = !((v$B3_18477_out0 && !v$A3_11217_out0) || (!v$B3_18477_out0) && v$A3_11217_out0);
assign v$G6_6784_out0 = ! v$B3_18461_out0;
assign v$G6_6785_out0 = ! v$B3_18462_out0;
assign v$G6_6787_out0 = ! v$B3_18464_out0;
assign v$G6_6788_out0 = ! v$B3_18465_out0;
assign v$G6_6796_out0 = ! v$B3_18473_out0;
assign v$G6_6797_out0 = ! v$B3_18474_out0;
assign v$G6_6799_out0 = ! v$B3_18476_out0;
assign v$G6_6800_out0 = ! v$B3_18477_out0;
assign v$_7872_out0 = { v$_10333_out0,v$_10333_out0 };
assign v$_7873_out0 = { v$_10334_out0,v$_10334_out0 };
assign v$A0$COMP$B0_8310_out0 = v$G24_16286_out0;
assign v$A0$COMP$B0_8311_out0 = v$G24_16287_out0;
assign v$A0$COMP$B0_8322_out0 = v$G24_16298_out0;
assign v$A0$COMP$B0_8323_out0 = v$G24_16299_out0;
assign v$G17_8488_out0 = !((v$A0_1886_out0 && !v$B0_3837_out0) || (!v$A0_1886_out0) && v$B0_3837_out0);
assign v$G17_8489_out0 = !((v$A0_1887_out0 && !v$B0_3838_out0) || (!v$A0_1887_out0) && v$B0_3838_out0);
assign v$G17_8491_out0 = !((v$A0_1889_out0 && !v$B0_3840_out0) || (!v$A0_1889_out0) && v$B0_3840_out0);
assign v$G17_8492_out0 = !((v$A0_1890_out0 && !v$B0_3841_out0) || (!v$A0_1890_out0) && v$B0_3841_out0);
assign v$G17_8500_out0 = !((v$A0_1898_out0 && !v$B0_3849_out0) || (!v$A0_1898_out0) && v$B0_3849_out0);
assign v$G17_8501_out0 = !((v$A0_1899_out0 && !v$B0_3850_out0) || (!v$A0_1899_out0) && v$B0_3850_out0);
assign v$G17_8503_out0 = !((v$A0_1901_out0 && !v$B0_3852_out0) || (!v$A0_1901_out0) && v$B0_3852_out0);
assign v$G17_8504_out0 = !((v$A0_1902_out0 && !v$B0_3853_out0) || (!v$A0_1902_out0) && v$B0_3853_out0);
assign v$G1_9761_out0 = v$LOWER$SAME_10635_out0 && v$HIGHER$SAME_15640_out0;
assign v$G1_9765_out0 = v$LOWER$SAME_10639_out0 && v$HIGHER$SAME_15644_out0;
assign v$G29_10754_out0 = v$A4$COMP$B4_7726_out0 || v$G30_1939_out0;
assign v$G29_10756_out0 = v$A4$COMP$B4_7728_out0 || v$G30_1951_out0;
assign v$G41_11374_out0 = v$G38_7609_out0 && v$G40_13945_out0;
assign v$G41_11377_out0 = v$G38_7612_out0 && v$G40_13948_out0;
assign v$G41_11386_out0 = v$G38_7621_out0 && v$G40_13957_out0;
assign v$G41_11389_out0 = v$G38_7624_out0 && v$G40_13960_out0;
assign v$G4_12406_out0 = v$G5_1268_out0 || v$S_17544_out0;
assign v$G4_12411_out0 = v$G5_1273_out0 || v$S_17555_out0;
assign v$G23_12741_out0 = ! v$B0_3837_out0;
assign v$G23_12742_out0 = ! v$B0_3838_out0;
assign v$G23_12744_out0 = ! v$B0_3840_out0;
assign v$G23_12745_out0 = ! v$B0_3841_out0;
assign v$G23_12753_out0 = ! v$B0_3849_out0;
assign v$G23_12754_out0 = ! v$B0_3850_out0;
assign v$G23_12756_out0 = ! v$B0_3852_out0;
assign v$G23_12757_out0 = ! v$B0_3853_out0;
assign v$G28_13591_out0 = v$A1XNORB1_16659_out0 && v$G25_11439_out0;
assign v$G28_13594_out0 = v$A1XNORB1_16662_out0 && v$G25_11442_out0;
assign v$G28_13603_out0 = v$A1XNORB1_16671_out0 && v$G25_11451_out0;
assign v$G28_13606_out0 = v$A1XNORB1_16674_out0 && v$G25_11454_out0;
assign v$G33_13676_out0 = !((v$A0_1886_out0 && !v$B0_3837_out0) || (!v$A0_1886_out0) && v$B0_3837_out0);
assign v$G33_13677_out0 = !((v$A0_1887_out0 && !v$B0_3838_out0) || (!v$A0_1887_out0) && v$B0_3838_out0);
assign v$G33_13679_out0 = !((v$A0_1889_out0 && !v$B0_3840_out0) || (!v$A0_1889_out0) && v$B0_3840_out0);
assign v$G33_13680_out0 = !((v$A0_1890_out0 && !v$B0_3841_out0) || (!v$A0_1890_out0) && v$B0_3841_out0);
assign v$G33_13688_out0 = !((v$A0_1898_out0 && !v$B0_3849_out0) || (!v$A0_1898_out0) && v$B0_3849_out0);
assign v$G33_13689_out0 = !((v$A0_1899_out0 && !v$B0_3850_out0) || (!v$A0_1899_out0) && v$B0_3850_out0);
assign v$G33_13691_out0 = !((v$A0_1901_out0 && !v$B0_3852_out0) || (!v$A0_1901_out0) && v$B0_3852_out0);
assign v$G33_13692_out0 = !((v$A0_1902_out0 && !v$B0_3853_out0) || (!v$A0_1902_out0) && v$B0_3853_out0);
assign v$G22_13912_out0 = v$A2XNORB2_4659_out0 && v$G20_10303_out0;
assign v$G22_13915_out0 = v$A2XNORB2_4662_out0 && v$G20_10306_out0;
assign v$G22_13924_out0 = v$A2XNORB2_4671_out0 && v$G20_10315_out0;
assign v$G22_13927_out0 = v$A2XNORB2_4674_out0 && v$G20_10318_out0;
assign v$NEXTSTATE_14112_out0 = v$G2_7901_out0;
assign v$NEXTSTATE_14115_out0 = v$G2_7904_out0;
assign v$G15_14223_out0 = !((v$A2_8372_out0 && !v$B2_17245_out0) || (!v$A2_8372_out0) && v$B2_17245_out0);
assign v$G15_14224_out0 = !((v$A2_8373_out0 && !v$B2_17246_out0) || (!v$A2_8373_out0) && v$B2_17246_out0);
assign v$G15_14226_out0 = !((v$A2_8375_out0 && !v$B2_17248_out0) || (!v$A2_8375_out0) && v$B2_17248_out0);
assign v$G15_14227_out0 = !((v$A2_8376_out0 && !v$B2_17249_out0) || (!v$A2_8376_out0) && v$B2_17249_out0);
assign v$G15_14235_out0 = !((v$A2_8384_out0 && !v$B2_17257_out0) || (!v$A2_8384_out0) && v$B2_17257_out0);
assign v$G15_14236_out0 = !((v$A2_8385_out0 && !v$B2_17258_out0) || (!v$A2_8385_out0) && v$B2_17258_out0);
assign v$G15_14238_out0 = !((v$A2_8387_out0 && !v$B2_17260_out0) || (!v$A2_8387_out0) && v$B2_17260_out0);
assign v$G15_14239_out0 = !((v$A2_8388_out0 && !v$B2_17261_out0) || (!v$A2_8388_out0) && v$B2_17261_out0);
assign v$Q_14759_out0 = v$G4_12405_out0;
assign v$Q_14770_out0 = v$G4_12410_out0;
assign v$G35_15123_out0 = !((v$A2_8372_out0 && !v$B2_17245_out0) || (!v$A2_8372_out0) && v$B2_17245_out0);
assign v$G35_15124_out0 = !((v$A2_8373_out0 && !v$B2_17246_out0) || (!v$A2_8373_out0) && v$B2_17246_out0);
assign v$G35_15126_out0 = !((v$A2_8375_out0 && !v$B2_17248_out0) || (!v$A2_8375_out0) && v$B2_17248_out0);
assign v$G35_15127_out0 = !((v$A2_8376_out0 && !v$B2_17249_out0) || (!v$A2_8376_out0) && v$B2_17249_out0);
assign v$G35_15135_out0 = !((v$A2_8384_out0 && !v$B2_17257_out0) || (!v$A2_8384_out0) && v$B2_17257_out0);
assign v$G35_15136_out0 = !((v$A2_8385_out0 && !v$B2_17258_out0) || (!v$A2_8385_out0) && v$B2_17258_out0);
assign v$G35_15138_out0 = !((v$A2_8387_out0 && !v$B2_17260_out0) || (!v$A2_8387_out0) && v$B2_17260_out0);
assign v$G35_15139_out0 = !((v$A2_8388_out0 && !v$B2_17261_out0) || (!v$A2_8388_out0) && v$B2_17261_out0);
assign v$G7_15414_out0 = v$G5_6084_out0 && v$G6_18041_out0;
assign v$MUX4_16602_out0 = v$EN_17563_out0 ? v$_1631_out0 : v$IN_9948_out0;
assign v$MUX4_16606_out0 = v$EN_17567_out0 ? v$_1635_out0 : v$IN_9952_out0;
assign v$G12_17095_out0 = ! v$B2_17245_out0;
assign v$G12_17096_out0 = ! v$B2_17246_out0;
assign v$G12_17098_out0 = ! v$B2_17248_out0;
assign v$G12_17099_out0 = ! v$B2_17249_out0;
assign v$G12_17107_out0 = ! v$B2_17257_out0;
assign v$G12_17108_out0 = ! v$B2_17258_out0;
assign v$G12_17110_out0 = ! v$B2_17260_out0;
assign v$G12_17111_out0 = ! v$B2_17261_out0;
assign v$EXP$SAME_17166_out0 = v$MUX4_12210_out0;
assign v$EXP$SAME_17167_out0 = v$MUX4_12211_out0;
assign v$G16_17474_out0 = !((v$A1_14944_out0 && !v$B1_14823_out0) || (!v$A1_14944_out0) && v$B1_14823_out0);
assign v$G16_17475_out0 = !((v$A1_14945_out0 && !v$B1_14824_out0) || (!v$A1_14945_out0) && v$B1_14824_out0);
assign v$G16_17477_out0 = !((v$A1_14947_out0 && !v$B1_14826_out0) || (!v$A1_14947_out0) && v$B1_14826_out0);
assign v$G16_17478_out0 = !((v$A1_14948_out0 && !v$B1_14827_out0) || (!v$A1_14948_out0) && v$B1_14827_out0);
assign v$G16_17486_out0 = !((v$A1_14956_out0 && !v$B1_14835_out0) || (!v$A1_14956_out0) && v$B1_14835_out0);
assign v$G16_17487_out0 = !((v$A1_14957_out0 && !v$B1_14836_out0) || (!v$A1_14957_out0) && v$B1_14836_out0);
assign v$G16_17489_out0 = !((v$A1_14959_out0 && !v$B1_14838_out0) || (!v$A1_14959_out0) && v$B1_14838_out0);
assign v$G16_17490_out0 = !((v$A1_14960_out0 && !v$B1_14839_out0) || (!v$A1_14960_out0) && v$B1_14839_out0);
assign v$G34_17932_out0 = !((v$A1_14944_out0 && !v$B1_14823_out0) || (!v$A1_14944_out0) && v$B1_14823_out0);
assign v$G34_17933_out0 = !((v$A1_14945_out0 && !v$B1_14824_out0) || (!v$A1_14945_out0) && v$B1_14824_out0);
assign v$G34_17935_out0 = !((v$A1_14947_out0 && !v$B1_14826_out0) || (!v$A1_14947_out0) && v$B1_14826_out0);
assign v$G34_17936_out0 = !((v$A1_14948_out0 && !v$B1_14827_out0) || (!v$A1_14948_out0) && v$B1_14827_out0);
assign v$G34_17944_out0 = !((v$A1_14956_out0 && !v$B1_14835_out0) || (!v$A1_14956_out0) && v$B1_14835_out0);
assign v$G34_17945_out0 = !((v$A1_14957_out0 && !v$B1_14836_out0) || (!v$A1_14957_out0) && v$B1_14836_out0);
assign v$G34_17947_out0 = !((v$A1_14959_out0 && !v$B1_14838_out0) || (!v$A1_14959_out0) && v$B1_14838_out0);
assign v$G34_17948_out0 = !((v$A1_14960_out0 && !v$B1_14839_out0) || (!v$A1_14960_out0) && v$B1_14839_out0);
assign v$G32_418_out0 = v$A1$COMP$B1_13087_out0 || v$A0$COMP$B0_8310_out0;
assign v$G32_419_out0 = v$A1$COMP$B1_13088_out0 || v$A0$COMP$B0_8311_out0;
assign v$G32_430_out0 = v$A1$COMP$B1_13099_out0 || v$A0$COMP$B0_8322_out0;
assign v$G32_431_out0 = v$A1$COMP$B1_13100_out0 || v$A0$COMP$B0_8323_out0;
assign v$A0XNORB0_1584_out0 = v$G17_8488_out0;
assign v$A0XNORB0_1585_out0 = v$G17_8489_out0;
assign v$A0XNORB0_1587_out0 = v$G17_8491_out0;
assign v$A0XNORB0_1588_out0 = v$G17_8492_out0;
assign v$A0XNORB0_1596_out0 = v$G17_8500_out0;
assign v$A0XNORB0_1597_out0 = v$G17_8501_out0;
assign v$A0XNORB0_1599_out0 = v$G17_8503_out0;
assign v$A0XNORB0_1600_out0 = v$G17_8504_out0;
assign v$A2$COMP$B2_2135_out0 = v$G13_4564_out0;
assign v$A2$COMP$B2_2138_out0 = v$G13_4567_out0;
assign v$A2$COMP$B2_2147_out0 = v$G13_4576_out0;
assign v$A2$COMP$B2_2150_out0 = v$G13_4579_out0;
assign v$MUX6_3072_out0 = v$FF1_14261_out0 ? v$LSBS_15901_out0 : v$_7872_out0;
assign v$MUX6_3073_out0 = v$FF1_14262_out0 ? v$LSBS_15902_out0 : v$_7873_out0;
assign v$HIGHER$OUT_4014_out0 = v$OUT_4090_out0;
assign v$HIGHER$OUT_4018_out0 = v$OUT_4106_out0;
assign v$OUT_4088_out0 = v$G29_10754_out0;
assign v$OUT_4104_out0 = v$G29_10756_out0;
assign v$LOWER$OUT_4383_out0 = v$OUT_4091_out0;
assign v$LOWER$OUT_4387_out0 = v$OUT_4107_out0;
assign v$A2XNORB2_4660_out0 = v$G15_14223_out0;
assign v$A2XNORB2_4661_out0 = v$G15_14224_out0;
assign v$A2XNORB2_4663_out0 = v$G15_14226_out0;
assign v$A2XNORB2_4664_out0 = v$G15_14227_out0;
assign v$A2XNORB2_4672_out0 = v$G15_14235_out0;
assign v$A2XNORB2_4673_out0 = v$G15_14236_out0;
assign v$A2XNORB2_4675_out0 = v$G15_14238_out0;
assign v$A2XNORB2_4676_out0 = v$G15_14239_out0;
assign v$G27_4989_out0 = v$A2XNORB2_4659_out0 && v$G28_13591_out0;
assign v$G27_4992_out0 = v$A2XNORB2_4662_out0 && v$G28_13594_out0;
assign v$G27_5001_out0 = v$A2XNORB2_4671_out0 && v$G28_13603_out0;
assign v$G27_5004_out0 = v$A2XNORB2_4674_out0 && v$G28_13606_out0;
assign v$G18_5188_out0 = v$A3XNORB3_15323_out0 && v$G22_13912_out0;
assign v$G18_5191_out0 = v$A3XNORB3_15326_out0 && v$G22_13915_out0;
assign v$G18_5200_out0 = v$A3XNORB3_15335_out0 && v$G22_13924_out0;
assign v$G18_5203_out0 = v$A3XNORB3_15338_out0 && v$G22_13927_out0;
assign v$G5_7216_out0 = v$A3_11201_out0 && v$G6_6784_out0;
assign v$G5_7217_out0 = v$A3_11202_out0 && v$G6_6785_out0;
assign v$G5_7219_out0 = v$A3_11204_out0 && v$G6_6787_out0;
assign v$G5_7220_out0 = v$A3_11205_out0 && v$G6_6788_out0;
assign v$G5_7228_out0 = v$A3_11213_out0 && v$G6_6796_out0;
assign v$G5_7229_out0 = v$A3_11214_out0 && v$G6_6797_out0;
assign v$G5_7231_out0 = v$A3_11216_out0 && v$G6_6799_out0;
assign v$G5_7232_out0 = v$A3_11217_out0 && v$G6_6800_out0;
assign v$G38_7610_out0 = v$G33_13676_out0 && v$G34_17932_out0;
assign v$G38_7611_out0 = v$G33_13677_out0 && v$G34_17933_out0;
assign v$G38_7613_out0 = v$G33_13679_out0 && v$G34_17935_out0;
assign v$G38_7614_out0 = v$G33_13680_out0 && v$G34_17936_out0;
assign v$G38_7622_out0 = v$G33_13688_out0 && v$G34_17944_out0;
assign v$G38_7623_out0 = v$G33_13689_out0 && v$G34_17945_out0;
assign v$G38_7625_out0 = v$G33_13691_out0 && v$G34_17947_out0;
assign v$G38_7626_out0 = v$G33_13692_out0 && v$G34_17948_out0;
assign v$TXFlag_8035_out0 = v$Q_14759_out0;
assign v$TXFlag_8036_out0 = v$Q_14770_out0;
assign v$IGNORE_8594_out0 = v$G7_15414_out0;
assign v$G20_10304_out0 = v$A1_14944_out0 && v$G21_3723_out0;
assign v$G20_10305_out0 = v$A1_14945_out0 && v$G21_3724_out0;
assign v$G20_10307_out0 = v$A1_14947_out0 && v$G21_3726_out0;
assign v$G20_10308_out0 = v$A1_14948_out0 && v$G21_3727_out0;
assign v$G20_10316_out0 = v$A1_14956_out0 && v$G21_3735_out0;
assign v$G20_10317_out0 = v$A1_14957_out0 && v$G21_3736_out0;
assign v$G20_10319_out0 = v$A1_14959_out0 && v$G21_3738_out0;
assign v$G20_10320_out0 = v$A1_14960_out0 && v$G21_3739_out0;
assign v$G29_10753_out0 = v$A4$COMP$B4_7725_out0 || v$G30_1936_out0;
assign v$G29_10755_out0 = v$A4$COMP$B4_7727_out0 || v$G30_1948_out0;
assign v$G25_11440_out0 = v$A0_1886_out0 && v$G23_12741_out0;
assign v$G25_11441_out0 = v$A0_1887_out0 && v$G23_12742_out0;
assign v$G25_11443_out0 = v$A0_1889_out0 && v$G23_12744_out0;
assign v$G25_11444_out0 = v$A0_1890_out0 && v$G23_12745_out0;
assign v$G25_11452_out0 = v$A0_1898_out0 && v$G23_12753_out0;
assign v$G25_11453_out0 = v$A0_1899_out0 && v$G23_12754_out0;
assign v$G25_11455_out0 = v$A0_1901_out0 && v$G23_12756_out0;
assign v$G25_11456_out0 = v$A0_1902_out0 && v$G23_12757_out0;
assign v$G4_12407_out0 = v$G5_1269_out0 || v$S_17545_out0;
assign v$G4_12408_out0 = v$G5_1270_out0 || v$S_17546_out0;
assign v$G4_12409_out0 = v$G5_1271_out0 || v$S_17547_out0;
assign v$G4_12412_out0 = v$G5_1274_out0 || v$S_17556_out0;
assign v$G4_12413_out0 = v$G5_1275_out0 || v$S_17557_out0;
assign v$G4_12414_out0 = v$G5_1276_out0 || v$S_17558_out0;
assign v$MUX2_12605_out0 = v$G3_2802_out0 ? v$_9821_out0 : v$MUX4_16602_out0;
assign v$MUX2_12609_out0 = v$G3_2806_out0 ? v$_9825_out0 : v$MUX4_16606_out0;
assign v$G40_13946_out0 = v$G35_15123_out0 && v$G36_6185_out0;
assign v$G40_13947_out0 = v$G35_15124_out0 && v$G36_6186_out0;
assign v$G40_13949_out0 = v$G35_15126_out0 && v$G36_6188_out0;
assign v$G40_13950_out0 = v$G35_15127_out0 && v$G36_6189_out0;
assign v$G40_13958_out0 = v$G35_15135_out0 && v$G36_6197_out0;
assign v$G40_13959_out0 = v$G35_15136_out0 && v$G36_6198_out0;
assign v$G40_13961_out0 = v$G35_15138_out0 && v$G36_6200_out0;
assign v$G40_13962_out0 = v$G35_15139_out0 && v$G36_6201_out0;
assign v$Q_14760_out0 = v$G4_12406_out0;
assign v$Q_14771_out0 = v$G4_12411_out0;
assign v$A3XNORB3_15324_out0 = v$G8_3908_out0;
assign v$A3XNORB3_15325_out0 = v$G8_3909_out0;
assign v$A3XNORB3_15327_out0 = v$G8_3911_out0;
assign v$A3XNORB3_15328_out0 = v$G8_3912_out0;
assign v$A3XNORB3_15336_out0 = v$G8_3920_out0;
assign v$A3XNORB3_15337_out0 = v$G8_3921_out0;
assign v$A3XNORB3_15339_out0 = v$G8_3923_out0;
assign v$A3XNORB3_15340_out0 = v$G8_3924_out0;
assign v$G11_16231_out0 = v$A2_8372_out0 && v$G12_17095_out0;
assign v$G11_16232_out0 = v$A2_8373_out0 && v$G12_17096_out0;
assign v$G11_16234_out0 = v$A2_8375_out0 && v$G12_17098_out0;
assign v$G11_16235_out0 = v$A2_8376_out0 && v$G12_17099_out0;
assign v$G11_16243_out0 = v$A2_8384_out0 && v$G12_17107_out0;
assign v$G11_16244_out0 = v$A2_8385_out0 && v$G12_17108_out0;
assign v$G11_16246_out0 = v$A2_8387_out0 && v$G12_17110_out0;
assign v$G11_16247_out0 = v$A2_8388_out0 && v$G12_17111_out0;
assign v$A1XNORB1_16660_out0 = v$G16_17474_out0;
assign v$A1XNORB1_16661_out0 = v$G16_17475_out0;
assign v$A1XNORB1_16663_out0 = v$G16_17477_out0;
assign v$A1XNORB1_16664_out0 = v$G16_17478_out0;
assign v$A1XNORB1_16672_out0 = v$G16_17486_out0;
assign v$A1XNORB1_16673_out0 = v$G16_17487_out0;
assign v$A1XNORB1_16675_out0 = v$G16_17489_out0;
assign v$A1XNORB1_16676_out0 = v$G16_17490_out0;
assign v$SAME_19333_out0 = v$G41_11374_out0;
assign v$SAME_19337_out0 = v$G41_11377_out0;
assign v$SAME_19342_out0 = v$G1_9761_out0;
assign v$SAME_19349_out0 = v$G41_11386_out0;
assign v$SAME_19353_out0 = v$G41_11389_out0;
assign v$SAME_19358_out0 = v$G1_9765_out0;
assign v$MUX3_3601_out0 = v$OUT_4088_out0 ? v$A$EXP_298_out0 : v$B$EXP_17296_out0;
assign v$MUX3_3605_out0 = v$OUT_4104_out0 ? v$A$EXP_302_out0 : v$B$EXP_17300_out0;
assign v$OUT_4084_out0 = v$G29_10753_out0;
assign v$OUT_4100_out0 = v$G29_10755_out0;
assign v$G13_4565_out0 = v$A3XNORB3_15324_out0 && v$G11_16231_out0;
assign v$G13_4566_out0 = v$A3XNORB3_15325_out0 && v$G11_16232_out0;
assign v$G13_4568_out0 = v$A3XNORB3_15327_out0 && v$G11_16234_out0;
assign v$G13_4569_out0 = v$A3XNORB3_15328_out0 && v$G11_16235_out0;
assign v$G13_4577_out0 = v$A3XNORB3_15336_out0 && v$G11_16243_out0;
assign v$G13_4578_out0 = v$A3XNORB3_15337_out0 && v$G11_16244_out0;
assign v$G13_4580_out0 = v$A3XNORB3_15339_out0 && v$G11_16246_out0;
assign v$G13_4581_out0 = v$A3XNORB3_15340_out0 && v$G11_16247_out0;
assign v$A3$COMP$B3_5161_out0 = v$G5_7216_out0;
assign v$A3$COMP$B3_5162_out0 = v$G5_7217_out0;
assign v$A3$COMP$B3_5164_out0 = v$G5_7219_out0;
assign v$A3$COMP$B3_5165_out0 = v$G5_7220_out0;
assign v$A3$COMP$B3_5173_out0 = v$G5_7228_out0;
assign v$A3$COMP$B3_5174_out0 = v$G5_7229_out0;
assign v$A3$COMP$B3_5176_out0 = v$G5_7231_out0;
assign v$A3$COMP$B3_5177_out0 = v$G5_7232_out0;
assign v$G3_9162_out0 = v$HIGHER$SAME_15641_out0 && v$LOWER$OUT_4383_out0;
assign v$G3_9166_out0 = v$HIGHER$SAME_15645_out0 && v$LOWER$OUT_4387_out0;
assign v$HIGHER$SAME_9460_out0 = v$SAME_19333_out0;
assign v$HIGHER$SAME_9461_out0 = v$SAME_19337_out0;
assign v$HIGHER$SAME_9462_out0 = v$SAME_19349_out0;
assign v$HIGHER$SAME_9463_out0 = v$SAME_19353_out0;
assign v$G41_11375_out0 = v$G38_7610_out0 && v$G40_13946_out0;
assign v$G41_11376_out0 = v$G38_7611_out0 && v$G40_13947_out0;
assign v$G41_11378_out0 = v$G38_7613_out0 && v$G40_13949_out0;
assign v$G41_11379_out0 = v$G38_7614_out0 && v$G40_13950_out0;
assign v$G41_11387_out0 = v$G38_7622_out0 && v$G40_13958_out0;
assign v$G41_11388_out0 = v$G38_7623_out0 && v$G40_13959_out0;
assign v$G41_11390_out0 = v$G38_7625_out0 && v$G40_13961_out0;
assign v$G41_11391_out0 = v$G38_7626_out0 && v$G40_13962_out0;
assign v$_12382_out0 = { v$_15239_out0,v$MUX6_3072_out0 };
assign v$_12386_out0 = { v$_15243_out0,v$MUX6_3073_out0 };
assign v$A1$COMP$B1_13080_out0 = v$G18_5188_out0;
assign v$A1$COMP$B1_13083_out0 = v$G18_5191_out0;
assign v$A1$COMP$B1_13092_out0 = v$G18_5200_out0;
assign v$A1$COMP$B1_13095_out0 = v$G18_5203_out0;
assign v$G28_13592_out0 = v$A1XNORB1_16660_out0 && v$G25_11440_out0;
assign v$G28_13593_out0 = v$A1XNORB1_16661_out0 && v$G25_11441_out0;
assign v$G28_13595_out0 = v$A1XNORB1_16663_out0 && v$G25_11443_out0;
assign v$G28_13596_out0 = v$A1XNORB1_16664_out0 && v$G25_11444_out0;
assign v$G28_13604_out0 = v$A1XNORB1_16672_out0 && v$G25_11452_out0;
assign v$G28_13605_out0 = v$A1XNORB1_16673_out0 && v$G25_11453_out0;
assign v$G28_13607_out0 = v$A1XNORB1_16675_out0 && v$G25_11455_out0;
assign v$G28_13608_out0 = v$A1XNORB1_16676_out0 && v$G25_11456_out0;
assign v$G22_13913_out0 = v$A2XNORB2_4660_out0 && v$G20_10304_out0;
assign v$G22_13914_out0 = v$A2XNORB2_4661_out0 && v$G20_10305_out0;
assign v$G22_13916_out0 = v$A2XNORB2_4663_out0 && v$G20_10307_out0;
assign v$G22_13917_out0 = v$A2XNORB2_4664_out0 && v$G20_10308_out0;
assign v$G22_13925_out0 = v$A2XNORB2_4672_out0 && v$G20_10316_out0;
assign v$G22_13926_out0 = v$A2XNORB2_4673_out0 && v$G20_10317_out0;
assign v$G22_13928_out0 = v$A2XNORB2_4675_out0 && v$G20_10319_out0;
assign v$G22_13929_out0 = v$A2XNORB2_4676_out0 && v$G20_10320_out0;
assign v$OUT_14343_out0 = v$OUT_4088_out0;
assign v$OUT_14347_out0 = v$OUT_4104_out0;
assign v$Q_14761_out0 = v$G4_12407_out0;
assign v$Q_14762_out0 = v$G4_12408_out0;
assign v$Q_14763_out0 = v$G4_12409_out0;
assign v$Q_14772_out0 = v$G4_12412_out0;
assign v$Q_14773_out0 = v$G4_12413_out0;
assign v$Q_14774_out0 = v$G4_12414_out0;
assign v$TXFlag_15829_out0 = v$TXFlag_8035_out0;
assign v$TXFlag_15830_out0 = v$TXFlag_8036_out0;
assign v$G31_16104_out0 = v$A2$COMP$B2_2142_out0 || v$G32_418_out0;
assign v$G31_16105_out0 = v$A2$COMP$B2_2143_out0 || v$G32_419_out0;
assign v$G31_16116_out0 = v$A2$COMP$B2_2154_out0 || v$G32_430_out0;
assign v$G31_16117_out0 = v$A2$COMP$B2_2155_out0 || v$G32_431_out0;
assign v$G24_16279_out0 = v$A3XNORB3_15323_out0 && v$G27_4989_out0;
assign v$G24_16282_out0 = v$A3XNORB3_15326_out0 && v$G27_4992_out0;
assign v$G24_16291_out0 = v$A3XNORB3_15335_out0 && v$G27_5001_out0;
assign v$G24_16294_out0 = v$A3XNORB3_15338_out0 && v$G27_5004_out0;
assign v$RXflag_16445_out0 = v$Q_14760_out0;
assign v$RXflag_16446_out0 = v$Q_14771_out0;
assign v$G6_17432_out0 = ! v$IGNORE_8594_out0;
assign v$MUX1_18539_out0 = v$OUT_4088_out0 ? v$B$EXP_17296_out0 : v$A$EXP_298_out0;
assign v$MUX1_18543_out0 = v$OUT_4104_out0 ? v$B$EXP_17300_out0 : v$A$EXP_302_out0;
assign v$SAME_18969_out0 = v$SAME_19342_out0;
assign v$SAME_18973_out0 = v$SAME_19358_out0;
assign v$G30_1937_out0 = v$A3$COMP$B3_5167_out0 || v$G31_16104_out0;
assign v$G30_1938_out0 = v$A3$COMP$B3_5168_out0 || v$G31_16105_out0;
assign v$G30_1949_out0 = v$A3$COMP$B3_5179_out0 || v$G31_16116_out0;
assign v$G30_1950_out0 = v$A3$COMP$B3_5180_out0 || v$G31_16117_out0;
assign v$A2$COMP$B2_2136_out0 = v$G13_4565_out0;
assign v$A2$COMP$B2_2137_out0 = v$G13_4566_out0;
assign v$A2$COMP$B2_2139_out0 = v$G13_4568_out0;
assign v$A2$COMP$B2_2140_out0 = v$G13_4569_out0;
assign v$A2$COMP$B2_2148_out0 = v$G13_4577_out0;
assign v$A2$COMP$B2_2149_out0 = v$G13_4578_out0;
assign v$A2$COMP$B2_2151_out0 = v$G13_4580_out0;
assign v$A2$COMP$B2_2152_out0 = v$G13_4581_out0;
assign v$MUX14_3166_out0 = v$IS$32$BIT_11362_out0 ? v$SAME_18969_out0 : v$SAME_18968_out0;
assign v$MUX14_3167_out0 = v$IS$32$BIT_11363_out0 ? v$SAME_18973_out0 : v$SAME_18972_out0;
assign v$MUX3_3599_out0 = v$OUT_4084_out0 ? v$A$EXP_296_out0 : v$B$EXP_17294_out0;
assign v$MUX3_3603_out0 = v$OUT_4100_out0 ? v$A$EXP_300_out0 : v$B$EXP_17298_out0;
assign v$Error_3949_out0 = v$Q_14763_out0;
assign v$Error_3950_out0 = v$Q_14774_out0;
assign v$TXoverflow_4265_out0 = v$Q_14761_out0;
assign v$TXoverflow_4266_out0 = v$Q_14772_out0;
assign v$G27_4990_out0 = v$A2XNORB2_4660_out0 && v$G28_13592_out0;
assign v$G27_4991_out0 = v$A2XNORB2_4661_out0 && v$G28_13593_out0;
assign v$G27_4993_out0 = v$A2XNORB2_4663_out0 && v$G28_13595_out0;
assign v$G27_4994_out0 = v$A2XNORB2_4664_out0 && v$G28_13596_out0;
assign v$G27_5002_out0 = v$A2XNORB2_4672_out0 && v$G28_13604_out0;
assign v$G27_5003_out0 = v$A2XNORB2_4673_out0 && v$G28_13605_out0;
assign v$G27_5005_out0 = v$A2XNORB2_4675_out0 && v$G28_13607_out0;
assign v$G27_5006_out0 = v$A2XNORB2_4676_out0 && v$G28_13608_out0;
assign v$G18_5189_out0 = v$A3XNORB3_15324_out0 && v$G22_13913_out0;
assign v$G18_5190_out0 = v$A3XNORB3_15325_out0 && v$G22_13914_out0;
assign v$G18_5192_out0 = v$A3XNORB3_15327_out0 && v$G22_13916_out0;
assign v$G18_5193_out0 = v$A3XNORB3_15328_out0 && v$G22_13917_out0;
assign v$G18_5201_out0 = v$A3XNORB3_15336_out0 && v$G22_13925_out0;
assign v$G18_5202_out0 = v$A3XNORB3_15337_out0 && v$G22_13926_out0;
assign v$G18_5204_out0 = v$A3XNORB3_15339_out0 && v$G22_13928_out0;
assign v$G18_5205_out0 = v$A3XNORB3_15340_out0 && v$G22_13929_out0;
assign v$MUX1_6916_out0 = v$G4_4188_out0 ? v$_12382_out0 : v$MUX2_12605_out0;
assign v$MUX1_6920_out0 = v$G4_4192_out0 ? v$_12386_out0 : v$MUX2_12609_out0;
assign v$XOR1_7918_out0 = v$C1_14150_out0 ^ v$MUX1_18539_out0;
assign v$XOR1_7922_out0 = v$C1_14154_out0 ^ v$MUX1_18543_out0;
assign v$A0$COMP$B0_8303_out0 = v$G24_16279_out0;
assign v$A0$COMP$B0_8306_out0 = v$G24_16282_out0;
assign v$A0$COMP$B0_8315_out0 = v$G24_16291_out0;
assign v$A0$COMP$B0_8318_out0 = v$G24_16294_out0;
assign v$RXoverflow_9918_out0 = v$Q_14762_out0;
assign v$RXoverflow_9919_out0 = v$Q_14773_out0;
assign v$RXFLAG_12700_out0 = v$RXflag_16445_out0;
assign v$RXFLAG_12701_out0 = v$RXflag_16446_out0;
assign v$G2_13478_out0 = v$HIGHER$OUT_4014_out0 || v$G3_9162_out0;
assign v$G2_13482_out0 = v$HIGHER$OUT_4018_out0 || v$G3_9166_out0;
assign v$OUT_14341_out0 = v$OUT_4084_out0;
assign v$OUT_14345_out0 = v$OUT_4100_out0;
assign v$TXFLAG_15295_out0 = v$TXFlag_15829_out0;
assign v$TXFLAG_15296_out0 = v$TXFlag_15830_out0;
assign v$G7_18265_out0 = v$G5_2865_out0 && v$G6_17432_out0;
assign v$MUX1_18537_out0 = v$OUT_4084_out0 ? v$B$EXP_17294_out0 : v$A$EXP_296_out0;
assign v$MUX1_18541_out0 = v$OUT_4100_out0 ? v$B$EXP_17298_out0 : v$A$EXP_300_out0;
assign v$SAME_19335_out0 = v$G41_11375_out0;
assign v$SAME_19336_out0 = v$G41_11376_out0;
assign v$SAME_19339_out0 = v$G41_11378_out0;
assign v$SAME_19340_out0 = v$G41_11379_out0;
assign v$SAME_19351_out0 = v$G41_11387_out0;
assign v$SAME_19352_out0 = v$G41_11388_out0;
assign v$SAME_19355_out0 = v$G41_11390_out0;
assign v$SAME_19356_out0 = v$G41_11391_out0;
assign v$G32_411_out0 = v$A1$COMP$B1_13080_out0 || v$A0$COMP$B0_8303_out0;
assign v$G32_414_out0 = v$A1$COMP$B1_13083_out0 || v$A0$COMP$B0_8306_out0;
assign v$G32_423_out0 = v$A1$COMP$B1_13092_out0 || v$A0$COMP$B0_8315_out0;
assign v$G32_426_out0 = v$A1$COMP$B1_13095_out0 || v$A0$COMP$B0_8318_out0;
assign v$EXP$SAME_1006_out0 = v$MUX14_3166_out0;
assign v$EXP$SAME_1007_out0 = v$MUX14_3167_out0;
assign v$MUX3_2124_out0 = v$G8_2052_out0 ? v$_13892_out0 : v$MUX1_6916_out0;
assign v$MUX3_2128_out0 = v$G8_2056_out0 ? v$_13896_out0 : v$MUX1_6920_out0;
assign v$TXFLAG_4060_out0 = v$TXFLAG_15295_out0;
assign v$TXFLAG_4061_out0 = v$TXFLAG_15296_out0;
assign v$OUT_4086_out0 = v$G30_1937_out0;
assign v$OUT_4087_out0 = v$G30_1938_out0;
assign v$OUT_4089_out0 = v$G2_13478_out0;
assign v$OUT_4102_out0 = v$G30_1949_out0;
assign v$OUT_4103_out0 = v$G30_1950_out0;
assign v$OUT_4105_out0 = v$G2_13482_out0;
assign {v$A1_6078_out1,v$A1_6078_out0 } = v$MUX3_3601_out0 + v$XOR1_7918_out0 + v$CIN_18828_out0;
assign {v$A1_6082_out1,v$A1_6082_out0 } = v$MUX3_3605_out0 + v$XOR1_7922_out0 + v$CIN_18832_out0;
assign v$XOR1_7916_out0 = v$C1_14148_out0 ^ v$MUX1_18537_out0;
assign v$XOR1_7920_out0 = v$C1_14152_out0 ^ v$MUX1_18541_out0;
assign v$_10339_out0 = { v$RXoverflow_9918_out0,v$Error_3949_out0 };
assign v$_10340_out0 = { v$RXoverflow_9919_out0,v$Error_3950_out0 };
assign v$LOWER$SAME_10633_out0 = v$SAME_19336_out0;
assign v$LOWER$SAME_10634_out0 = v$SAME_19340_out0;
assign v$LOWER$SAME_10637_out0 = v$SAME_19352_out0;
assign v$LOWER$SAME_10638_out0 = v$SAME_19356_out0;
assign v$A1$COMP$B1_13081_out0 = v$G18_5189_out0;
assign v$A1$COMP$B1_13082_out0 = v$G18_5190_out0;
assign v$A1$COMP$B1_13084_out0 = v$G18_5192_out0;
assign v$A1$COMP$B1_13085_out0 = v$G18_5193_out0;
assign v$A1$COMP$B1_13093_out0 = v$G18_5201_out0;
assign v$A1$COMP$B1_13094_out0 = v$G18_5202_out0;
assign v$A1$COMP$B1_13096_out0 = v$G18_5204_out0;
assign v$A1$COMP$B1_13097_out0 = v$G18_5205_out0;
assign v$RXFLAG_15620_out0 = v$RXFLAG_12700_out0;
assign v$RXFLAG_15621_out0 = v$RXFLAG_12701_out0;
assign v$HIGHER$SAME_15638_out0 = v$SAME_19335_out0;
assign v$HIGHER$SAME_15639_out0 = v$SAME_19339_out0;
assign v$HIGHER$SAME_15642_out0 = v$SAME_19351_out0;
assign v$HIGHER$SAME_15643_out0 = v$SAME_19355_out0;
assign v$_15881_out0 = { v$TXFlag_8035_out0,v$TXoverflow_4265_out0 };
assign v$_15882_out0 = { v$TXFlag_8036_out0,v$TXoverflow_4266_out0 };
assign v$G24_16280_out0 = v$A3XNORB3_15324_out0 && v$G27_4990_out0;
assign v$G24_16281_out0 = v$A3XNORB3_15325_out0 && v$G27_4991_out0;
assign v$G24_16283_out0 = v$A3XNORB3_15327_out0 && v$G27_4993_out0;
assign v$G24_16284_out0 = v$A3XNORB3_15328_out0 && v$G27_4994_out0;
assign v$G24_16292_out0 = v$A3XNORB3_15336_out0 && v$G27_5002_out0;
assign v$G24_16293_out0 = v$A3XNORB3_15337_out0 && v$G27_5003_out0;
assign v$G24_16295_out0 = v$A3XNORB3_15339_out0 && v$G27_5005_out0;
assign v$G24_16296_out0 = v$A3XNORB3_15340_out0 && v$G27_5006_out0;
assign v$RAMWEN_18576_out0 = v$G7_18265_out0;
assign v$F_2133_out0 = v$TXFLAG_4060_out0;
assign v$F_2134_out0 = v$TXFLAG_4061_out0;
assign v$OUT_3399_out0 = v$MUX3_2124_out0;
assign v$OUT_3403_out0 = v$MUX3_2128_out0;
assign v$MUX3_3602_out0 = v$OUT_4089_out0 ? v$A$EXP_299_out0 : v$B$EXP_17297_out0;
assign v$MUX3_3606_out0 = v$OUT_4105_out0 ? v$A$EXP_303_out0 : v$B$EXP_17301_out0;
assign v$HIGHER$OUT_4013_out0 = v$OUT_4086_out0;
assign v$HIGHER$OUT_4017_out0 = v$OUT_4102_out0;
assign v$LOWER$OUT_4382_out0 = v$OUT_4087_out0;
assign v$LOWER$OUT_4386_out0 = v$OUT_4103_out0;
assign {v$A1_6076_out1,v$A1_6076_out0 } = v$MUX3_3599_out0 + v$XOR1_7916_out0 + v$CIN_18826_out0;
assign {v$A1_6080_out1,v$A1_6080_out0 } = v$MUX3_3603_out0 + v$XOR1_7920_out0 + v$CIN_18830_out0;
assign v$A0$COMP$B0_8304_out0 = v$G24_16280_out0;
assign v$A0$COMP$B0_8305_out0 = v$G24_16281_out0;
assign v$A0$COMP$B0_8307_out0 = v$G24_16283_out0;
assign v$A0$COMP$B0_8308_out0 = v$G24_16284_out0;
assign v$A0$COMP$B0_8316_out0 = v$G24_16292_out0;
assign v$A0$COMP$B0_8317_out0 = v$G24_16293_out0;
assign v$A0$COMP$B0_8319_out0 = v$G24_16295_out0;
assign v$A0$COMP$B0_8320_out0 = v$G24_16296_out0;
assign v$DIFF_9416_out0 = v$A1_6078_out0;
assign v$DIFF_9420_out0 = v$A1_6082_out0;
assign v$G1_9759_out0 = v$LOWER$SAME_10633_out0 && v$HIGHER$SAME_15638_out0;
assign v$G1_9760_out0 = v$LOWER$SAME_10634_out0 && v$HIGHER$SAME_15639_out0;
assign v$G1_9763_out0 = v$LOWER$SAME_10637_out0 && v$HIGHER$SAME_15642_out0;
assign v$G1_9764_out0 = v$LOWER$SAME_10638_out0 && v$HIGHER$SAME_15643_out0;
assign v$OUT_14344_out0 = v$OUT_4089_out0;
assign v$OUT_14348_out0 = v$OUT_4105_out0;
assign v$NOT$USED1_14985_out0 = v$A1_6078_out1;
assign v$NOT$USED1_14989_out0 = v$A1_6082_out1;
assign v$G31_16097_out0 = v$A2$COMP$B2_2135_out0 || v$G32_411_out0;
assign v$G31_16100_out0 = v$A2$COMP$B2_2138_out0 || v$G32_414_out0;
assign v$G31_16109_out0 = v$A2$COMP$B2_2147_out0 || v$G32_423_out0;
assign v$G31_16112_out0 = v$A2$COMP$B2_2150_out0 || v$G32_426_out0;
assign v$MUX1_18540_out0 = v$OUT_4089_out0 ? v$B$EXP_17297_out0 : v$A$EXP_299_out0;
assign v$MUX1_18544_out0 = v$OUT_4105_out0 ? v$B$EXP_17301_out0 : v$A$EXP_303_out0;
assign v$_19155_out0 = { v$RXflag_16445_out0,v$_10339_out0 };
assign v$_19156_out0 = { v$RXflag_16446_out0,v$_10340_out0 };
assign v$G32_412_out0 = v$A1$COMP$B1_13081_out0 || v$A0$COMP$B0_8304_out0;
assign v$G32_413_out0 = v$A1$COMP$B1_13082_out0 || v$A0$COMP$B0_8305_out0;
assign v$G32_415_out0 = v$A1$COMP$B1_13084_out0 || v$A0$COMP$B0_8307_out0;
assign v$G32_416_out0 = v$A1$COMP$B1_13085_out0 || v$A0$COMP$B0_8308_out0;
assign v$G32_424_out0 = v$A1$COMP$B1_13093_out0 || v$A0$COMP$B0_8316_out0;
assign v$G32_425_out0 = v$A1$COMP$B1_13094_out0 || v$A0$COMP$B0_8317_out0;
assign v$G32_427_out0 = v$A1$COMP$B1_13096_out0 || v$A0$COMP$B0_8319_out0;
assign v$G32_428_out0 = v$A1$COMP$B1_13097_out0 || v$A0$COMP$B0_8320_out0;
assign v$G30_1930_out0 = v$A3$COMP$B3_5160_out0 || v$G31_16097_out0;
assign v$G30_1933_out0 = v$A3$COMP$B3_5163_out0 || v$G31_16100_out0;
assign v$G30_1942_out0 = v$A3$COMP$B3_5172_out0 || v$G31_16109_out0;
assign v$G30_1945_out0 = v$A3$COMP$B3_5175_out0 || v$G31_16112_out0;
assign v$G51_3675_out0 = v$NQ1_11550_out0 && v$F_2133_out0;
assign v$G51_3676_out0 = v$NQ1_11551_out0 && v$F_2134_out0;
assign v$G28_3947_out0 = ! v$F_2133_out0;
assign v$G28_3948_out0 = ! v$F_2134_out0;
assign v$IN_4527_out0 = v$OUT_3399_out0;
assign v$IN_4531_out0 = v$OUT_3403_out0;
assign v$_6592_out0 = { v$_15881_out0,v$_19155_out0 };
assign v$_6593_out0 = { v$_15882_out0,v$_19156_out0 };
assign v$XOR1_7919_out0 = v$C1_14151_out0 ^ v$MUX1_18540_out0;
assign v$XOR1_7923_out0 = v$C1_14155_out0 ^ v$MUX1_18544_out0;
assign v$G3_9161_out0 = v$HIGHER$SAME_15640_out0 && v$LOWER$OUT_4382_out0;
assign v$G3_9165_out0 = v$HIGHER$SAME_15644_out0 && v$LOWER$OUT_4386_out0;
assign v$DIFF_9414_out0 = v$A1_6076_out0;
assign v$DIFF_9418_out0 = v$A1_6080_out0;
assign v$NOT$USED1_14983_out0 = v$A1_6076_out1;
assign v$NOT$USED1_14987_out0 = v$A1_6080_out1;
assign v$MUX5_16091_out0 = v$IS$32$BITS_3203_out0 ? v$OUT_14344_out0 : v$OUT_14343_out0;
assign v$MUX5_16092_out0 = v$IS$32$BITS_3204_out0 ? v$OUT_14348_out0 : v$OUT_14347_out0;
assign v$_18048_out0 = { v$DIFF_9416_out0,v$C2_13910_out0 };
assign v$_18049_out0 = { v$DIFF_9420_out0,v$C2_13911_out0 };
assign v$SAME_19334_out0 = v$G1_9759_out0;
assign v$SAME_19338_out0 = v$G1_9760_out0;
assign v$SAME_19350_out0 = v$G1_9763_out0;
assign v$SAME_19354_out0 = v$G1_9764_out0;
assign v$LOWER$SAME_3975_out0 = v$SAME_19334_out0;
assign v$LOWER$SAME_3976_out0 = v$SAME_19338_out0;
assign v$LOWER$SAME_3977_out0 = v$SAME_19350_out0;
assign v$LOWER$SAME_3978_out0 = v$SAME_19354_out0;
assign v$OUT_4076_out0 = v$G30_1930_out0;
assign v$OUT_4080_out0 = v$G30_1933_out0;
assign v$OUT_4092_out0 = v$G30_1942_out0;
assign v$OUT_4096_out0 = v$G30_1945_out0;
assign {v$A1_6079_out1,v$A1_6079_out0 } = v$MUX3_3602_out0 + v$XOR1_7919_out0 + v$CIN_18829_out0;
assign {v$A1_6083_out1,v$A1_6083_out0 } = v$MUX3_3606_out0 + v$XOR1_7923_out0 + v$CIN_18833_out0;
assign v$_7938_out0 = { v$DIFF_9414_out0,v$C4_6859_out0 };
assign v$_7939_out0 = { v$DIFF_9418_out0,v$C4_6860_out0 };
assign v$A$EXP$LARGER_9815_out0 = v$MUX5_16091_out0;
assign v$A$EXP$LARGER_9816_out0 = v$MUX5_16092_out0;
assign v$IN_9949_out0 = v$IN_4527_out0;
assign v$IN_9953_out0 = v$IN_4531_out0;
assign v$G49_11564_out0 = v$G50_17963_out0 || v$G51_3675_out0;
assign v$G49_11565_out0 = v$G50_17964_out0 || v$G51_3676_out0;
assign v$G2_13477_out0 = v$HIGHER$OUT_4013_out0 || v$G3_9161_out0;
assign v$G2_13481_out0 = v$HIGHER$OUT_4017_out0 || v$G3_9165_out0;
assign v$NF_15164_out0 = v$G28_3947_out0;
assign v$NF_15165_out0 = v$G28_3948_out0;
assign v$G31_16098_out0 = v$A2$COMP$B2_2136_out0 || v$G32_412_out0;
assign v$G31_16099_out0 = v$A2$COMP$B2_2137_out0 || v$G32_413_out0;
assign v$G31_16101_out0 = v$A2$COMP$B2_2139_out0 || v$G32_415_out0;
assign v$G31_16102_out0 = v$A2$COMP$B2_2140_out0 || v$G32_416_out0;
assign v$G31_16110_out0 = v$A2$COMP$B2_2148_out0 || v$G32_424_out0;
assign v$G31_16111_out0 = v$A2$COMP$B2_2149_out0 || v$G32_425_out0;
assign v$G31_16113_out0 = v$A2$COMP$B2_2151_out0 || v$G32_427_out0;
assign v$G31_16114_out0 = v$A2$COMP$B2_2152_out0 || v$G32_428_out0;
assign v$_16778_out0 = { v$_6592_out0,v$C1_17454_out0 };
assign v$_16779_out0 = { v$_6593_out0,v$C1_17455_out0 };
assign v$G30_1931_out0 = v$A3$COMP$B3_5161_out0 || v$G31_16098_out0;
assign v$G30_1932_out0 = v$A3$COMP$B3_5162_out0 || v$G31_16099_out0;
assign v$G30_1934_out0 = v$A3$COMP$B3_5164_out0 || v$G31_16101_out0;
assign v$G30_1935_out0 = v$A3$COMP$B3_5165_out0 || v$G31_16102_out0;
assign v$G30_1943_out0 = v$A3$COMP$B3_5173_out0 || v$G31_16110_out0;
assign v$G30_1944_out0 = v$A3$COMP$B3_5174_out0 || v$G31_16111_out0;
assign v$G30_1946_out0 = v$A3$COMP$B3_5176_out0 || v$G31_16113_out0;
assign v$G30_1947_out0 = v$A3$COMP$B3_5177_out0 || v$G31_16114_out0;
assign v$G2_2058_out0 = v$EXP$SAME_17166_out0 || v$A$EXP$LARGER_9815_out0;
assign v$G2_2059_out0 = v$EXP$SAME_17167_out0 || v$A$EXP$LARGER_9816_out0;
assign v$Status_3973_out0 = v$_16778_out0;
assign v$Status_3974_out0 = v$_16779_out0;
assign v$OUT_4085_out0 = v$G2_13477_out0;
assign v$OUT_4101_out0 = v$G2_13481_out0;
assign v$_5016_out0 = v$IN_9949_out0[7:0];
assign v$_5020_out0 = v$IN_9953_out0[7:0];
assign v$_7794_out0 = v$IN_9949_out0[15:15];
assign v$_7795_out0 = v$IN_9953_out0[15:15];
assign v$HIGHER$OUT_8106_out0 = v$OUT_4076_out0;
assign v$HIGHER$OUT_8107_out0 = v$OUT_4080_out0;
assign v$HIGHER$OUT_8108_out0 = v$OUT_4092_out0;
assign v$HIGHER$OUT_8109_out0 = v$OUT_4096_out0;
assign v$DIFF_9417_out0 = v$A1_6079_out0;
assign v$DIFF_9421_out0 = v$A1_6083_out0;
assign v$_13855_out0 = v$IN_9949_out0[7:0];
assign v$_13858_out0 = v$IN_9953_out0[7:0];
assign v$_14705_out0 = v$IN_9949_out0[7:0];
assign v$_14706_out0 = v$IN_9953_out0[7:0];
assign v$NOT$USED1_14986_out0 = v$A1_6079_out1;
assign v$NOT$USED1_14990_out0 = v$A1_6083_out1;
assign v$_15204_out0 = v$IN_9949_out0[15:8];
assign v$_15208_out0 = v$IN_9953_out0[15:8];
assign v$_15240_out0 = v$IN_9949_out0[15:8];
assign v$_15244_out0 = v$IN_9953_out0[15:8];
assign v$IS$A$LARGER_15264_out0 = v$A$EXP$LARGER_9815_out0;
assign v$IS$A$LARGER_15265_out0 = v$A$EXP$LARGER_9816_out0;
assign v$G4_15927_out0 = v$EXP$SAME_17166_out0 || v$A$EXP$LARGER_9815_out0;
assign v$G4_15928_out0 = v$EXP$SAME_17167_out0 || v$A$EXP$LARGER_9816_out0;
assign v$_17371_out0 = v$IN_9949_out0[15:8];
assign v$_17375_out0 = v$IN_9953_out0[15:8];
assign v$G1_18090_out0 = v$LOWER$SAME_3975_out0 && v$HIGHER$SAME_9460_out0;
assign v$G1_18091_out0 = v$LOWER$SAME_3976_out0 && v$HIGHER$SAME_9461_out0;
assign v$G1_18092_out0 = v$LOWER$SAME_3977_out0 && v$HIGHER$SAME_9462_out0;
assign v$G1_18093_out0 = v$LOWER$SAME_3978_out0 && v$HIGHER$SAME_9463_out0;
assign v$G48_19127_out0 = v$NQ0_16214_out0 && v$G49_11564_out0;
assign v$G48_19128_out0 = v$NQ0_16215_out0 && v$G49_11565_out0;
assign v$_1632_out0 = { v$C1_8290_out0,v$_5016_out0 };
assign v$_1636_out0 = { v$C1_8294_out0,v$_5020_out0 };
assign v$MUX2_1765_out0 = v$IS$A$LARGER_15264_out0 ? v$SEL4_2485_out0 : v$SEL3_12468_out0;
assign v$MUX2_1766_out0 = v$IS$A$LARGER_15265_out0 ? v$SEL4_2486_out0 : v$SEL3_12469_out0;
assign v$MUX1_2096_out0 = v$IS$A$LARGER_15264_out0 ? v$SEL1_16347_out0 : v$SEL2_11519_out0;
assign v$MUX1_2097_out0 = v$IS$A$LARGER_15265_out0 ? v$SEL1_16348_out0 : v$SEL2_11520_out0;
assign v$MUX3_3600_out0 = v$OUT_4085_out0 ? v$A$EXP_297_out0 : v$B$EXP_17295_out0;
assign v$MUX3_3604_out0 = v$OUT_4101_out0 ? v$A$EXP_301_out0 : v$B$EXP_17299_out0;
assign v$OUT_4078_out0 = v$G30_1931_out0;
assign v$OUT_4079_out0 = v$G30_1932_out0;
assign v$OUT_4082_out0 = v$G30_1934_out0;
assign v$OUT_4083_out0 = v$G30_1935_out0;
assign v$OUT_4094_out0 = v$G30_1943_out0;
assign v$OUT_4095_out0 = v$G30_1944_out0;
assign v$OUT_4098_out0 = v$G30_1946_out0;
assign v$OUT_4099_out0 = v$G30_1947_out0;
assign v$MUX1_4198_out0 = v$G2_2058_out0 ? v$B_6781_out0 : v$A_2497_out0;
assign v$MUX1_4199_out0 = v$G2_2059_out0 ? v$B_6782_out0 : v$A_2498_out0;
assign v$MUX6_8275_out0 = v$IS$32$BITS_3203_out0 ? v$DIFF_9417_out0 : v$_18048_out0;
assign v$MUX6_8276_out0 = v$IS$32$BITS_3204_out0 ? v$DIFF_9421_out0 : v$_18049_out0;
assign v$STATUS_9155_out0 = v$Status_3973_out0;
assign v$STATUS_9156_out0 = v$Status_3974_out0;
assign v$SAME_9249_out0 = v$G1_18090_out0;
assign v$SAME_9250_out0 = v$G1_18091_out0;
assign v$SAME_9251_out0 = v$G1_18092_out0;
assign v$SAME_9252_out0 = v$G1_18093_out0;
assign v$_9822_out0 = { v$_17371_out0,v$LSBS_8263_out0 };
assign v$_9826_out0 = { v$_17375_out0,v$LSBS_8264_out0 };
assign v$_13893_out0 = { v$_15204_out0,v$_13855_out0 };
assign v$_13897_out0 = { v$_15208_out0,v$_13858_out0 };
assign v$MUX6_14288_out0 = v$S_18561_out0 ? v$_14705_out0 : v$C1_14033_out0;
assign v$MUX6_14289_out0 = v$S_18562_out0 ? v$_14706_out0 : v$C1_14034_out0;
assign v$OUT_14342_out0 = v$OUT_4085_out0;
assign v$OUT_14346_out0 = v$OUT_4101_out0;
assign v$MUX2_15790_out0 = v$G2_2058_out0 ? v$A_2497_out0 : v$B_6781_out0;
assign v$MUX2_15791_out0 = v$G2_2059_out0 ? v$A_2498_out0 : v$B_6782_out0;
assign v$MUX10_17440_out0 = v$G4_15927_out0 ? v$A_2497_out0 : v$B_6781_out0;
assign v$MUX10_17441_out0 = v$G4_15928_out0 ? v$A_2498_out0 : v$B_6782_out0;
assign v$G5_18490_out0 = v$G6_3383_out0 || v$G48_19127_out0;
assign v$G5_18491_out0 = v$G6_3384_out0 || v$G48_19128_out0;
assign v$MUX1_18538_out0 = v$OUT_4085_out0 ? v$B$EXP_17295_out0 : v$A$EXP_297_out0;
assign v$MUX1_18542_out0 = v$OUT_4101_out0 ? v$B$EXP_17299_out0 : v$A$EXP_301_out0;
assign v$MUX9_18555_out0 = v$G4_15927_out0 ? v$B_6781_out0 : v$A_2497_out0;
assign v$MUX9_18556_out0 = v$G4_15928_out0 ? v$B_6782_out0 : v$A_2498_out0;
assign v$_18585_out0 = { v$_7794_out0,v$_7794_out0 };
assign v$_18586_out0 = { v$_7795_out0,v$_7795_out0 };
assign v$SEL10_3221_out0 = v$MUX9_18555_out0[14:10];
assign v$SEL10_3222_out0 = v$MUX9_18556_out0[14:10];
assign v$SEL9_3955_out0 = v$MUX10_17440_out0[14:10];
assign v$SEL9_3956_out0 = v$MUX10_17441_out0[14:10];
assign v$HIGHER$OUT_4011_out0 = v$OUT_4078_out0;
assign v$HIGHER$OUT_4012_out0 = v$OUT_4082_out0;
assign v$HIGHER$OUT_4015_out0 = v$OUT_4094_out0;
assign v$HIGHER$OUT_4016_out0 = v$OUT_4098_out0;
assign v$LOWER$OUT_4380_out0 = v$OUT_4079_out0;
assign v$LOWER$OUT_4381_out0 = v$OUT_4083_out0;
assign v$LOWER$OUT_4384_out0 = v$OUT_4095_out0;
assign v$LOWER$OUT_4385_out0 = v$OUT_4099_out0;
assign v$MUX2_5066_out0 = v$IS$32$BIT_11362_out0 ? v$OUT_14342_out0 : v$OUT_14341_out0;
assign v$MUX2_5067_out0 = v$IS$32$BIT_11363_out0 ? v$OUT_14346_out0 : v$OUT_14345_out0;
assign v$XOR1_7917_out0 = v$C1_14149_out0 ^ v$MUX1_18538_out0;
assign v$XOR1_7921_out0 = v$C1_14153_out0 ^ v$MUX1_18542_out0;
assign v$MUX1_7971_out0 = v$G47_1685_out0 ? v$C1_1623_out0 : v$G5_18490_out0;
assign v$MUX1_7972_out0 = v$G47_1686_out0 ? v$C1_1624_out0 : v$G5_18491_out0;
assign v$SAME$H_9245_out0 = v$SAME_9249_out0;
assign v$SAME$H_9246_out0 = v$SAME_9251_out0;
assign v$_11523_out0 = { v$MUX2_1765_out0,v$C2_3818_out0 };
assign v$_11524_out0 = { v$MUX2_1766_out0,v$C2_3819_out0 };
assign v$SEL4_12764_out0 = v$MUX2_15790_out0[14:7];
assign v$SEL4_12765_out0 = v$MUX2_15791_out0[14:7];
assign v$EXP$DIFF_13064_out0 = v$MUX6_8275_out0;
assign v$EXP$DIFF_13065_out0 = v$MUX6_8276_out0;
assign v$_14703_out0 = { v$MUX1_2096_out0,v$C1_4520_out0 };
assign v$_14704_out0 = { v$MUX1_2097_out0,v$C1_4521_out0 };
assign v$MUX4_16603_out0 = v$EN_17564_out0 ? v$_1632_out0 : v$IN_9949_out0;
assign v$MUX4_16607_out0 = v$EN_17568_out0 ? v$_1636_out0 : v$IN_9953_out0;
assign v$SAME$L_17063_out0 = v$SAME_9250_out0;
assign v$SAME$L_17064_out0 = v$SAME_9252_out0;
assign v$_18052_out0 = { v$_18585_out0,v$_18585_out0 };
assign v$_18053_out0 = { v$_18586_out0,v$_18586_out0 };
assign v$MUX2_18372_out0 = v$FF2_9793_out0 ? v$STATUS_9155_out0 : v$RXBYTE_10010_out0;
assign v$MUX2_18373_out0 = v$FF2_9794_out0 ? v$STATUS_9156_out0 : v$RXBYTE_10011_out0;
assign v$SEL3_18423_out0 = v$MUX1_4198_out0[14:7];
assign v$SEL3_18424_out0 = v$MUX1_4199_out0[14:7];
assign v$SMALLER$EXP_3150_out0 = v$SEL10_3221_out0;
assign v$SMALLER$EXP_3151_out0 = v$SEL3_18423_out0;
assign v$SMALLER$EXP_3152_out0 = v$SEL10_3222_out0;
assign v$SMALLER$EXP_3153_out0 = v$SEL3_18424_out0;
assign {v$A1_6077_out1,v$A1_6077_out0 } = v$MUX3_3600_out0 + v$XOR1_7917_out0 + v$CIN_18827_out0;
assign {v$A1_6081_out1,v$A1_6081_out0 } = v$MUX3_3604_out0 + v$XOR1_7921_out0 + v$CIN_18831_out0;
assign v$_7193_out0 = { v$MUX2_18372_out0,v$C1_15419_out0 };
assign v$_7194_out0 = { v$MUX2_18373_out0,v$C1_15420_out0 };
assign v$G3_9159_out0 = v$HIGHER$SAME_15638_out0 && v$LOWER$OUT_4380_out0;
assign v$G3_9160_out0 = v$HIGHER$SAME_15639_out0 && v$LOWER$OUT_4381_out0;
assign v$G3_9163_out0 = v$HIGHER$SAME_15642_out0 && v$LOWER$OUT_4384_out0;
assign v$G3_9164_out0 = v$HIGHER$SAME_15643_out0 && v$LOWER$OUT_4385_out0;
assign v$LARGER$EXP_10729_out0 = v$SEL9_3955_out0;
assign v$LARGER$EXP_10730_out0 = v$SEL4_12764_out0;
assign v$LARGER$EXP_10731_out0 = v$SEL9_3956_out0;
assign v$LARGER$EXP_10732_out0 = v$SEL4_12765_out0;
assign v$MUX2_12606_out0 = v$G3_2803_out0 ? v$_9822_out0 : v$MUX4_16603_out0;
assign v$MUX2_12610_out0 = v$G3_2807_out0 ? v$_9826_out0 : v$MUX4_16607_out0;
assign v$IN_13746_out0 = v$_11523_out0;
assign v$IN_13750_out0 = v$_11524_out0;
assign v$_14916_out0 = { v$_18052_out0,v$_18052_out0 };
assign v$_14917_out0 = { v$_18053_out0,v$_18053_out0 };
assign v$EXP$DIFF_14934_out0 = v$EXP$DIFF_13064_out0;
assign v$EXP$DIFF_14935_out0 = v$EXP$DIFF_13065_out0;
assign v$SEL5_16783_out0 = v$_14703_out0[23:13];
assign v$SEL5_16784_out0 = v$_14704_out0[23:13];
assign v$Q0P_17393_out0 = v$MUX1_7971_out0;
assign v$Q0P_17394_out0 = v$MUX1_7972_out0;
assign v$DIFF_18144_out0 = v$EXP$DIFF_13064_out0;
assign v$DIFF_18145_out0 = v$EXP$DIFF_13064_out0;
assign v$DIFF_18146_out0 = v$EXP$DIFF_13065_out0;
assign v$DIFF_18147_out0 = v$EXP$DIFF_13065_out0;
assign v$A$EXP$LARGER_18846_out0 = v$MUX2_5066_out0;
assign v$A$EXP$LARGER_18847_out0 = v$MUX2_5067_out0;
assign v$G4_18881_out0 = v$SAME$L_17063_out0 && v$SAME$H_9245_out0;
assign v$G4_18882_out0 = v$SAME$L_17064_out0 && v$SAME$H_9246_out0;
assign v$MUX1_2159_out0 = v$FF1_11566_out0 ? v$_7193_out0 : v$RAMDOUT_17399_out0;
assign v$MUX1_2160_out0 = v$FF1_11567_out0 ? v$_7194_out0 : v$RAMDOUT_17400_out0;
assign v$IN_5387_out0 = v$IN_13746_out0;
assign v$IN_5418_out0 = v$IN_13750_out0;
assign v$SAME_6530_out0 = v$G4_18881_out0;
assign v$SAME_6531_out0 = v$G4_18882_out0;
assign v$DIFF_9415_out0 = v$A1_6077_out0;
assign v$DIFF_9419_out0 = v$A1_6081_out0;
assign v$_10464_out0 = { v$C4_2644_out0,v$SEL5_16783_out0 };
assign v$_10465_out0 = { v$C4_2645_out0,v$SEL5_16784_out0 };
assign v$G2_13475_out0 = v$HIGHER$OUT_4011_out0 || v$G3_9159_out0;
assign v$G2_13476_out0 = v$HIGHER$OUT_4012_out0 || v$G3_9160_out0;
assign v$G2_13479_out0 = v$HIGHER$OUT_4015_out0 || v$G3_9163_out0;
assign v$G2_13480_out0 = v$HIGHER$OUT_4016_out0 || v$G3_9164_out0;
assign v$MUX5_13753_out0 = v$FF1_8531_out0 ? v$LSBS_8263_out0 : v$_14916_out0;
assign v$MUX5_13754_out0 = v$FF1_8532_out0 ? v$LSBS_8264_out0 : v$_14917_out0;
assign v$N_14681_out0 = v$DIFF_18144_out0;
assign v$N_14682_out0 = v$DIFF_18145_out0;
assign v$N_14683_out0 = v$DIFF_18146_out0;
assign v$N_14684_out0 = v$DIFF_18147_out0;
assign v$NOT$USED1_14984_out0 = v$A1_6077_out1;
assign v$NOT$USED1_14988_out0 = v$A1_6081_out1;
assign v$_16748_out0 = { v$Q0P_17393_out0,v$Q1P_6027_out0 };
assign v$_16749_out0 = { v$Q0P_17394_out0,v$Q1P_6028_out0 };
assign v$EXP$DIFF_18281_out0 = v$EXP$DIFF_14934_out0;
assign v$EXP$DIFF_18282_out0 = v$EXP$DIFF_14935_out0;
assign v$MANTISA$SAME_2630_out0 = v$SAME_6530_out0;
assign v$MANTISA$SAME_2631_out0 = v$SAME_6531_out0;
assign v$MUX3_3320_out0 = v$IS$32$BITS_4307_out0 ? v$_14703_out0 : v$_10464_out0;
assign v$MUX3_3321_out0 = v$IS$32$BITS_4308_out0 ? v$_14704_out0 : v$_10465_out0;
assign v$RAMDOutOut_3407_out0 = v$MUX1_2159_out0;
assign v$RAMDOutOut_3408_out0 = v$MUX1_2160_out0;
assign v$IN_4041_out0 = v$IN_5387_out0;
assign v$IN_4050_out0 = v$IN_5418_out0;
assign v$OUT_4077_out0 = v$G2_13475_out0;
assign v$OUT_4081_out0 = v$G2_13476_out0;
assign v$OUT_4093_out0 = v$G2_13479_out0;
assign v$OUT_4097_out0 = v$G2_13480_out0;
assign v$SEL26_5050_out0 = v$N_14681_out0[7:5];
assign v$SEL26_5051_out0 = v$N_14682_out0[7:5];
assign v$SEL26_5052_out0 = v$N_14683_out0[7:5];
assign v$SEL26_5053_out0 = v$N_14684_out0[7:5];
assign v$SHIFT$AMOUNT_7705_out0 = v$EXP$DIFF_18281_out0;
assign v$SHIFT$AMOUNT_7709_out0 = v$EXP$DIFF_18282_out0;
assign v$_9807_out0 = { v$_16748_out0,v$_2866_out0 };
assign v$_9808_out0 = { v$_16749_out0,v$_2867_out0 };
assign v$MUX13_10825_out0 = v$IS$32$BIT_11362_out0 ? v$DIFF_9415_out0 : v$_7938_out0;
assign v$MUX13_10826_out0 = v$IS$32$BIT_11363_out0 ? v$DIFF_9419_out0 : v$_7939_out0;
assign v$_12383_out0 = { v$_15240_out0,v$MUX5_13753_out0 };
assign v$_12387_out0 = { v$_15244_out0,v$MUX5_13754_out0 };
assign v$SEL25_14039_out0 = v$N_14681_out0[4:0];
assign v$SEL25_14040_out0 = v$N_14682_out0[4:0];
assign v$SEL25_14041_out0 = v$N_14683_out0[4:0];
assign v$SEL25_14042_out0 = v$N_14684_out0[4:0];
assign v$SEL3_1284_out0 = v$SHIFT$AMOUNT_7705_out0[2:2];
assign v$SEL3_1288_out0 = v$SHIFT$AMOUNT_7709_out0[2:2];
assign v$SEL1_2478_out0 = v$SHIFT$AMOUNT_7705_out0[0:0];
assign v$SEL1_2482_out0 = v$SHIFT$AMOUNT_7709_out0[0:0];
assign v$OP1_4258_out0 = v$MUX3_3320_out0;
assign v$OP1_4259_out0 = v$MUX3_3321_out0;
assign v$SEL4_5155_out0 = v$SHIFT$AMOUNT_7705_out0[3:3];
assign v$SEL4_5159_out0 = v$SHIFT$AMOUNT_7709_out0[3:3];
assign v$SEL7_6599_out0 = v$SHIFT$AMOUNT_7705_out0[5:5];
assign v$SEL7_6603_out0 = v$SHIFT$AMOUNT_7709_out0[5:5];
assign v$LOWER$OUT_6665_out0 = v$OUT_4077_out0;
assign v$LOWER$OUT_6666_out0 = v$OUT_4081_out0;
assign v$LOWER$OUT_6667_out0 = v$OUT_4093_out0;
assign v$LOWER$OUT_6668_out0 = v$OUT_4097_out0;
assign v$MUX1_6917_out0 = v$G4_4189_out0 ? v$_12383_out0 : v$MUX2_12606_out0;
assign v$MUX1_6921_out0 = v$G4_4193_out0 ? v$_12387_out0 : v$MUX2_12610_out0;
assign v$SEL1_9068_out0 = v$IN_4041_out0[23:1];
assign v$SEL1_9099_out0 = v$IN_4050_out0[23:1];
assign v$SEL5_12784_out0 = v$SHIFT$AMOUNT_7705_out0[4:4];
assign v$SEL5_12788_out0 = v$SHIFT$AMOUNT_7709_out0[4:4];
assign v$DIFF_13242_out0 = v$MUX13_10825_out0;
assign v$DIFF_13243_out0 = v$MUX13_10826_out0;
assign v$SEL6_14368_out0 = v$SHIFT$AMOUNT_7705_out0[6:6];
assign v$SEL6_14372_out0 = v$SHIFT$AMOUNT_7709_out0[6:6];
assign v$SEL1_15996_out0 = v$IN_4041_out0[22:0];
assign v$SEL1_16027_out0 = v$IN_4050_out0[22:0];
assign v$N_16856_out0 = v$SEL25_14039_out0;
assign v$N_16857_out0 = v$SEL25_14040_out0;
assign v$N_16858_out0 = v$SEL25_14041_out0;
assign v$N_16859_out0 = v$SEL25_14042_out0;
assign v$SEL8_17193_out0 = v$SHIFT$AMOUNT_7705_out0[7:7];
assign v$SEL8_17197_out0 = v$SHIFT$AMOUNT_7709_out0[7:7];
assign v$NUPPER_18007_out0 = v$SEL26_5050_out0;
assign v$NUPPER_18008_out0 = v$SEL26_5051_out0;
assign v$NUPPER_18009_out0 = v$SEL26_5052_out0;
assign v$NUPPER_18010_out0 = v$SEL26_5053_out0;
assign v$UART$DOUT_18104_out0 = v$RAMDOutOut_3407_out0;
assign v$UART$DOUT_18105_out0 = v$RAMDOutOut_3408_out0;
assign v$SEL2_18963_out0 = v$SHIFT$AMOUNT_7705_out0[1:1];
assign v$SEL2_18967_out0 = v$SHIFT$AMOUNT_7709_out0[1:1];
assign v$DIFF_304_out0 = v$DIFF_13242_out0;
assign v$DIFF_305_out0 = v$DIFF_13243_out0;
assign v$EN_1500_out0 = v$SEL5_12784_out0;
assign v$EN_1501_out0 = v$SEL4_5155_out0;
assign v$EN_1510_out0 = v$SEL5_12788_out0;
assign v$EN_1511_out0 = v$SEL4_5159_out0;
assign v$EQ3_1977_out0 = v$N_16856_out0 == 5'h2;
assign v$EQ3_1978_out0 = v$N_16857_out0 == 5'h2;
assign v$EQ3_1979_out0 = v$N_16858_out0 == 5'h2;
assign v$EQ3_1980_out0 = v$N_16859_out0 == 5'h2;
assign v$MUX3_2125_out0 = v$G8_2053_out0 ? v$_13893_out0 : v$MUX1_6917_out0;
assign v$MUX3_2129_out0 = v$G8_2057_out0 ? v$_13897_out0 : v$MUX1_6921_out0;
assign v$EQ24_2732_out0 = v$N_16856_out0 == 5'h17;
assign v$EQ24_2733_out0 = v$N_16857_out0 == 5'h17;
assign v$EQ24_2734_out0 = v$N_16858_out0 == 5'h17;
assign v$EQ24_2735_out0 = v$N_16859_out0 == 5'h17;
assign v$EQ22_3060_out0 = v$N_16856_out0 == 5'h15;
assign v$EQ22_3061_out0 = v$N_16857_out0 == 5'h15;
assign v$EQ22_3062_out0 = v$N_16858_out0 == 5'h15;
assign v$EQ22_3063_out0 = v$N_16859_out0 == 5'h15;
assign v$EQ23_3415_out0 = v$N_16856_out0 == 5'h16;
assign v$EQ23_3416_out0 = v$N_16857_out0 == 5'h16;
assign v$EQ23_3417_out0 = v$N_16858_out0 == 5'h16;
assign v$EQ23_3418_out0 = v$N_16859_out0 == 5'h16;
assign v$EQ5_3537_out0 = v$N_16856_out0 == 5'h4;
assign v$EQ5_3538_out0 = v$N_16857_out0 == 5'h4;
assign v$EQ5_3539_out0 = v$N_16858_out0 == 5'h4;
assign v$EQ5_3540_out0 = v$N_16859_out0 == 5'h4;
assign v$EQ21_3547_out0 = v$N_16856_out0 == 5'h14;
assign v$EQ21_3548_out0 = v$N_16857_out0 == 5'h14;
assign v$EQ21_3549_out0 = v$N_16858_out0 == 5'h14;
assign v$EQ21_3550_out0 = v$N_16859_out0 == 5'h14;
assign v$A_3673_out0 = v$OP1_4258_out0;
assign v$A_3674_out0 = v$OP1_4259_out0;
assign v$EQ7_4242_out0 = v$N_16856_out0 == 5'h6;
assign v$EQ7_4243_out0 = v$N_16857_out0 == 5'h6;
assign v$EQ7_4244_out0 = v$N_16858_out0 == 5'h6;
assign v$EQ7_4245_out0 = v$N_16859_out0 == 5'h6;
assign v$_4428_out0 = { v$C2_126_out0,v$SEL1_15996_out0 };
assign v$_4459_out0 = { v$C2_157_out0,v$SEL1_16027_out0 };
assign v$EN_4967_out0 = v$SEL3_1284_out0;
assign v$EN_4973_out0 = v$SEL3_1288_out0;
assign v$EN_5431_out0 = v$SEL1_2478_out0;
assign v$EN_5437_out0 = v$SEL1_2482_out0;
assign v$EQ14_5642_out0 = v$N_16856_out0 == 5'hd;
assign v$EQ14_5643_out0 = v$N_16857_out0 == 5'hd;
assign v$EQ14_5644_out0 = v$N_16858_out0 == 5'hd;
assign v$EQ14_5645_out0 = v$N_16859_out0 == 5'hd;
assign v$EQ6_5666_out0 = v$N_16856_out0 == 5'h5;
assign v$EQ6_5667_out0 = v$N_16857_out0 == 5'h5;
assign v$EQ6_5668_out0 = v$N_16858_out0 == 5'h5;
assign v$EQ6_5669_out0 = v$N_16859_out0 == 5'h5;
assign v$EQ19_5682_out0 = v$N_16856_out0 == 5'h12;
assign v$EQ19_5683_out0 = v$N_16857_out0 == 5'h12;
assign v$EQ19_5684_out0 = v$N_16858_out0 == 5'h12;
assign v$EQ19_5685_out0 = v$N_16859_out0 == 5'h12;
assign v$EQ17_6155_out0 = v$N_16856_out0 == 5'h10;
assign v$EQ17_6156_out0 = v$N_16857_out0 == 5'h10;
assign v$EQ17_6157_out0 = v$N_16858_out0 == 5'h10;
assign v$EQ17_6158_out0 = v$N_16859_out0 == 5'h10;
assign v$EQ10_6169_out0 = v$N_16856_out0 == 5'h8;
assign v$EQ10_6170_out0 = v$N_16857_out0 == 5'h8;
assign v$EQ10_6171_out0 = v$N_16858_out0 == 5'h8;
assign v$EQ10_6172_out0 = v$N_16859_out0 == 5'h8;
assign v$EQ11_6408_out0 = v$N_16856_out0 == 5'ha;
assign v$EQ11_6409_out0 = v$N_16857_out0 == 5'ha;
assign v$EQ11_6410_out0 = v$N_16858_out0 == 5'ha;
assign v$EQ11_6411_out0 = v$N_16859_out0 == 5'ha;
assign v$SEL28_7645_out0 = v$NUPPER_18007_out0[1:1];
assign v$SEL28_7646_out0 = v$NUPPER_18008_out0[1:1];
assign v$SEL28_7647_out0 = v$NUPPER_18009_out0[1:1];
assign v$SEL28_7648_out0 = v$NUPPER_18010_out0[1:1];
assign v$EN_8203_out0 = v$SEL2_18963_out0;
assign v$EN_8209_out0 = v$SEL2_18967_out0;
assign v$RAMDOUT_8245_out0 = v$UART$DOUT_18104_out0;
assign v$RAMDOUT_8246_out0 = v$UART$DOUT_18105_out0;
assign v$EQ16_8597_out0 = v$N_16856_out0 == 5'hf;
assign v$EQ16_8598_out0 = v$N_16857_out0 == 5'hf;
assign v$EQ16_8599_out0 = v$N_16858_out0 == 5'hf;
assign v$EQ16_8600_out0 = v$N_16859_out0 == 5'hf;
assign v$_9329_out0 = { v$SEL1_9068_out0,v$C1_6264_out0 };
assign v$_9360_out0 = { v$SEL1_9099_out0,v$C1_6295_out0 };
assign v$EQ13_9893_out0 = v$N_16856_out0 == 5'hc;
assign v$EQ13_9894_out0 = v$N_16857_out0 == 5'hc;
assign v$EQ13_9895_out0 = v$N_16858_out0 == 5'hc;
assign v$EQ13_9896_out0 = v$N_16859_out0 == 5'hc;
assign v$EQ20_10370_out0 = v$N_16856_out0 == 5'h13;
assign v$EQ20_10371_out0 = v$N_16857_out0 == 5'h13;
assign v$EQ20_10372_out0 = v$N_16858_out0 == 5'h13;
assign v$EQ20_10373_out0 = v$N_16859_out0 == 5'h13;
assign v$EQ18_13375_out0 = v$N_16856_out0 == 5'h11;
assign v$EQ18_13376_out0 = v$N_16857_out0 == 5'h11;
assign v$EQ18_13377_out0 = v$N_16858_out0 == 5'h11;
assign v$EQ18_13378_out0 = v$N_16859_out0 == 5'h11;
assign v$EQ1_13999_out0 = v$N_16856_out0 == 5'h0;
assign v$EQ1_14000_out0 = v$N_16857_out0 == 5'h0;
assign v$EQ1_14001_out0 = v$N_16858_out0 == 5'h0;
assign v$EQ1_14002_out0 = v$N_16859_out0 == 5'h0;
assign v$EQ9_14361_out0 = v$N_16856_out0 == 5'h9;
assign v$EQ9_14362_out0 = v$N_16857_out0 == 5'h9;
assign v$EQ9_14363_out0 = v$N_16858_out0 == 5'h9;
assign v$EQ9_14364_out0 = v$N_16859_out0 == 5'h9;
assign v$EQ12_14427_out0 = v$N_16856_out0 == 5'hb;
assign v$EQ12_14428_out0 = v$N_16857_out0 == 5'hb;
assign v$EQ12_14429_out0 = v$N_16858_out0 == 5'hb;
assign v$EQ12_14430_out0 = v$N_16859_out0 == 5'hb;
assign v$EQ2_14810_out0 = v$N_16856_out0 == 5'h1;
assign v$EQ2_14811_out0 = v$N_16857_out0 == 5'h1;
assign v$EQ2_14812_out0 = v$N_16858_out0 == 5'h1;
assign v$EQ2_14813_out0 = v$N_16859_out0 == 5'h1;
assign v$EQ8_15018_out0 = v$N_16856_out0 == 5'h7;
assign v$EQ8_15019_out0 = v$N_16857_out0 == 5'h7;
assign v$EQ8_15020_out0 = v$N_16858_out0 == 5'h7;
assign v$EQ8_15021_out0 = v$N_16859_out0 == 5'h7;
assign v$EQ15_16574_out0 = v$N_16856_out0 == 5'he;
assign v$EQ15_16575_out0 = v$N_16857_out0 == 5'he;
assign v$EQ15_16576_out0 = v$N_16858_out0 == 5'he;
assign v$EQ15_16577_out0 = v$N_16859_out0 == 5'he;
assign v$G1_16646_out0 = v$SEL7_6599_out0 || v$SEL6_14368_out0;
assign v$G1_16650_out0 = v$SEL7_6603_out0 || v$SEL6_14372_out0;
assign v$SEL27_16918_out0 = v$NUPPER_18007_out0[0:0];
assign v$SEL27_16919_out0 = v$NUPPER_18008_out0[0:0];
assign v$SEL27_16920_out0 = v$NUPPER_18009_out0[0:0];
assign v$SEL27_16921_out0 = v$NUPPER_18010_out0[0:0];
assign v$SEL29_17214_out0 = v$NUPPER_18007_out0[2:2];
assign v$SEL29_17215_out0 = v$NUPPER_18008_out0[2:2];
assign v$SEL29_17216_out0 = v$NUPPER_18009_out0[2:2];
assign v$SEL29_17217_out0 = v$NUPPER_18010_out0[2:2];
assign v$G2_18840_out0 = v$HIGHER$SAME_9460_out0 && v$LOWER$OUT_6665_out0;
assign v$G2_18841_out0 = v$HIGHER$SAME_9461_out0 && v$LOWER$OUT_6666_out0;
assign v$G2_18842_out0 = v$HIGHER$SAME_9462_out0 && v$LOWER$OUT_6667_out0;
assign v$G2_18843_out0 = v$HIGHER$SAME_9463_out0 && v$LOWER$OUT_6668_out0;
assign v$EQ4_19209_out0 = v$N_16856_out0 == 5'h3;
assign v$EQ4_19210_out0 = v$N_16857_out0 == 5'h3;
assign v$EQ4_19211_out0 = v$N_16858_out0 == 5'h3;
assign v$EQ4_19212_out0 = v$N_16859_out0 == 5'h3;
assign v$RAMDOUT_68_out0 = v$RAMDOUT_8245_out0;
assign v$RAMDOUT_69_out0 = v$RAMDOUT_8246_out0;
assign v$MUX1_2565_out0 = v$LEFT$SHIT_3277_out0 ? v$_4428_out0 : v$_9329_out0;
assign v$MUX1_2596_out0 = v$LEFT$SHIT_3308_out0 ? v$_4459_out0 : v$_9360_out0;
assign v$DIFF_3044_out0 = v$DIFF_304_out0;
assign v$DIFF_3045_out0 = v$DIFF_305_out0;
assign v$OUT_3400_out0 = v$MUX3_2125_out0;
assign v$OUT_3404_out0 = v$MUX3_2129_out0;
assign v$G1_9137_out0 = v$SEL27_16918_out0 || v$SEL28_7645_out0;
assign v$G1_9138_out0 = v$SEL27_16919_out0 || v$SEL28_7646_out0;
assign v$G1_9139_out0 = v$SEL27_16920_out0 || v$SEL28_7647_out0;
assign v$G1_9140_out0 = v$SEL27_16921_out0 || v$SEL28_7648_out0;
assign v$G3_13637_out0 = v$HIGHER$OUT_8106_out0 || v$G2_18840_out0;
assign v$G3_13638_out0 = v$HIGHER$OUT_8107_out0 || v$G2_18841_out0;
assign v$G3_13639_out0 = v$HIGHER$OUT_8108_out0 || v$G2_18842_out0;
assign v$G3_13640_out0 = v$HIGHER$OUT_8109_out0 || v$G2_18843_out0;
assign v$A_14857_out0 = v$A_3673_out0;
assign v$A_14858_out0 = v$A_3674_out0;
assign v$G2_18057_out0 = v$G1_16646_out0 || v$SEL8_17193_out0;
assign v$G2_18061_out0 = v$G1_16650_out0 || v$SEL8_17197_out0;
assign v$RAMDOUT_5664_out0 = v$RAMDOUT_68_out0;
assign v$RAMDOUT_5665_out0 = v$RAMDOUT_69_out0;
assign v$SHIFT$AMOUNT_7702_out0 = v$DIFF_3044_out0;
assign v$SHIFT$AMOUNT_7703_out0 = v$DIFF_3044_out0;
assign v$SHIFT$AMOUNT_7706_out0 = v$DIFF_3045_out0;
assign v$SHIFT$AMOUNT_7707_out0 = v$DIFF_3045_out0;
assign v$OUT_9267_out0 = v$G3_13637_out0;
assign v$OUT_9268_out0 = v$G3_13638_out0;
assign v$OUT_9269_out0 = v$G3_13639_out0;
assign v$OUT_9270_out0 = v$G3_13640_out0;
assign v$SEL5_10785_out0 = v$A_14857_out0[23:1];
assign v$SEL5_10786_out0 = v$A_14858_out0[23:1];
assign v$G2_12476_out0 = v$G1_9137_out0 || v$SEL29_17214_out0;
assign v$G2_12477_out0 = v$G1_9138_out0 || v$SEL29_17215_out0;
assign v$G2_12478_out0 = v$G1_9139_out0 || v$SEL29_17216_out0;
assign v$G2_12479_out0 = v$G1_9140_out0 || v$SEL29_17217_out0;
assign v$OUT_15104_out0 = v$OUT_3400_out0;
assign v$OUT_15105_out0 = v$OUT_3404_out0;
assign v$MUX2_19189_out0 = v$EN_5431_out0 ? v$MUX1_2565_out0 : v$IN_4041_out0;
assign v$MUX2_19195_out0 = v$EN_5437_out0 ? v$MUX1_2596_out0 : v$IN_4050_out0;
assign v$SEL3_1281_out0 = v$SHIFT$AMOUNT_7702_out0[2:2];
assign v$SEL3_1282_out0 = v$SHIFT$AMOUNT_7703_out0[2:2];
assign v$SEL3_1285_out0 = v$SHIFT$AMOUNT_7706_out0[2:2];
assign v$SEL3_1286_out0 = v$SHIFT$AMOUNT_7707_out0[2:2];
assign v$_1303_out0 = { v$SEL5_10785_out0,v$C6_9182_out0 };
assign v$_1304_out0 = { v$SEL5_10786_out0,v$C6_9183_out0 };
assign v$SEL1_2475_out0 = v$SHIFT$AMOUNT_7702_out0[0:0];
assign v$SEL1_2476_out0 = v$SHIFT$AMOUNT_7703_out0[0:0];
assign v$SEL1_2479_out0 = v$SHIFT$AMOUNT_7706_out0[0:0];
assign v$SEL1_2480_out0 = v$SHIFT$AMOUNT_7707_out0[0:0];
assign v$G3_4935_out0 = v$OUT_9268_out0 && v$SAME$H_9245_out0;
assign v$G3_4936_out0 = v$OUT_9270_out0 && v$SAME$H_9246_out0;
assign v$SEL4_5152_out0 = v$SHIFT$AMOUNT_7702_out0[3:3];
assign v$SEL4_5153_out0 = v$SHIFT$AMOUNT_7703_out0[3:3];
assign v$SEL4_5156_out0 = v$SHIFT$AMOUNT_7706_out0[3:3];
assign v$SEL4_5157_out0 = v$SHIFT$AMOUNT_7707_out0[3:3];
assign v$SEL7_6596_out0 = v$SHIFT$AMOUNT_7702_out0[5:5];
assign v$SEL7_6597_out0 = v$SHIFT$AMOUNT_7703_out0[5:5];
assign v$SEL7_6600_out0 = v$SHIFT$AMOUNT_7706_out0[5:5];
assign v$SEL7_6601_out0 = v$SHIFT$AMOUNT_7707_out0[5:5];
assign v$OP2_10643_out0 = v$OUT_15104_out0;
assign v$OP2_10644_out0 = v$OUT_15105_out0;
assign v$MUX2_12557_out0 = v$G24_18545_out0 ? v$RAMDOUT_5664_out0 : v$RMN_6420_out0;
assign v$MUX2_12558_out0 = v$G24_18546_out0 ? v$RAMDOUT_5665_out0 : v$RMN_6421_out0;
assign v$SEL5_12781_out0 = v$SHIFT$AMOUNT_7702_out0[4:4];
assign v$SEL5_12782_out0 = v$SHIFT$AMOUNT_7703_out0[4:4];
assign v$SEL5_12785_out0 = v$SHIFT$AMOUNT_7706_out0[4:4];
assign v$SEL5_12786_out0 = v$SHIFT$AMOUNT_7707_out0[4:4];
assign v$SEL6_14365_out0 = v$SHIFT$AMOUNT_7702_out0[6:6];
assign v$SEL6_14366_out0 = v$SHIFT$AMOUNT_7703_out0[6:6];
assign v$SEL6_14369_out0 = v$SHIFT$AMOUNT_7706_out0[6:6];
assign v$SEL6_14370_out0 = v$SHIFT$AMOUNT_7707_out0[6:6];
assign v$OUT_15537_out0 = v$MUX2_19189_out0;
assign v$OUT_15568_out0 = v$MUX2_19195_out0;
assign v$SEL8_17190_out0 = v$SHIFT$AMOUNT_7702_out0[7:7];
assign v$SEL8_17191_out0 = v$SHIFT$AMOUNT_7703_out0[7:7];
assign v$SEL8_17194_out0 = v$SHIFT$AMOUNT_7706_out0[7:7];
assign v$SEL8_17195_out0 = v$SHIFT$AMOUNT_7707_out0[7:7];
assign v$SEL2_18960_out0 = v$SHIFT$AMOUNT_7702_out0[1:1];
assign v$SEL2_18961_out0 = v$SHIFT$AMOUNT_7703_out0[1:1];
assign v$SEL2_18964_out0 = v$SHIFT$AMOUNT_7706_out0[1:1];
assign v$SEL2_18965_out0 = v$SHIFT$AMOUNT_7707_out0[1:1];
assign v$EN_1493_out0 = v$SEL5_12781_out0;
assign v$EN_1494_out0 = v$SEL4_5152_out0;
assign v$EN_1495_out0 = v$SEL5_12782_out0;
assign v$EN_1496_out0 = v$SEL4_5153_out0;
assign v$EN_1503_out0 = v$SEL5_12785_out0;
assign v$EN_1504_out0 = v$SEL4_5156_out0;
assign v$EN_1505_out0 = v$SEL5_12786_out0;
assign v$EN_1506_out0 = v$SEL4_5157_out0;
assign v$EN_4963_out0 = v$SEL3_1281_out0;
assign v$EN_4964_out0 = v$SEL3_1282_out0;
assign v$EN_4969_out0 = v$SEL3_1285_out0;
assign v$EN_4970_out0 = v$SEL3_1286_out0;
assign v$IN_5389_out0 = v$OUT_15537_out0;
assign v$IN_5420_out0 = v$OUT_15568_out0;
assign v$EN_5427_out0 = v$SEL1_2475_out0;
assign v$EN_5428_out0 = v$SEL1_2476_out0;
assign v$EN_5433_out0 = v$SEL1_2479_out0;
assign v$EN_5434_out0 = v$SEL1_2480_out0;
assign v$EN_8199_out0 = v$SEL2_18960_out0;
assign v$EN_8200_out0 = v$SEL2_18961_out0;
assign v$EN_8205_out0 = v$SEL2_18964_out0;
assign v$EN_8206_out0 = v$SEL2_18965_out0;
assign v$OP2_15675_out0 = v$OP2_10643_out0;
assign v$OP2_15676_out0 = v$OP2_10644_out0;
assign v$G1_16179_out0 = v$G3_4935_out0 || v$OUT_9267_out0;
assign v$G1_16180_out0 = v$G3_4936_out0 || v$OUT_9269_out0;
assign v$G1_16643_out0 = v$SEL7_6596_out0 || v$SEL6_14365_out0;
assign v$G1_16644_out0 = v$SEL7_6597_out0 || v$SEL6_14366_out0;
assign v$G1_16647_out0 = v$SEL7_6600_out0 || v$SEL6_14369_out0;
assign v$G1_16648_out0 = v$SEL7_6601_out0 || v$SEL6_14370_out0;
assign v$REGDIN_18984_out0 = v$MUX2_12557_out0;
assign v$REGDIN_18985_out0 = v$MUX2_12558_out0;
assign v$OUT_4021_out0 = v$G1_16179_out0;
assign v$OUT_4022_out0 = v$G1_16180_out0;
assign v$OP2_7906_out0 = v$OP2_15675_out0;
assign v$OP2_7907_out0 = v$OP2_15676_out0;
assign v$IN_12356_out0 = v$IN_5389_out0;
assign v$IN_12362_out0 = v$IN_5420_out0;
assign v$REGDIN_17124_out0 = v$REGDIN_18984_out0;
assign v$REGDIN_17125_out0 = v$REGDIN_18985_out0;
assign v$G2_18054_out0 = v$G1_16643_out0 || v$SEL8_17190_out0;
assign v$G2_18055_out0 = v$G1_16644_out0 || v$SEL8_17191_out0;
assign v$G2_18058_out0 = v$G1_16647_out0 || v$SEL8_17194_out0;
assign v$G2_18059_out0 = v$G1_16648_out0 || v$SEL8_17195_out0;
assign v$SEL1_9070_out0 = v$IN_12356_out0[23:2];
assign v$SEL1_9101_out0 = v$IN_12362_out0[23:2];
assign v$XOR1_9920_out0 = v$OP2_7906_out0 ^ v$MUX1_18336_out0;
assign v$XOR1_9921_out0 = v$OP2_7907_out0 ^ v$MUX1_18337_out0;
assign v$B_12288_out0 = v$OP2_7906_out0;
assign v$B_12289_out0 = v$OP2_7907_out0;
assign v$SEL1_15998_out0 = v$IN_12356_out0[21:0];
assign v$SEL1_16029_out0 = v$IN_12362_out0[21:0];
assign v$A$MANTISA$LARGER_16641_out0 = v$OUT_4021_out0;
assign v$A$MANTISA$LARGER_16642_out0 = v$OUT_4022_out0;
assign v$_4430_out0 = { v$C2_128_out0,v$SEL1_15998_out0 };
assign v$_4461_out0 = { v$C2_159_out0,v$SEL1_16029_out0 };
assign v$_9331_out0 = { v$SEL1_9070_out0,v$C1_6266_out0 };
assign v$_9362_out0 = { v$SEL1_9101_out0,v$C1_6297_out0 };
assign {v$A1_9805_out1,v$A1_9805_out0 } = v$OP1_5658_out0 + v$XOR1_9920_out0 + v$MUX2_12801_out0;
assign {v$A1_9806_out1,v$A1_9806_out0 } = v$OP1_5659_out0 + v$XOR1_9921_out0 + v$MUX2_12802_out0;
assign v$B_10432_out0 = v$B_12288_out0;
assign v$B_10433_out0 = v$B_12289_out0;
assign v$G7_19251_out0 = v$A$MANTISA$LARGER_16641_out0 && v$EXP$SAME_1006_out0;
assign v$G7_19252_out0 = v$A$MANTISA$LARGER_16642_out0 && v$EXP$SAME_1007_out0;
assign v$MUX1_2567_out0 = v$LEFT$SHIT_3279_out0 ? v$_4430_out0 : v$_9331_out0;
assign v$MUX1_2598_out0 = v$LEFT$SHIT_3310_out0 ? v$_4461_out0 : v$_9362_out0;
assign v$ADDEROUT_3704_out0 = v$A1_9805_out0;
assign v$ADDEROUT_3705_out0 = v$A1_9806_out0;
assign v$_5447_out0 = v$B_10432_out0[7:4];
assign v$_5448_out0 = v$B_10433_out0[7:4];
assign v$_6594_out0 = v$B_10432_out0[11:8];
assign v$_6595_out0 = v$B_10433_out0[11:8];
assign v$G9_17527_out0 = v$A$EXP$LARGER_18846_out0 || v$G7_19251_out0;
assign v$G9_17528_out0 = v$A$EXP$LARGER_18847_out0 || v$G7_19252_out0;
assign v$_18850_out0 = v$B_10432_out0[15:12];
assign v$_18851_out0 = v$B_10433_out0[15:12];
assign v$_19217_out0 = v$B_10432_out0[3:0];
assign v$_19218_out0 = v$B_10433_out0[3:0];
assign v$_56_out0 = v$_19217_out0[1:0];
assign v$_56_out1 = v$_19217_out0[3:2];
assign v$_57_out0 = v$_19218_out0[1:0];
assign v$_57_out1 = v$_19218_out0[3:2];
assign v$_237_out0 = v$_5447_out0[1:0];
assign v$_237_out1 = v$_5447_out0[3:2];
assign v$_238_out0 = v$_5448_out0[1:0];
assign v$_238_out1 = v$_5448_out0[3:2];
assign v$_1625_out0 = v$_18850_out0[1:0];
assign v$_1625_out1 = v$_18850_out0[3:2];
assign v$_1626_out0 = v$_18851_out0[1:0];
assign v$_1626_out1 = v$_18851_out0[3:2];
assign v$MUX2_2674_out0 = v$EN_8203_out0 ? v$MUX1_2567_out0 : v$IN_12356_out0;
assign v$MUX2_2680_out0 = v$EN_8209_out0 ? v$MUX1_2598_out0 : v$IN_12362_out0;
assign v$_7786_out0 = v$_6594_out0[1:0];
assign v$_7786_out1 = v$_6594_out0[3:2];
assign v$_7787_out0 = v$_6595_out0[1:0];
assign v$_7787_out1 = v$_6595_out0[3:2];
assign v$IS$A$LARGER_17444_out0 = v$G9_17527_out0;
assign v$IS$A$LARGER_17445_out0 = v$G9_17528_out0;
assign v$G8_255_out0 = v$IS$A$LARGER_17444_out0 || v$IS$SUB_4611_out0;
assign v$G8_256_out0 = v$IS$A$LARGER_17445_out0 || v$IS$SUB_4612_out0;
assign v$MUX11_1353_out0 = v$IS$A$LARGER_17444_out0 ? v$SEL5_326_out0 : v$G1_15752_out0;
assign v$MUX11_1354_out0 = v$IS$A$LARGER_17445_out0 ? v$SEL5_327_out0 : v$G1_15753_out0;
assign v$_5255_out0 = v$_56_out1[0:0];
assign v$_5255_out1 = v$_56_out1[1:1];
assign v$_5256_out0 = v$_57_out1[0:0];
assign v$_5256_out1 = v$_57_out1[1:1];
assign v$MUX15_7291_out0 = v$IS$A$LARGER_17444_out0 ? v$A_3465_out0 : v$B_18356_out0;
assign v$MUX15_7292_out0 = v$IS$A$LARGER_17445_out0 ? v$A_3466_out0 : v$B_18357_out0;
assign v$IS$A$LARGER_7361_out0 = v$IS$A$LARGER_17444_out0;
assign v$IS$A$LARGER_7362_out0 = v$IS$A$LARGER_17445_out0;
assign v$_7710_out0 = v$_237_out1[0:0];
assign v$_7710_out1 = v$_237_out1[1:1];
assign v$_7711_out0 = v$_238_out1[0:0];
assign v$_7711_out1 = v$_238_out1[1:1];
assign v$_9398_out0 = v$_237_out0[0:0];
assign v$_9398_out1 = v$_237_out0[1:1];
assign v$_9399_out0 = v$_238_out0[0:0];
assign v$_9399_out1 = v$_238_out0[1:1];
assign v$_9437_out0 = v$_7786_out0[0:0];
assign v$_9437_out1 = v$_7786_out0[1:1];
assign v$_9438_out0 = v$_7787_out0[0:0];
assign v$_9438_out1 = v$_7787_out0[1:1];
assign v$_15249_out0 = v$_56_out0[0:0];
assign v$_15249_out1 = v$_56_out0[1:1];
assign v$_15250_out0 = v$_57_out0[0:0];
assign v$_15250_out1 = v$_57_out0[1:1];
assign v$OUT_15539_out0 = v$MUX2_2674_out0;
assign v$OUT_15570_out0 = v$MUX2_2680_out0;
assign v$_15788_out0 = v$_1625_out0[0:0];
assign v$_15788_out1 = v$_1625_out0[1:1];
assign v$_15789_out0 = v$_1626_out0[0:0];
assign v$_15789_out1 = v$_1626_out0[1:1];
assign v$_15905_out0 = v$_1625_out1[0:0];
assign v$_15905_out1 = v$_1625_out1[1:1];
assign v$_15906_out0 = v$_1626_out1[0:0];
assign v$_15906_out1 = v$_1626_out1[1:1];
assign v$G2_16133_out0 = v$IS$A$LARGER_17444_out0 && v$IS$SUB_4611_out0;
assign v$G2_16134_out0 = v$IS$A$LARGER_17445_out0 && v$IS$SUB_4612_out0;
assign v$_16750_out0 = v$_7786_out1[0:0];
assign v$_16750_out1 = v$_7786_out1[1:1];
assign v$_16751_out0 = v$_7787_out1[0:0];
assign v$_16751_out1 = v$_7787_out1[1:1];
assign v$MUX16_19139_out0 = v$IS$A$LARGER_17444_out0 ? v$A_3465_out0 : v$B_18356_out0;
assign v$MUX16_19140_out0 = v$IS$A$LARGER_17445_out0 ? v$A_3466_out0 : v$B_18357_out0;
assign v$G14_1831_out0 = v$_17170_out1 && v$_15788_out1;
assign v$G14_1832_out0 = v$_17171_out1 && v$_15789_out1;
assign v$G13_1847_out0 = v$_17170_out0 && v$_15788_out0;
assign v$G13_1848_out0 = v$_17171_out0 && v$_15789_out0;
assign v$G5_2440_out0 = v$_4176_out0 && v$_9398_out0;
assign v$G5_2441_out0 = v$_4177_out0 && v$_9399_out0;
assign v$G6_2452_out0 = v$_4176_out1 && v$_9398_out1;
assign v$G6_2453_out0 = v$_4177_out1 && v$_9399_out1;
assign v$G9_3651_out0 = v$_346_out0 && v$_9437_out0;
assign v$G9_3652_out0 = v$_347_out0 && v$_9438_out0;
assign v$A$IS$OP1_5221_out0 = v$G8_255_out0;
assign v$A$IS$OP1_5222_out0 = v$G8_256_out0;
assign v$IN_5388_out0 = v$OUT_15539_out0;
assign v$IN_5419_out0 = v$OUT_15570_out0;
assign v$SEL17_5630_out0 = v$MUX16_19139_out0[14:7];
assign v$SEL17_5631_out0 = v$MUX16_19140_out0[14:7];
assign v$G11_8511_out0 = v$_5108_out0 && v$_16750_out0;
assign v$G11_8512_out0 = v$_5109_out0 && v$_16751_out0;
assign v$G2_9406_out0 = v$_11568_out1 && v$_15249_out1;
assign v$G2_9407_out0 = v$_11569_out1 && v$_15250_out1;
assign v$G8_9410_out0 = v$_10697_out1 && v$_7710_out1;
assign v$G8_9411_out0 = v$_10698_out1 && v$_7711_out1;
assign v$IS$A$LARGER_10896_out0 = v$IS$A$LARGER_7361_out0;
assign v$IS$A$LARGER_10897_out0 = v$IS$A$LARGER_7362_out0;
assign v$G4_12443_out0 = v$G2_16133_out0 && v$G5_16393_out0;
assign v$G4_12444_out0 = v$G2_16134_out0 && v$G5_16394_out0;
assign v$SUBTRACTION$SIGN_12445_out0 = v$MUX11_1353_out0;
assign v$SUBTRACTION$SIGN_12446_out0 = v$MUX11_1354_out0;
assign v$G1_12690_out0 = v$_11568_out0 && v$_15249_out0;
assign v$G1_12691_out0 = v$_11569_out0 && v$_15250_out0;
assign v$G7_12768_out0 = v$_10697_out0 && v$_7710_out0;
assign v$G7_12769_out0 = v$_10698_out0 && v$_7711_out0;
assign v$G3_13520_out0 = v$_5646_out0 && v$_5255_out0;
assign v$G3_13521_out0 = v$_5647_out0 && v$_5256_out0;
assign v$G12_14383_out0 = v$_5108_out1 && v$_16750_out1;
assign v$G12_14384_out0 = v$_5109_out1 && v$_16751_out1;
assign v$G4_15100_out0 = v$_5646_out1 && v$_5255_out1;
assign v$G4_15101_out0 = v$_5647_out1 && v$_5256_out1;
assign v$G15_15183_out0 = v$_3332_out0 && v$_15905_out0;
assign v$G15_15184_out0 = v$_3333_out0 && v$_15906_out0;
assign v$SEL3_18385_out0 = v$MUX15_7291_out0[14:7];
assign v$SEL3_18386_out0 = v$MUX15_7292_out0[14:7];
assign v$SEL18_18852_out0 = v$MUX16_19139_out0[14:10];
assign v$SEL18_18853_out0 = v$MUX16_19140_out0[14:10];
assign v$G10_19095_out0 = v$_346_out1 && v$_9437_out1;
assign v$G10_19096_out0 = v$_347_out1 && v$_9438_out1;
assign v$G16_19392_out0 = v$_3332_out1 && v$_15905_out1;
assign v$G16_19393_out0 = v$_3333_out1 && v$_15906_out1;
assign v$MUX9_2652_out0 = v$A$IS$OP1_5221_out0 ? v$B$MANTISA_16181_out0 : v$A$MANTISA_3937_out0;
assign v$MUX9_2653_out0 = v$A$IS$OP1_5222_out0 ? v$B$MANTISA_16182_out0 : v$A$MANTISA_3938_out0;
assign v$_3363_out0 = { v$G15_15183_out0,v$G16_19392_out0 };
assign v$_3364_out0 = { v$G15_15184_out0,v$G16_19393_out0 };
assign v$_9831_out0 = { v$G7_12768_out0,v$G8_9410_out0 };
assign v$_9832_out0 = { v$G7_12769_out0,v$G8_9411_out0 };
assign v$_11481_out0 = { v$G3_13520_out0,v$G4_15100_out0 };
assign v$_11482_out0 = { v$G3_13521_out0,v$G4_15101_out0 };
assign v$SINGLE$PRECISION$EXPONENT_11558_out0 = v$SEL3_18385_out0;
assign v$SINGLE$PRECISION$EXPONENT_11559_out0 = v$SEL3_18386_out0;
assign v$MUX3_13369_out0 = v$A$IS$OP1_5221_out0 ? v$A$MANTISA_3937_out0 : v$B$MANTISA_16181_out0;
assign v$MUX3_13370_out0 = v$A$IS$OP1_5222_out0 ? v$A$MANTISA_3938_out0 : v$B$MANTISA_16182_out0;
assign v$EXPONENT_14267_out0 = v$SEL17_5630_out0;
assign v$EXPONENT_14268_out0 = v$SEL17_5631_out0;
assign v$_14779_out0 = { v$G1_12690_out0,v$G2_9406_out0 };
assign v$_14780_out0 = { v$G1_12691_out0,v$G2_9407_out0 };
assign v$_14814_out0 = { v$G5_2440_out0,v$G6_2452_out0 };
assign v$_14815_out0 = { v$G5_2441_out0,v$G6_2453_out0 };
assign v$IN_16200_out0 = v$IN_5388_out0;
assign v$IN_16206_out0 = v$IN_5419_out0;
assign v$G1_16383_out0 = ! v$IS$A$LARGER_10896_out0;
assign v$G1_16384_out0 = ! v$IS$A$LARGER_10897_out0;
assign v$_16610_out0 = { v$G11_8511_out0,v$G12_14383_out0 };
assign v$_16611_out0 = { v$G11_8512_out0,v$G12_14384_out0 };
assign v$EXPONENT_16622_out0 = v$SEL18_18852_out0;
assign v$EXPONENT_16623_out0 = v$SEL18_18853_out0;
assign v$_17395_out0 = { v$G9_3651_out0,v$G10_19095_out0 };
assign v$_17396_out0 = { v$G9_3652_out0,v$G10_19096_out0 };
assign v$MUX4_18328_out0 = v$G4_12443_out0 ? v$A_3465_out0 : v$B_18356_out0;
assign v$MUX4_18329_out0 = v$G4_12444_out0 ? v$A_3466_out0 : v$B_18357_out0;
assign v$_19177_out0 = { v$G13_1847_out0,v$G14_1831_out0 };
assign v$_19178_out0 = { v$G13_1848_out0,v$G14_1832_out0 };
assign v$_267_out0 = { v$_19177_out0,v$_3363_out0 };
assign v$_268_out0 = { v$_19178_out0,v$_3364_out0 };
assign v$EXPONENT_1521_out0 = v$SINGLE$PRECISION$EXPONENT_11558_out0;
assign v$EXPONENT_1522_out0 = v$SINGLE$PRECISION$EXPONENT_11559_out0;
assign v$_3887_out0 = { v$_17395_out0,v$_16610_out0 };
assign v$_3888_out0 = { v$_17396_out0,v$_16611_out0 };
assign v$SEL1_9069_out0 = v$IN_16200_out0[23:4];
assign v$SEL1_9100_out0 = v$IN_16206_out0[23:4];
assign v$OP1$MANTISA_9449_out0 = v$MUX3_13369_out0;
assign v$OP1$MANTISA_9450_out0 = v$MUX3_13370_out0;
assign v$SEL1_9839_out0 = v$MUX4_18328_out0[14:10];
assign v$SEL1_9840_out0 = v$MUX4_18329_out0[14:10];
assign v$OP2$MANTISA_9922_out0 = v$MUX9_2652_out0;
assign v$OP2$MANTISA_9923_out0 = v$MUX9_2653_out0;
assign v$_13589_out0 = { v$_14814_out0,v$_9831_out0 };
assign v$_13590_out0 = { v$_14815_out0,v$_9832_out0 };
assign v$SEL1_15997_out0 = v$IN_16200_out0[19:0];
assign v$SEL1_16028_out0 = v$IN_16206_out0[19:0];
assign v$G2_17128_out0 = v$IS$SUB_13643_out0 && v$G1_16383_out0;
assign v$G2_17129_out0 = v$IS$SUB_13644_out0 && v$G1_16384_out0;
assign v$_17497_out0 = { v$_14779_out0,v$_11481_out0 };
assign v$_17498_out0 = { v$_14780_out0,v$_11482_out0 };
assign v$C0_208_out0 = v$_17497_out0;
assign v$C0_209_out0 = v$_17498_out0;
assign v$OP2$MANTISA_2853_out0 = v$OP2$MANTISA_9922_out0;
assign v$OP2$MANTISA_2854_out0 = v$OP2$MANTISA_9923_out0;
assign v$C12_3507_out0 = v$_267_out0;
assign v$C12_3508_out0 = v$_268_out0;
assign v$OP1$MANTISA_3971_out0 = v$OP1$MANTISA_9449_out0;
assign v$OP1$MANTISA_3972_out0 = v$OP1$MANTISA_9450_out0;
assign v$_4429_out0 = { v$C2_127_out0,v$SEL1_15997_out0 };
assign v$_4460_out0 = { v$C2_158_out0,v$SEL1_16028_out0 };
assign v$NEED$SHIFT$OP1_5034_out0 = v$G2_17128_out0;
assign v$NEED$SHIFT$OP1_5035_out0 = v$G2_17129_out0;
assign v$HALF$PRECISION$EXPONENT_6622_out0 = v$SEL1_9839_out0;
assign v$HALF$PRECISION$EXPONENT_6623_out0 = v$SEL1_9840_out0;
assign v$C8_8637_out0 = v$_3887_out0;
assign v$C8_8638_out0 = v$_3888_out0;
assign v$_9330_out0 = { v$SEL1_9069_out0,v$C1_6265_out0 };
assign v$_9361_out0 = { v$SEL1_9100_out0,v$C1_6296_out0 };
assign v$C4_11272_out0 = v$_13589_out0;
assign v$C4_11273_out0 = v$_13590_out0;
assign v$MUX1_2566_out0 = v$LEFT$SHIT_3278_out0 ? v$_4429_out0 : v$_9330_out0;
assign v$MUX1_2597_out0 = v$LEFT$SHIT_3309_out0 ? v$_4460_out0 : v$_9361_out0;
assign v$OP2$MANTISA_3710_out0 = v$OP2$MANTISA_2853_out0;
assign v$OP2$MANTISA_3711_out0 = v$OP2$MANTISA_2854_out0;
assign v$_3866_out0 = { v$C0_208_out0,v$C4_11272_out0 };
assign v$_3867_out0 = { v$C0_209_out0,v$C4_11273_out0 };
assign v$_9369_out0 = { v$C8_8637_out0,v$C12_3507_out0 };
assign v$_9370_out0 = { v$C8_8638_out0,v$C12_3508_out0 };
assign v$OP1$MANTISA_12378_out0 = v$OP1$MANTISA_3971_out0;
assign v$OP1$MANTISA_12379_out0 = v$OP1$MANTISA_3972_out0;
assign v$EXPONENT_17014_out0 = v$HALF$PRECISION$EXPONENT_6622_out0;
assign v$EXPONENT_17015_out0 = v$HALF$PRECISION$EXPONENT_6623_out0;
assign v$IN_13743_out0 = v$OP2$MANTISA_3710_out0;
assign v$IN_13744_out0 = v$OP1$MANTISA_12378_out0;
assign v$IN_13747_out0 = v$OP2$MANTISA_3711_out0;
assign v$IN_13748_out0 = v$OP1$MANTISA_12379_out0;
assign v$MUX2_15821_out0 = v$EN_4967_out0 ? v$MUX1_2566_out0 : v$IN_16200_out0;
assign v$MUX2_15827_out0 = v$EN_4973_out0 ? v$MUX1_2597_out0 : v$IN_16206_out0;
assign v$_16987_out0 = { v$_3866_out0,v$_9369_out0 };
assign v$_16988_out0 = { v$_3867_out0,v$_9370_out0 };
assign v$IN_5367_out0 = v$IN_13743_out0;
assign v$IN_5372_out0 = v$IN_13744_out0;
assign v$IN_5398_out0 = v$IN_13747_out0;
assign v$IN_5403_out0 = v$IN_13748_out0;
assign v$OUT_15538_out0 = v$MUX2_15821_out0;
assign v$OUT_15569_out0 = v$MUX2_15827_out0;
assign v$C_18715_out0 = v$_16987_out0;
assign v$C_18716_out0 = v$_16988_out0;
assign v$IN_4036_out0 = v$IN_5367_out0;
assign v$IN_4037_out0 = v$IN_5372_out0;
assign v$IN_4045_out0 = v$IN_5398_out0;
assign v$IN_4046_out0 = v$IN_5403_out0;
assign v$IN_5386_out0 = v$OUT_15538_out0;
assign v$IN_5417_out0 = v$OUT_15569_out0;
assign v$ANDOUT_7689_out0 = v$C_18715_out0;
assign v$ANDOUT_7690_out0 = v$C_18716_out0;
assign v$MUX3_4062_out0 = v$G6_6224_out0 ? v$ANDOUT_7689_out0 : v$ADDEROUT_3704_out0;
assign v$MUX3_4063_out0 = v$G6_6225_out0 ? v$ANDOUT_7690_out0 : v$ADDEROUT_3705_out0;
assign v$IN_5241_out0 = v$IN_5386_out0;
assign v$IN_5251_out0 = v$IN_5417_out0;
assign v$SEL1_9048_out0 = v$IN_4036_out0[23:1];
assign v$SEL1_9053_out0 = v$IN_4037_out0[23:1];
assign v$SEL1_9079_out0 = v$IN_4045_out0[23:1];
assign v$SEL1_9084_out0 = v$IN_4046_out0[23:1];
assign v$SEL1_15976_out0 = v$IN_4036_out0[22:0];
assign v$SEL1_15981_out0 = v$IN_4037_out0[22:0];
assign v$SEL1_16007_out0 = v$IN_4045_out0[22:0];
assign v$SEL1_16012_out0 = v$IN_4046_out0[22:0];
assign v$_4408_out0 = { v$C2_106_out0,v$SEL1_15976_out0 };
assign v$_4413_out0 = { v$C2_111_out0,v$SEL1_15981_out0 };
assign v$_4439_out0 = { v$C2_137_out0,v$SEL1_16007_out0 };
assign v$_4444_out0 = { v$C2_142_out0,v$SEL1_16012_out0 };
assign v$MUX4_6214_out0 = v$EQ1_2712_out0 ? v$OP2_7906_out0 : v$MUX3_4062_out0;
assign v$MUX4_6215_out0 = v$EQ1_2713_out0 ? v$OP2_7907_out0 : v$MUX3_4063_out0;
assign v$SEL1_9067_out0 = v$IN_5241_out0[23:8];
assign v$SEL1_9098_out0 = v$IN_5251_out0[23:8];
assign v$_9309_out0 = { v$SEL1_9048_out0,v$C1_6244_out0 };
assign v$_9314_out0 = { v$SEL1_9053_out0,v$C1_6249_out0 };
assign v$_9340_out0 = { v$SEL1_9079_out0,v$C1_6275_out0 };
assign v$_9345_out0 = { v$SEL1_9084_out0,v$C1_6280_out0 };
assign v$SEL1_15995_out0 = v$IN_5241_out0[15:0];
assign v$SEL1_16026_out0 = v$IN_5251_out0[15:0];
assign v$MUX1_2545_out0 = v$LEFT$SHIT_3257_out0 ? v$_4408_out0 : v$_9309_out0;
assign v$MUX1_2550_out0 = v$LEFT$SHIT_3262_out0 ? v$_4413_out0 : v$_9314_out0;
assign v$MUX1_2576_out0 = v$LEFT$SHIT_3288_out0 ? v$_4439_out0 : v$_9340_out0;
assign v$MUX1_2581_out0 = v$LEFT$SHIT_3293_out0 ? v$_4444_out0 : v$_9345_out0;
assign v$_4427_out0 = { v$C2_125_out0,v$SEL1_15995_out0 };
assign v$_4458_out0 = { v$C2_156_out0,v$SEL1_16026_out0 };
assign v$_9328_out0 = { v$SEL1_9067_out0,v$C1_6263_out0 };
assign v$_9359_out0 = { v$SEL1_9098_out0,v$C1_6294_out0 };
assign v$ALUOUT_18679_out0 = v$MUX4_6214_out0;
assign v$ALUOUT_18680_out0 = v$MUX4_6215_out0;
assign v$MUX1_2564_out0 = v$LEFT$SHIT_3276_out0 ? v$_4427_out0 : v$_9328_out0;
assign v$MUX1_2595_out0 = v$LEFT$SHIT_3307_out0 ? v$_4458_out0 : v$_9359_out0;
assign v$ALUOUT_7203_out0 = v$ALUOUT_18679_out0;
assign v$ALUOUT_7204_out0 = v$ALUOUT_18680_out0;
assign v$MUX2_19185_out0 = v$EN_5427_out0 ? v$MUX1_2545_out0 : v$IN_4036_out0;
assign v$MUX2_19186_out0 = v$EN_5428_out0 ? v$MUX1_2550_out0 : v$IN_4037_out0;
assign v$MUX2_19191_out0 = v$EN_5433_out0 ? v$MUX1_2576_out0 : v$IN_4045_out0;
assign v$MUX2_19192_out0 = v$EN_5434_out0 ? v$MUX1_2581_out0 : v$IN_4046_out0;
assign v$MUX4_46_out0 = v$IR2$15_7754_out0 ? v$ALUOUT_7203_out0 : v$REGDIN_17124_out0;
assign v$MUX4_47_out0 = v$IR2$15_7755_out0 ? v$ALUOUT_7204_out0 : v$REGDIN_17125_out0;
assign v$MUX2_2696_out0 = v$EN_1501_out0 ? v$MUX1_2564_out0 : v$IN_5241_out0;
assign v$MUX2_2706_out0 = v$EN_1511_out0 ? v$MUX1_2595_out0 : v$IN_5251_out0;
assign v$OUT_15517_out0 = v$MUX2_19185_out0;
assign v$OUT_15522_out0 = v$MUX2_19186_out0;
assign v$OUT_15548_out0 = v$MUX2_19191_out0;
assign v$OUT_15553_out0 = v$MUX2_19192_out0;
assign v$ALUOUT_17162_out0 = v$ALUOUT_7203_out0;
assign v$ALUOUT_17163_out0 = v$ALUOUT_7204_out0;
assign v$IN_5369_out0 = v$OUT_15517_out0;
assign v$IN_5374_out0 = v$OUT_15522_out0;
assign v$IN_5400_out0 = v$OUT_15548_out0;
assign v$IN_5405_out0 = v$OUT_15553_out0;
assign v$ALUOUT_10671_out0 = v$ALUOUT_17162_out0;
assign v$ALUOUT_10672_out0 = v$ALUOUT_17163_out0;
assign v$OUT_15536_out0 = v$MUX2_2696_out0;
assign v$OUT_15567_out0 = v$MUX2_2706_out0;
assign v$IN_5385_out0 = v$OUT_15536_out0;
assign v$IN_5416_out0 = v$OUT_15567_out0;
assign v$_9123_out0 = v$ALUOUT_10671_out0[15:15];
assign v$_9124_out0 = v$ALUOUT_10672_out0[15:15];
assign v$IN_12352_out0 = v$IN_5369_out0;
assign v$IN_12353_out0 = v$IN_5374_out0;
assign v$IN_12358_out0 = v$IN_5400_out0;
assign v$IN_12359_out0 = v$IN_5405_out0;
assign v$EQ1_16882_out0 = v$ALUOUT_10671_out0 == 16'h0;
assign v$EQ1_16883_out0 = v$ALUOUT_10672_out0 == 16'h0;
assign v$IN_5240_out0 = v$IN_5385_out0;
assign v$IN_5250_out0 = v$IN_5416_out0;
assign v$SEL1_9050_out0 = v$IN_12352_out0[23:2];
assign v$SEL1_9055_out0 = v$IN_12353_out0[23:2];
assign v$SEL1_9081_out0 = v$IN_12358_out0[23:2];
assign v$SEL1_9086_out0 = v$IN_12359_out0[23:2];
assign v$G18_14176_out0 = v$_9123_out0 && v$IR2$VALID_13833_out0;
assign v$G18_14177_out0 = v$_9124_out0 && v$IR2$VALID_13834_out0;
assign v$G17_14419_out0 = v$EQ1_16882_out0 && v$IR2$VALID_13833_out0;
assign v$G17_14420_out0 = v$EQ1_16883_out0 && v$IR2$VALID_13834_out0;
assign v$SEL1_15978_out0 = v$IN_12352_out0[21:0];
assign v$SEL1_15983_out0 = v$IN_12353_out0[21:0];
assign v$SEL1_16009_out0 = v$IN_12358_out0[21:0];
assign v$SEL1_16014_out0 = v$IN_12359_out0[21:0];
assign v$MUX3_1579_out0 = v$G18_14176_out0 ? v$G18_14176_out0 : v$REG2_12370_out0;
assign v$MUX3_1580_out0 = v$G18_14177_out0 ? v$G18_14177_out0 : v$REG2_12371_out0;
assign v$_4410_out0 = { v$C2_108_out0,v$SEL1_15978_out0 };
assign v$_4415_out0 = { v$C2_113_out0,v$SEL1_15983_out0 };
assign v$_4441_out0 = { v$C2_139_out0,v$SEL1_16009_out0 };
assign v$_4446_out0 = { v$C2_144_out0,v$SEL1_16014_out0 };
assign v$SEL1_9066_out0 = v$IN_5240_out0[23:16];
assign v$SEL1_9097_out0 = v$IN_5250_out0[23:16];
assign v$_9311_out0 = { v$SEL1_9050_out0,v$C1_6246_out0 };
assign v$_9316_out0 = { v$SEL1_9055_out0,v$C1_6251_out0 };
assign v$_9342_out0 = { v$SEL1_9081_out0,v$C1_6277_out0 };
assign v$_9347_out0 = { v$SEL1_9086_out0,v$C1_6282_out0 };
assign v$MUX4_13221_out0 = v$G17_14419_out0 ? v$G17_14419_out0 : v$REG3_18364_out0;
assign v$MUX4_13222_out0 = v$G17_14420_out0 ? v$G17_14420_out0 : v$REG3_18365_out0;
assign v$SEL1_15994_out0 = v$IN_5240_out0[7:0];
assign v$SEL1_16025_out0 = v$IN_5250_out0[7:0];
assign v$MUX1_2547_out0 = v$LEFT$SHIT_3259_out0 ? v$_4410_out0 : v$_9311_out0;
assign v$MUX1_2552_out0 = v$LEFT$SHIT_3264_out0 ? v$_4415_out0 : v$_9316_out0;
assign v$MUX1_2578_out0 = v$LEFT$SHIT_3290_out0 ? v$_4441_out0 : v$_9342_out0;
assign v$MUX1_2583_out0 = v$LEFT$SHIT_3295_out0 ? v$_4446_out0 : v$_9347_out0;
assign v$EQ_3889_out0 = v$MUX4_13221_out0;
assign v$EQ_3890_out0 = v$MUX4_13222_out0;
assign v$_4426_out0 = { v$C2_124_out0,v$SEL1_15994_out0 };
assign v$_4457_out0 = { v$C2_155_out0,v$SEL1_16025_out0 };
assign v$_9327_out0 = { v$SEL1_9066_out0,v$C1_6262_out0 };
assign v$_9358_out0 = { v$SEL1_9097_out0,v$C1_6293_out0 };
assign v$MI_12694_out0 = v$MUX3_1579_out0;
assign v$MI_12695_out0 = v$MUX3_1580_out0;
assign v$EQ_450_out0 = v$EQ_3889_out0;
assign v$EQ_451_out0 = v$EQ_3890_out0;
assign v$MUX1_2563_out0 = v$LEFT$SHIT_3275_out0 ? v$_4426_out0 : v$_9327_out0;
assign v$MUX1_2594_out0 = v$LEFT$SHIT_3306_out0 ? v$_4457_out0 : v$_9358_out0;
assign v$MUX2_2670_out0 = v$EN_8199_out0 ? v$MUX1_2547_out0 : v$IN_12352_out0;
assign v$MUX2_2671_out0 = v$EN_8200_out0 ? v$MUX1_2552_out0 : v$IN_12353_out0;
assign v$MUX2_2676_out0 = v$EN_8205_out0 ? v$MUX1_2578_out0 : v$IN_12358_out0;
assign v$MUX2_2677_out0 = v$EN_8206_out0 ? v$MUX1_2583_out0 : v$IN_12359_out0;
assign v$MI_6504_out0 = v$MI_12694_out0;
assign v$MI_6505_out0 = v$MI_12695_out0;
assign v$MI_2609_out0 = v$MI_6504_out0;
assign v$MI_2610_out0 = v$MI_6505_out0;
assign v$MUX2_2695_out0 = v$EN_1500_out0 ? v$MUX1_2563_out0 : v$IN_5240_out0;
assign v$MUX2_2705_out0 = v$EN_1510_out0 ? v$MUX1_2594_out0 : v$IN_5250_out0;
assign v$EQ_6416_out0 = v$EQ_450_out0;
assign v$EQ_6417_out0 = v$EQ_451_out0;
assign v$OUT_15519_out0 = v$MUX2_2670_out0;
assign v$OUT_15524_out0 = v$MUX2_2671_out0;
assign v$OUT_15550_out0 = v$MUX2_2676_out0;
assign v$OUT_15555_out0 = v$MUX2_2677_out0;
assign v$EQ_3677_out0 = v$EQ_6416_out0;
assign v$EQ_3678_out0 = v$EQ_6417_out0;
assign v$IN_5368_out0 = v$OUT_15519_out0;
assign v$IN_5373_out0 = v$OUT_15524_out0;
assign v$IN_5399_out0 = v$OUT_15550_out0;
assign v$IN_5404_out0 = v$OUT_15555_out0;
assign v$MI_8756_out0 = v$MI_2609_out0;
assign v$MI_8757_out0 = v$MI_2610_out0;
assign v$OUT_15535_out0 = v$MUX2_2695_out0;
assign v$OUT_15566_out0 = v$MUX2_2705_out0;
assign v$MUX1_12194_out0 = v$G2_18057_out0 ? v$C1_4626_out0 : v$OUT_15535_out0;
assign v$MUX1_12198_out0 = v$G2_18061_out0 ? v$C1_4630_out0 : v$OUT_15566_out0;
assign v$MI_13060_out0 = v$MI_8756_out0;
assign v$MI_13061_out0 = v$MI_8757_out0;
assign v$EQ_14007_out0 = v$EQ_3677_out0;
assign v$EQ_14008_out0 = v$EQ_3678_out0;
assign v$IN_16196_out0 = v$IN_5368_out0;
assign v$IN_16197_out0 = v$IN_5373_out0;
assign v$IN_16202_out0 = v$IN_5399_out0;
assign v$IN_16203_out0 = v$IN_5404_out0;
assign v$SEL1_9049_out0 = v$IN_16196_out0[23:4];
assign v$SEL1_9054_out0 = v$IN_16197_out0[23:4];
assign v$SEL1_9080_out0 = v$IN_16202_out0[23:4];
assign v$SEL1_9085_out0 = v$IN_16203_out0[23:4];
assign v$OUT_10439_out0 = v$MUX1_12194_out0;
assign v$OUT_10443_out0 = v$MUX1_12198_out0;
assign v$MI_12451_out0 = v$MI_13060_out0;
assign v$MI_12452_out0 = v$MI_13061_out0;
assign v$EQ_15177_out0 = v$EQ_14007_out0;
assign v$EQ_15178_out0 = v$EQ_14008_out0;
assign v$SEL1_15977_out0 = v$IN_16196_out0[19:0];
assign v$SEL1_15982_out0 = v$IN_16197_out0[19:0];
assign v$SEL1_16008_out0 = v$IN_16202_out0[19:0];
assign v$SEL1_16013_out0 = v$IN_16203_out0[19:0];
assign v$G20_2788_out0 = v$G22_15929_out0 || v$EQ_15177_out0;
assign v$G20_2789_out0 = v$G22_15930_out0 || v$EQ_15178_out0;
assign v$OP2_4320_out0 = v$OUT_10439_out0;
assign v$OP2_4321_out0 = v$OUT_10443_out0;
assign v$_4409_out0 = { v$C2_107_out0,v$SEL1_15977_out0 };
assign v$_4414_out0 = { v$C2_112_out0,v$SEL1_15982_out0 };
assign v$_4440_out0 = { v$C2_138_out0,v$SEL1_16008_out0 };
assign v$_4445_out0 = { v$C2_143_out0,v$SEL1_16013_out0 };
assign v$_9310_out0 = { v$SEL1_9049_out0,v$C1_6245_out0 };
assign v$_9315_out0 = { v$SEL1_9054_out0,v$C1_6250_out0 };
assign v$_9341_out0 = { v$SEL1_9080_out0,v$C1_6276_out0 };
assign v$_9346_out0 = { v$SEL1_9085_out0,v$C1_6281_out0 };
assign v$G25_13323_out0 = v$JEQ_1833_out0 && v$EQ_15177_out0;
assign v$G25_13324_out0 = v$JEQ_1834_out0 && v$EQ_15178_out0;
assign v$G19_14605_out0 = v$JMI_13727_out0 && v$MI_12451_out0;
assign v$G19_14606_out0 = v$JMI_13728_out0 && v$MI_12452_out0;
assign v$G24_734_out0 = v$JLS_17065_out0 && v$G20_2788_out0;
assign v$G24_735_out0 = v$JLS_17066_out0 && v$G20_2789_out0;
assign v$MUX1_2546_out0 = v$LEFT$SHIT_3258_out0 ? v$_4409_out0 : v$_9310_out0;
assign v$MUX1_2551_out0 = v$LEFT$SHIT_3263_out0 ? v$_4414_out0 : v$_9315_out0;
assign v$MUX1_2577_out0 = v$LEFT$SHIT_3289_out0 ? v$_4440_out0 : v$_9341_out0;
assign v$MUX1_2582_out0 = v$LEFT$SHIT_3294_out0 ? v$_4445_out0 : v$_9346_out0;
assign v$B_14138_out0 = v$OP2_4320_out0;
assign v$B_14139_out0 = v$OP2_4321_out0;
assign v$G21_15897_out0 = v$G19_14605_out0 || v$G25_13323_out0;
assign v$G21_15898_out0 = v$G19_14606_out0 || v$G25_13324_out0;
assign v$B_80_out0 = v$B_14138_out0;
assign v$B_81_out0 = v$B_14139_out0;
assign v$G15_5719_out0 = v$JMP_4500_out0 || v$G21_15897_out0;
assign v$G15_5720_out0 = v$JMP_4501_out0 || v$G21_15898_out0;
assign v$MUX2_15817_out0 = v$EN_4963_out0 ? v$MUX1_2546_out0 : v$IN_16196_out0;
assign v$MUX2_15818_out0 = v$EN_4964_out0 ? v$MUX1_2551_out0 : v$IN_16197_out0;
assign v$MUX2_15823_out0 = v$EN_4969_out0 ? v$MUX1_2577_out0 : v$IN_16202_out0;
assign v$MUX2_15824_out0 = v$EN_4970_out0 ? v$MUX1_2582_out0 : v$IN_16203_out0;
assign v$MUX1_3094_out0 = v$START_4398_out0 ? v$B_80_out0 : v$B$SHIFTED_14379_out0;
assign v$MUX1_3095_out0 = v$START_4399_out0 ? v$B_81_out0 : v$B$SHIFTED_14380_out0;
assign v$MUX4_8416_out0 = v$START_4398_out0 ? v$B_80_out0 : v$B$SHIFTED_14379_out0;
assign v$MUX4_8417_out0 = v$START_4399_out0 ? v$B_81_out0 : v$B$SHIFTED_14380_out0;
assign v$OUT_15518_out0 = v$MUX2_15817_out0;
assign v$OUT_15523_out0 = v$MUX2_15818_out0;
assign v$OUT_15549_out0 = v$MUX2_15823_out0;
assign v$OUT_15554_out0 = v$MUX2_15824_out0;
assign v$G23_18289_out0 = v$G15_5719_out0 || v$G17_5699_out0;
assign v$G23_18290_out0 = v$G15_5720_out0 || v$G17_5700_out0;
assign v$G16_1476_out0 = v$G23_18289_out0 || v$G24_734_out0;
assign v$G16_1477_out0 = v$G23_18290_out0 || v$G24_735_out0;
assign v$IN_5366_out0 = v$OUT_15518_out0;
assign v$IN_5371_out0 = v$OUT_15523_out0;
assign v$IN_5395_out0 = v$MUX4_8416_out0;
assign v$IN_5397_out0 = v$OUT_15549_out0;
assign v$IN_5402_out0 = v$OUT_15554_out0;
assign v$IN_5426_out0 = v$MUX4_8417_out0;
assign v$OP2_13046_out0 = v$MUX1_3094_out0;
assign v$OP2_13047_out0 = v$MUX1_3095_out0;
assign v$SEL1_1437_out0 = v$OP2_13046_out0[0:0];
assign v$SEL1_1438_out0 = v$OP2_13047_out0[0:0];
assign v$IN_4044_out0 = v$IN_5395_out0;
assign v$IN_4053_out0 = v$IN_5426_out0;
assign v$IN_5234_out0 = v$IN_5366_out0;
assign v$IN_5236_out0 = v$IN_5371_out0;
assign v$IN_5244_out0 = v$IN_5397_out0;
assign v$IN_5246_out0 = v$IN_5402_out0;
assign v$TAKEJUMP_11294_out0 = v$G16_1476_out0;
assign v$TAKEJUMP_11295_out0 = v$G16_1477_out0;
assign v$SEL3_19268_out0 = v$OP2_13046_out0[0:0];
assign v$SEL3_19269_out0 = v$OP2_13047_out0[0:0];
assign v$SEL1_9047_out0 = v$IN_5234_out0[23:8];
assign v$SEL1_9052_out0 = v$IN_5236_out0[23:8];
assign v$SEL1_9076_out0 = v$IN_4044_out0[23:1];
assign v$SEL1_9078_out0 = v$IN_5244_out0[23:8];
assign v$SEL1_9083_out0 = v$IN_5246_out0[23:8];
assign v$SEL1_9107_out0 = v$IN_4053_out0[23:1];
assign v$MUX5_10765_out0 = v$SEL3_19268_out0 ? v$_1303_out0 : v$C4_18589_out0;
assign v$MUX5_10766_out0 = v$SEL3_19269_out0 ? v$_1304_out0 : v$C4_18590_out0;
assign v$MUX2_13050_out0 = v$SEL1_1437_out0 ? v$A_14857_out0 : v$C3_19045_out0;
assign v$MUX2_13051_out0 = v$SEL1_1438_out0 ? v$A_14858_out0 : v$C3_19046_out0;
assign v$G26_14220_out0 = v$G29_8174_out0 || v$TAKEJUMP_11294_out0;
assign v$G26_14221_out0 = v$G29_8175_out0 || v$TAKEJUMP_11295_out0;
assign v$SEL1_15975_out0 = v$IN_5234_out0[15:0];
assign v$SEL1_15980_out0 = v$IN_5236_out0[15:0];
assign v$SEL1_16004_out0 = v$IN_4044_out0[22:0];
assign v$SEL1_16006_out0 = v$IN_5244_out0[15:0];
assign v$SEL1_16011_out0 = v$IN_5246_out0[15:0];
assign v$SEL1_16035_out0 = v$IN_4053_out0[22:0];
assign v$_4407_out0 = { v$C2_105_out0,v$SEL1_15975_out0 };
assign v$_4412_out0 = { v$C2_110_out0,v$SEL1_15980_out0 };
assign v$_4436_out0 = { v$C2_134_out0,v$SEL1_16004_out0 };
assign v$_4438_out0 = { v$C2_136_out0,v$SEL1_16006_out0 };
assign v$_4443_out0 = { v$C2_141_out0,v$SEL1_16011_out0 };
assign v$_4467_out0 = { v$C2_165_out0,v$SEL1_16035_out0 };
assign v$B2_8722_out0 = v$MUX2_13050_out0;
assign v$B2_8725_out0 = v$MUX2_13051_out0;
assign v$_9308_out0 = { v$SEL1_9047_out0,v$C1_6243_out0 };
assign v$_9313_out0 = { v$SEL1_9052_out0,v$C1_6248_out0 };
assign v$_9337_out0 = { v$SEL1_9076_out0,v$C1_6272_out0 };
assign v$_9339_out0 = { v$SEL1_9078_out0,v$C1_6274_out0 };
assign v$_9344_out0 = { v$SEL1_9083_out0,v$C1_6279_out0 };
assign v$_9368_out0 = { v$SEL1_9107_out0,v$C1_6303_out0 };
assign v$MUX8_12853_out0 = v$G26_14220_out0 ? v$MUX5_17586_out0 : v$PCINTERRUPT_18413_out0;
assign v$MUX8_12854_out0 = v$G26_14221_out0 ? v$MUX5_17587_out0 : v$PCINTERRUPT_18414_out0;
assign v$MUX3_18515_out0 = v$START_4398_out0 ? v$MUX5_10765_out0 : v$RESULT_5279_out0;
assign v$MUX3_18516_out0 = v$START_4399_out0 ? v$MUX5_10766_out0 : v$RESULT_5280_out0;
assign v$MUX1_2544_out0 = v$LEFT$SHIT_3256_out0 ? v$_4407_out0 : v$_9308_out0;
assign v$MUX1_2549_out0 = v$LEFT$SHIT_3261_out0 ? v$_4412_out0 : v$_9313_out0;
assign v$MUX1_2573_out0 = v$LEFT$SHIT_3285_out0 ? v$_4436_out0 : v$_9337_out0;
assign v$MUX1_2575_out0 = v$LEFT$SHIT_3287_out0 ? v$_4438_out0 : v$_9339_out0;
assign v$MUX1_2580_out0 = v$LEFT$SHIT_3292_out0 ? v$_4443_out0 : v$_9344_out0;
assign v$MUX1_2604_out0 = v$LEFT$SHIT_3316_out0 ? v$_4467_out0 : v$_9368_out0;
assign v$MUX2_3903_out0 = v$ININTERRUPT_1277_out0 ? v$MUX8_12853_out0 : v$PCNORMAL_13337_out0;
assign v$MUX2_3904_out0 = v$ININTERRUPT_1278_out0 ? v$MUX8_12854_out0 : v$PCNORMAL_13338_out0;
assign v$_4142_out0 = v$B2_8722_out0[11:0];
assign v$_4142_out1 = v$B2_8722_out0[23:12];
assign v$_4145_out0 = v$B2_8725_out0[11:0];
assign v$_4145_out1 = v$B2_8725_out0[23:12];
assign v$A1_14172_out0 = v$MUX3_18515_out0;
assign v$A1_14175_out0 = v$MUX3_18516_out0;
assign v$_1371_out0 = v$_4142_out1[5:0];
assign v$_1371_out1 = v$_4142_out1[11:6];
assign v$_1374_out0 = v$_4145_out1[5:0];
assign v$_1374_out1 = v$_4145_out1[11:6];
assign v$_1679_out0 = v$_4142_out0[5:0];
assign v$_1679_out1 = v$_4142_out0[11:6];
assign v$_1682_out0 = v$_4145_out0[5:0];
assign v$_1682_out1 = v$_4145_out0[11:6];
assign v$MUX4_1731_out0 = v$TAKEJUMP_11294_out0 ? v$N_18899_out0 : v$MUX2_3903_out0;
assign v$MUX4_1732_out0 = v$TAKEJUMP_11295_out0 ? v$N_18900_out0 : v$MUX2_3904_out0;
assign v$MUX2_2689_out0 = v$EN_1494_out0 ? v$MUX1_2544_out0 : v$IN_5234_out0;
assign v$MUX2_2691_out0 = v$EN_1496_out0 ? v$MUX1_2549_out0 : v$IN_5236_out0;
assign v$MUX2_2699_out0 = v$EN_1504_out0 ? v$MUX1_2575_out0 : v$IN_5244_out0;
assign v$MUX2_2701_out0 = v$EN_1506_out0 ? v$MUX1_2580_out0 : v$IN_5246_out0;
assign v$_7862_out0 = v$A1_14172_out0[11:0];
assign v$_7862_out1 = v$A1_14172_out0[23:12];
assign v$_7865_out0 = v$A1_14175_out0[11:0];
assign v$_7865_out1 = v$A1_14175_out0[23:12];
assign v$MUX2_15436_out0 = v$EN_4056_out0 ? v$MUX1_2573_out0 : v$IN_4044_out0;
assign v$MUX2_15439_out0 = v$EN_4059_out0 ? v$MUX1_2604_out0 : v$IN_4053_out0;
assign v$PC_3365_out0 = v$MUX4_1731_out0;
assign v$PC_3366_out0 = v$MUX4_1732_out0;
assign v$_10358_out0 = v$_1371_out1[2:0];
assign v$_10358_out1 = v$_1371_out1[5:3];
assign v$_10361_out0 = v$_1374_out1[2:0];
assign v$_10361_out1 = v$_1374_out1[5:3];
assign v$_13563_out0 = v$_1679_out1[2:0];
assign v$_13563_out1 = v$_1679_out1[5:3];
assign v$_13566_out0 = v$_1682_out1[2:0];
assign v$_13566_out1 = v$_1682_out1[5:3];
assign v$_14326_out0 = v$_1679_out0[2:0];
assign v$_14326_out1 = v$_1679_out0[5:3];
assign v$_14329_out0 = v$_1682_out0[2:0];
assign v$_14329_out1 = v$_1682_out0[5:3];
assign v$OUT_15516_out0 = v$MUX2_2689_out0;
assign v$OUT_15521_out0 = v$MUX2_2691_out0;
assign v$OUT_15545_out0 = v$MUX2_15436_out0;
assign v$OUT_15547_out0 = v$MUX2_2699_out0;
assign v$OUT_15552_out0 = v$MUX2_2701_out0;
assign v$OUT_15576_out0 = v$MUX2_15439_out0;
assign v$_16725_out0 = v$_7862_out0[5:0];
assign v$_16725_out1 = v$_7862_out0[11:6];
assign v$_16728_out0 = v$_7865_out0[5:0];
assign v$_16728_out1 = v$_7865_out0[11:6];
assign v$_17624_out0 = v$_7862_out1[5:0];
assign v$_17624_out1 = v$_7862_out1[11:6];
assign v$_17627_out0 = v$_7865_out1[5:0];
assign v$_17627_out1 = v$_7865_out1[11:6];
assign v$_18342_out0 = v$_1371_out0[2:0];
assign v$_18342_out1 = v$_1371_out0[5:3];
assign v$_18345_out0 = v$_1374_out0[2:0];
assign v$_18345_out1 = v$_1374_out0[5:3];
assign v$NEXTINSTRUCTIONADDRESS_19015_out0 = v$MUX4_1731_out0;
assign v$NEXTINSTRUCTIONADDRESS_19016_out0 = v$MUX4_1732_out0;
assign v$_2026_out0 = v$_17624_out1[2:0];
assign v$_2026_out1 = v$_17624_out1[5:3];
assign v$_2029_out0 = v$_17627_out1[2:0];
assign v$_2029_out1 = v$_17627_out1[5:3];
assign v$_3131_out0 = v$_14326_out0[0:0];
assign v$_3131_out1 = v$_14326_out0[2:2];
assign v$_3134_out0 = v$_14329_out0[0:0];
assign v$_3134_out1 = v$_14329_out0[2:2];
assign v$IN_5365_out0 = v$OUT_15516_out0;
assign v$IN_5370_out0 = v$OUT_15521_out0;
assign v$IN_5396_out0 = v$OUT_15547_out0;
assign v$IN_5401_out0 = v$OUT_15552_out0;
assign v$PCNEXT_6889_out0 = v$NEXTINSTRUCTIONADDRESS_19015_out0;
assign v$PCNEXT_6890_out0 = v$NEXTINSTRUCTIONADDRESS_19016_out0;
assign v$_8090_out0 = v$_18342_out0[0:0];
assign v$_8090_out1 = v$_18342_out0[2:2];
assign v$_8093_out0 = v$_18345_out0[0:0];
assign v$_8093_out1 = v$_18345_out0[2:2];
assign v$_9391_out0 = v$_10358_out1[0:0];
assign v$_9391_out1 = v$_10358_out1[2:2];
assign v$_9394_out0 = v$_10361_out1[0:0];
assign v$_9394_out1 = v$_10361_out1[2:2];
assign v$_10476_out0 = v$_17624_out0[2:0];
assign v$_10476_out1 = v$_17624_out0[5:3];
assign v$_10479_out0 = v$_17627_out0[2:0];
assign v$_10479_out1 = v$_17627_out0[5:3];
assign v$_11266_out0 = v$_13563_out1[0:0];
assign v$_11266_out1 = v$_13563_out1[2:2];
assign v$_11269_out0 = v$_13566_out1[0:0];
assign v$_11269_out1 = v$_13566_out1[2:2];
assign v$_14357_out0 = v$_16725_out0[2:0];
assign v$_14357_out1 = v$_16725_out0[5:3];
assign v$_14360_out0 = v$_16728_out0[2:0];
assign v$_14360_out1 = v$_16728_out0[5:3];
assign {v$A1_15427_out1,v$A1_15427_out0 } = v$PC_3365_out0 + v$C1_16546_out0 + v$EN_9408_out0;
assign {v$A1_15428_out1,v$A1_15428_out0 } = v$PC_3366_out0 + v$C1_16547_out0 + v$EN_9409_out0;
assign v$_15760_out0 = v$_10358_out0[0:0];
assign v$_15760_out1 = v$_10358_out0[2:2];
assign v$_15763_out0 = v$_10361_out0[0:0];
assign v$_15763_out1 = v$_10361_out0[2:2];
assign v$_16878_out0 = v$_18342_out1[0:0];
assign v$_16878_out1 = v$_18342_out1[2:2];
assign v$_16881_out0 = v$_18345_out1[0:0];
assign v$_16881_out1 = v$_18345_out1[2:2];
assign v$_17363_out0 = v$_14326_out1[0:0];
assign v$_17363_out1 = v$_14326_out1[2:2];
assign v$_17366_out0 = v$_14329_out1[0:0];
assign v$_17366_out1 = v$_14329_out1[2:2];
assign v$_18789_out0 = v$_13563_out0[0:0];
assign v$_18789_out1 = v$_13563_out0[2:2];
assign v$_18792_out0 = v$_13566_out0[0:0];
assign v$_18792_out1 = v$_13566_out0[2:2];
assign v$_19029_out0 = v$_16725_out1[2:0];
assign v$_19029_out1 = v$_16725_out1[5:3];
assign v$_19032_out0 = v$_16728_out1[2:0];
assign v$_19032_out1 = v$_16728_out1[5:3];
assign v$_1464_out0 = v$_19029_out0[0:0];
assign v$_1464_out1 = v$_19029_out0[2:2];
assign v$_1467_out0 = v$_19032_out0[0:0];
assign v$_1467_out1 = v$_19032_out0[2:2];
assign v$_1517_out0 = v$_14357_out1[0:0];
assign v$_1517_out1 = v$_14357_out1[2:2];
assign v$_1520_out0 = v$_14360_out1[0:0];
assign v$_1520_out1 = v$_14360_out1[2:2];
assign v$_2016_out0 = v$_2026_out1[0:0];
assign v$_2016_out1 = v$_2026_out1[2:2];
assign v$_2019_out0 = v$_2029_out1[0:0];
assign v$_2019_out1 = v$_2029_out1[2:2];
assign v$PC$NEXT0_2098_out0 = v$PCNEXT_6890_out0;
assign v$B12_2116_out0 = v$_8090_out0;
assign v$B12_2119_out0 = v$_8093_out0;
assign v$B0_3423_out0 = v$_3131_out0;
assign v$B0_3426_out0 = v$_3134_out0;
assign v$PC$NEXT1_3697_out0 = v$PCNEXT_6889_out0;
assign v$B9_4222_out0 = v$_11266_out0;
assign v$B9_4225_out0 = v$_11269_out0;
assign v$IN_5233_out0 = v$IN_5365_out0;
assign v$IN_5235_out0 = v$IN_5370_out0;
assign v$IN_5243_out0 = v$IN_5396_out0;
assign v$IN_5245_out0 = v$IN_5401_out0;
assign v$IGNORE_5650_out0 = v$A1_15427_out1;
assign v$IGNORE_5651_out0 = v$A1_15428_out1;
assign v$_7178_out0 = v$_18789_out1[0:0];
assign v$_7178_out1 = v$_18789_out1[1:1];
assign v$_7181_out0 = v$_18792_out1[0:0];
assign v$_7181_out1 = v$_18792_out1[1:1];
assign v$_7260_out0 = v$_17363_out1[0:0];
assign v$_7260_out1 = v$_17363_out1[1:1];
assign v$_7263_out0 = v$_17366_out1[0:0];
assign v$_7263_out1 = v$_17366_out1[1:1];
assign v$_7357_out0 = v$_14357_out0[0:0];
assign v$_7357_out1 = v$_14357_out0[2:2];
assign v$_7360_out0 = v$_14360_out0[0:0];
assign v$_7360_out1 = v$_14360_out0[2:2];
assign v$_9755_out0 = v$_9391_out1[0:0];
assign v$_9755_out1 = v$_9391_out1[1:1];
assign v$_9758_out0 = v$_9394_out1[0:0];
assign v$_9758_out1 = v$_9394_out1[1:1];
assign v$B3_9847_out0 = v$_17363_out0;
assign v$B3_9850_out0 = v$_17366_out0;
assign v$_9875_out0 = v$_11266_out1[0:0];
assign v$_9875_out1 = v$_11266_out1[1:1];
assign v$_9878_out0 = v$_11269_out1[0:0];
assign v$_9878_out1 = v$_11269_out1[1:1];
assign v$B15_10448_out0 = v$_16878_out0;
assign v$B15_10451_out0 = v$_16881_out0;
assign v$_10900_out0 = v$_10476_out0[0:0];
assign v$_10900_out1 = v$_10476_out0[2:2];
assign v$_10903_out0 = v$_10479_out0[0:0];
assign v$_10903_out1 = v$_10479_out0[2:2];
assign v$B18_11370_out0 = v$_15760_out0;
assign v$B18_11373_out0 = v$_15763_out0;
assign v$_11415_out0 = v$_19029_out1[0:0];
assign v$_11415_out1 = v$_19029_out1[2:2];
assign v$_11418_out0 = v$_19032_out1[0:0];
assign v$_11418_out1 = v$_19032_out1[2:2];
assign v$_11533_out0 = v$_3131_out1[0:0];
assign v$_11533_out1 = v$_3131_out1[1:1];
assign v$_11536_out0 = v$_3134_out1[0:0];
assign v$_11536_out1 = v$_3134_out1[1:1];
assign v$_11598_out0 = v$_2026_out0[0:0];
assign v$_11598_out1 = v$_2026_out0[2:2];
assign v$_11601_out0 = v$_2029_out0[0:0];
assign v$_11601_out1 = v$_2029_out0[2:2];
assign v$_13760_out0 = v$_16878_out1[0:0];
assign v$_13760_out1 = v$_16878_out1[1:1];
assign v$_13763_out0 = v$_16881_out1[0:0];
assign v$_13763_out1 = v$_16881_out1[1:1];
assign v$B6_13885_out0 = v$_18789_out0;
assign v$B6_13888_out0 = v$_18792_out0;
assign v$SUM_14246_out0 = v$A1_15427_out0;
assign v$SUM_14247_out0 = v$A1_15428_out0;
assign v$_16744_out0 = v$_10476_out1[0:0];
assign v$_16744_out1 = v$_10476_out1[2:2];
assign v$_16747_out0 = v$_10479_out1[0:0];
assign v$_16747_out1 = v$_10479_out1[2:2];
assign v$_17210_out0 = v$_15760_out1[0:0];
assign v$_17210_out1 = v$_15760_out1[1:1];
assign v$_17213_out0 = v$_15763_out1[0:0];
assign v$_17213_out1 = v$_15763_out1[1:1];
assign v$_17967_out0 = v$_8090_out1[0:0];
assign v$_17967_out1 = v$_8090_out1[1:1];
assign v$_17970_out0 = v$_8093_out1[0:0];
assign v$_17970_out1 = v$_8093_out1[1:1];
assign v$B21_18691_out0 = v$_9391_out0;
assign v$B21_18694_out0 = v$_9394_out0;
assign v$A6_322_out0 = v$_1464_out0;
assign v$A6_325_out0 = v$_1467_out0;
assign v$B23_1443_out0 = v$_9755_out1;
assign v$B23_1446_out0 = v$_9758_out1;
assign v$A21_2794_out0 = v$_2016_out0;
assign v$A21_2797_out0 = v$_2019_out0;
assign v$ADDRESS_2829_out0 = v$PC$NEXT1_3697_out0;
assign v$B_2944_out0 = v$B6_13885_out0;
assign v$B_2945_out0 = v$B3_9847_out0;
assign v$B_2946_out0 = v$B21_18691_out0;
assign v$B_2947_out0 = v$B9_4222_out0;
assign v$B_2948_out0 = v$B15_10448_out0;
assign v$B_2952_out0 = v$B12_2116_out0;
assign v$B_2956_out0 = v$B0_3423_out0;
assign v$B_2961_out0 = v$B18_11370_out0;
assign v$B_3016_out0 = v$B6_13888_out0;
assign v$B_3017_out0 = v$B3_9850_out0;
assign v$B_3018_out0 = v$B21_18694_out0;
assign v$B_3019_out0 = v$B9_4225_out0;
assign v$B_3020_out0 = v$B15_10451_out0;
assign v$B_3024_out0 = v$B12_2119_out0;
assign v$B_3028_out0 = v$B0_3426_out0;
assign v$B_3033_out0 = v$B18_11373_out0;
assign v$B2_3328_out0 = v$_11533_out1;
assign v$B2_3331_out0 = v$_11536_out1;
assign v$A12_3357_out0 = v$_10900_out0;
assign v$A12_3360_out0 = v$_10903_out0;
assign v$A9_3645_out0 = v$_11415_out0;
assign v$A9_3648_out0 = v$_11418_out0;
assign v$B20_4114_out0 = v$_17210_out1;
assign v$B20_4117_out0 = v$_17213_out1;
assign v$B14_4160_out0 = v$_17967_out1;
assign v$B14_4163_out0 = v$_17970_out1;
assign v$A0_4470_out0 = v$_7357_out0;
assign v$A0_4473_out0 = v$_7360_out0;
assign v$_6230_out0 = v$_16744_out1[0:0];
assign v$_6230_out1 = v$_16744_out1[1:1];
assign v$_6233_out0 = v$_16747_out1[0:0];
assign v$_6233_out1 = v$_16747_out1[1:1];
assign v$_7678_out0 = v$_1517_out1[0:0];
assign v$_7678_out1 = v$_1517_out1[1:1];
assign v$_7681_out0 = v$_1520_out1[0:0];
assign v$_7681_out1 = v$_1520_out1[1:1];
assign v$PC0_8220_out0 = v$PC$NEXT0_2098_out0;
assign v$B1_8428_out0 = v$_11533_out0;
assign v$B1_8431_out0 = v$_11536_out0;
assign v$B13_9024_out0 = v$_17967_out0;
assign v$B13_9027_out0 = v$_17970_out0;
assign v$SEL1_9046_out0 = v$IN_5233_out0[23:16];
assign v$SEL1_9051_out0 = v$IN_5235_out0[23:16];
assign v$SEL1_9077_out0 = v$IN_5243_out0[23:16];
assign v$SEL1_9082_out0 = v$IN_5245_out0[23:16];
assign v$B11_9445_out0 = v$_9875_out1;
assign v$B11_9448_out0 = v$_9878_out1;
assign v$B10_10299_out0 = v$_9875_out0;
assign v$B10_10302_out0 = v$_9878_out0;
assign v$_10741_out0 = v$_2016_out1[0:0];
assign v$_10741_out1 = v$_2016_out1[1:1];
assign v$_10744_out0 = v$_2019_out1[0:0];
assign v$_10744_out1 = v$_2019_out1[1:1];
assign v$B22_11302_out0 = v$_9755_out0;
assign v$B22_11305_out0 = v$_9758_out0;
assign v$_12180_out0 = v$_7357_out1[0:0];
assign v$_12180_out1 = v$_7357_out1[1:1];
assign v$_12183_out0 = v$_7360_out1[0:0];
assign v$_12183_out1 = v$_7360_out1[1:1];
assign v$PC1_12778_out0 = v$PC$NEXT1_3697_out0;
assign v$B8_13717_out0 = v$_7178_out1;
assign v$B8_13720_out0 = v$_7181_out1;
assign v$A3_15211_out0 = v$_1517_out0;
assign v$A3_15214_out0 = v$_1520_out0;
assign v$B4_15268_out0 = v$_7260_out0;
assign v$B4_15271_out0 = v$_7263_out0;
assign v$ADDRESS_15794_out0 = v$PC$NEXT0_2098_out0;
assign v$SEL1_15974_out0 = v$IN_5233_out0[7:0];
assign v$SEL1_15979_out0 = v$IN_5235_out0[7:0];
assign v$SEL1_16005_out0 = v$IN_5243_out0[7:0];
assign v$SEL1_16010_out0 = v$IN_5245_out0[7:0];
assign v$B17_16127_out0 = v$_13760_out1;
assign v$B17_16130_out0 = v$_13763_out1;
assign v$_16341_out0 = v$_1464_out1[0:0];
assign v$_16341_out1 = v$_1464_out1[1:1];
assign v$_16344_out0 = v$_1467_out1[0:0];
assign v$_16344_out1 = v$_1467_out1[1:1];
assign v$_16793_out0 = v$_10900_out1[0:0];
assign v$_16793_out1 = v$_10900_out1[1:1];
assign v$_16796_out0 = v$_10903_out1[0:0];
assign v$_16796_out1 = v$_10903_out1[1:1];
assign v$B16_17036_out0 = v$_13760_out0;
assign v$B16_17039_out0 = v$_13763_out0;
assign v$_17324_out0 = v$_11598_out1[0:0];
assign v$_17324_out1 = v$_11598_out1[1:1];
assign v$_17327_out0 = v$_11601_out1[0:0];
assign v$_17327_out1 = v$_11601_out1[1:1];
assign v$B19_17412_out0 = v$_17210_out0;
assign v$B19_17415_out0 = v$_17213_out0;
assign v$B7_17636_out0 = v$_7178_out0;
assign v$B7_17639_out0 = v$_7181_out0;
assign v$A15_17959_out0 = v$_16744_out0;
assign v$A15_17962_out0 = v$_16747_out0;
assign v$A18_18302_out0 = v$_11598_out0;
assign v$A18_18305_out0 = v$_11601_out0;
assign v$_18368_out0 = v$_11415_out1[0:0];
assign v$_18368_out1 = v$_11415_out1[1:1];
assign v$_18371_out0 = v$_11418_out1[0:0];
assign v$_18371_out1 = v$_11418_out1[1:1];
assign v$B5_18980_out0 = v$_7260_out1;
assign v$B5_18983_out0 = v$_7263_out1;
assign v$A14_740_out0 = v$_16793_out1;
assign v$A14_743_out0 = v$_16796_out1;
assign v$A19_1365_out0 = v$_17324_out0;
assign v$A19_1368_out0 = v$_17327_out0;
assign v$A10_1705_out0 = v$_18368_out0;
assign v$A10_1708_out0 = v$_18371_out0;
assign v$A1_1871_out0 = v$_12180_out0;
assign v$A1_1874_out0 = v$_12183_out0;
assign v$_2613_out0 = v$ADDRESS_15794_out0[9:0];
assign v$_2613_out1 = v$ADDRESS_15794_out0[11:2];
assign v$_2810_out0 = v$ADDRESS_2829_out0[9:0];
assign v$_2810_out1 = v$ADDRESS_2829_out0[11:2];
assign v$B_2949_out0 = v$B7_17636_out0;
assign v$B_2950_out0 = v$B1_8428_out0;
assign v$B_2951_out0 = v$B14_4160_out0;
assign v$B_2953_out0 = v$B8_13717_out0;
assign v$B_2954_out0 = v$B17_16127_out0;
assign v$B_2955_out0 = v$B23_1443_out0;
assign v$B_2957_out0 = v$B13_9024_out0;
assign v$B_2958_out0 = v$B4_15268_out0;
assign v$B_2959_out0 = v$B19_17412_out0;
assign v$B_2960_out0 = v$B22_11302_out0;
assign v$B_2962_out0 = v$B10_10299_out0;
assign v$B_2963_out0 = v$B20_4114_out0;
assign v$B_2964_out0 = v$B2_3328_out0;
assign v$B_2965_out0 = v$B11_9445_out0;
assign v$B_2966_out0 = v$B5_18980_out0;
assign v$B_2967_out0 = v$B16_17036_out0;
assign v$B_3021_out0 = v$B7_17639_out0;
assign v$B_3022_out0 = v$B1_8431_out0;
assign v$B_3023_out0 = v$B14_4163_out0;
assign v$B_3025_out0 = v$B8_13720_out0;
assign v$B_3026_out0 = v$B17_16130_out0;
assign v$B_3027_out0 = v$B23_1446_out0;
assign v$B_3029_out0 = v$B13_9027_out0;
assign v$B_3030_out0 = v$B4_15271_out0;
assign v$B_3031_out0 = v$B19_17415_out0;
assign v$B_3032_out0 = v$B22_11305_out0;
assign v$B_3034_out0 = v$B10_10302_out0;
assign v$B_3035_out0 = v$B20_4117_out0;
assign v$B_3036_out0 = v$B2_3331_out0;
assign v$B_3037_out0 = v$B11_9448_out0;
assign v$B_3038_out0 = v$B5_18983_out0;
assign v$B_3039_out0 = v$B16_17039_out0;
assign v$_4406_out0 = { v$C2_104_out0,v$SEL1_15974_out0 };
assign v$_4411_out0 = { v$C2_109_out0,v$SEL1_15979_out0 };
assign v$_4437_out0 = { v$C2_135_out0,v$SEL1_16005_out0 };
assign v$_4442_out0 = { v$C2_140_out0,v$SEL1_16010_out0 };
assign v$A22_4592_out0 = v$_10741_out0;
assign v$A22_4595_out0 = v$_10744_out0;
assign v$A20_4605_out0 = v$_17324_out1;
assign v$A20_4608_out0 = v$_17327_out1;
assign v$A23_5283_out0 = v$_10741_out1;
assign v$A23_5286_out0 = v$_10744_out1;
assign v$A5_6903_out0 = v$_7678_out1;
assign v$A5_6906_out0 = v$_7681_out1;
assign v$A_7439_out0 = v$A6_322_out0;
assign v$A_7440_out0 = v$A3_15211_out0;
assign v$A_7441_out0 = v$A21_2794_out0;
assign v$A_7442_out0 = v$A9_3645_out0;
assign v$A_7443_out0 = v$A15_17959_out0;
assign v$A_7447_out0 = v$A12_3357_out0;
assign v$A_7451_out0 = v$A0_4470_out0;
assign v$A_7456_out0 = v$A18_18302_out0;
assign v$A_7511_out0 = v$A6_325_out0;
assign v$A_7512_out0 = v$A3_15214_out0;
assign v$A_7513_out0 = v$A21_2797_out0;
assign v$A_7514_out0 = v$A9_3648_out0;
assign v$A_7515_out0 = v$A15_17962_out0;
assign v$A_7519_out0 = v$A12_3360_out0;
assign v$A_7523_out0 = v$A0_4473_out0;
assign v$A_7528_out0 = v$A18_18305_out0;
assign v$_9307_out0 = { v$SEL1_9046_out0,v$C1_6242_out0 };
assign v$_9312_out0 = { v$SEL1_9051_out0,v$C1_6247_out0 };
assign v$_9338_out0 = { v$SEL1_9077_out0,v$C1_6273_out0 };
assign v$_9343_out0 = { v$SEL1_9082_out0,v$C1_6278_out0 };
assign v$A11_10388_out0 = v$_18368_out1;
assign v$A11_10391_out0 = v$_18371_out1;
assign {v$A1A_12226_out1,v$A1A_12226_out0 } = v$A0_4470_out0 + v$B0_3423_out0 + v$C1_4635_out0;
assign {v$A1A_12229_out1,v$A1A_12229_out0 } = v$A0_4473_out0 + v$B0_3426_out0 + v$C1_4638_out0;
assign v$A16_14193_out0 = v$_6230_out0;
assign v$A16_14196_out0 = v$_6233_out0;
assign v$A13_14447_out0 = v$_16793_out0;
assign v$A13_14450_out0 = v$_16796_out0;
assign v$A7_15893_out0 = v$_16341_out0;
assign v$A7_15896_out0 = v$_16344_out0;
assign v$A17_17344_out0 = v$_6230_out1;
assign v$A17_17347_out0 = v$_6233_out1;
assign v$A4_18140_out0 = v$_7678_out0;
assign v$A4_18143_out0 = v$_7681_out0;
assign v$A8_18699_out0 = v$_16341_out1;
assign v$A8_18702_out0 = v$_16344_out1;
assign v$A2_18870_out0 = v$_12180_out1;
assign v$A2_18873_out0 = v$_12183_out1;
assign v$MUX1_2543_out0 = v$LEFT$SHIT_3255_out0 ? v$_4406_out0 : v$_9307_out0;
assign v$MUX1_2548_out0 = v$LEFT$SHIT_3260_out0 ? v$_4411_out0 : v$_9312_out0;
assign v$MUX1_2574_out0 = v$LEFT$SHIT_3286_out0 ? v$_4437_out0 : v$_9338_out0;
assign v$MUX1_2579_out0 = v$LEFT$SHIT_3291_out0 ? v$_4442_out0 : v$_9343_out0;
assign v$G2_5526_out0 = ((v$A_7439_out0 && !v$B_2944_out0) || (!v$A_7439_out0) && v$B_2944_out0);
assign v$G2_5527_out0 = ((v$A_7440_out0 && !v$B_2945_out0) || (!v$A_7440_out0) && v$B_2945_out0);
assign v$G2_5528_out0 = ((v$A_7441_out0 && !v$B_2946_out0) || (!v$A_7441_out0) && v$B_2946_out0);
assign v$G2_5529_out0 = ((v$A_7442_out0 && !v$B_2947_out0) || (!v$A_7442_out0) && v$B_2947_out0);
assign v$G2_5530_out0 = ((v$A_7443_out0 && !v$B_2948_out0) || (!v$A_7443_out0) && v$B_2948_out0);
assign v$G2_5534_out0 = ((v$A_7447_out0 && !v$B_2952_out0) || (!v$A_7447_out0) && v$B_2952_out0);
assign v$G2_5538_out0 = ((v$A_7451_out0 && !v$B_2956_out0) || (!v$A_7451_out0) && v$B_2956_out0);
assign v$G2_5543_out0 = ((v$A_7456_out0 && !v$B_2961_out0) || (!v$A_7456_out0) && v$B_2961_out0);
assign v$G2_5598_out0 = ((v$A_7511_out0 && !v$B_3016_out0) || (!v$A_7511_out0) && v$B_3016_out0);
assign v$G2_5599_out0 = ((v$A_7512_out0 && !v$B_3017_out0) || (!v$A_7512_out0) && v$B_3017_out0);
assign v$G2_5600_out0 = ((v$A_7513_out0 && !v$B_3018_out0) || (!v$A_7513_out0) && v$B_3018_out0);
assign v$G2_5601_out0 = ((v$A_7514_out0 && !v$B_3019_out0) || (!v$A_7514_out0) && v$B_3019_out0);
assign v$G2_5602_out0 = ((v$A_7515_out0 && !v$B_3020_out0) || (!v$A_7515_out0) && v$B_3020_out0);
assign v$G2_5606_out0 = ((v$A_7519_out0 && !v$B_3024_out0) || (!v$A_7519_out0) && v$B_3024_out0);
assign v$G2_5610_out0 = ((v$A_7523_out0 && !v$B_3028_out0) || (!v$A_7523_out0) && v$B_3028_out0);
assign v$G2_5615_out0 = ((v$A_7528_out0 && !v$B_3033_out0) || (!v$A_7528_out0) && v$B_3033_out0);
assign v$A_7444_out0 = v$A7_15893_out0;
assign v$A_7445_out0 = v$A1_1871_out0;
assign v$A_7446_out0 = v$A14_740_out0;
assign v$A_7448_out0 = v$A8_18699_out0;
assign v$A_7449_out0 = v$A17_17344_out0;
assign v$A_7450_out0 = v$A23_5283_out0;
assign v$A_7452_out0 = v$A13_14447_out0;
assign v$A_7453_out0 = v$A4_18140_out0;
assign v$A_7454_out0 = v$A19_1365_out0;
assign v$A_7455_out0 = v$A22_4592_out0;
assign v$A_7457_out0 = v$A10_1705_out0;
assign v$A_7458_out0 = v$A20_4605_out0;
assign v$A_7459_out0 = v$A2_18870_out0;
assign v$A_7460_out0 = v$A11_10388_out0;
assign v$A_7461_out0 = v$A5_6903_out0;
assign v$A_7462_out0 = v$A16_14193_out0;
assign v$A_7516_out0 = v$A7_15896_out0;
assign v$A_7517_out0 = v$A1_1874_out0;
assign v$A_7518_out0 = v$A14_743_out0;
assign v$A_7520_out0 = v$A8_18702_out0;
assign v$A_7521_out0 = v$A17_17347_out0;
assign v$A_7522_out0 = v$A23_5286_out0;
assign v$A_7524_out0 = v$A13_14450_out0;
assign v$A_7525_out0 = v$A4_18143_out0;
assign v$A_7526_out0 = v$A19_1368_out0;
assign v$A_7527_out0 = v$A22_4595_out0;
assign v$A_7529_out0 = v$A10_1708_out0;
assign v$A_7530_out0 = v$A20_4608_out0;
assign v$A_7531_out0 = v$A2_18873_out0;
assign v$A_7532_out0 = v$A11_10391_out0;
assign v$A_7533_out0 = v$A5_6906_out0;
assign v$A_7534_out0 = v$A16_14196_out0;
assign v$END_12506_out0 = v$_2613_out1;
assign v$END_12724_out0 = v$_2810_out1;
assign v$G1_12950_out0 = v$A_7439_out0 && v$B_2944_out0;
assign v$G1_12951_out0 = v$A_7440_out0 && v$B_2945_out0;
assign v$G1_12952_out0 = v$A_7441_out0 && v$B_2946_out0;
assign v$G1_12953_out0 = v$A_7442_out0 && v$B_2947_out0;
assign v$G1_12954_out0 = v$A_7443_out0 && v$B_2948_out0;
assign v$G1_12958_out0 = v$A_7447_out0 && v$B_2952_out0;
assign v$G1_12962_out0 = v$A_7451_out0 && v$B_2956_out0;
assign v$G1_12967_out0 = v$A_7456_out0 && v$B_2961_out0;
assign v$G1_13022_out0 = v$A_7511_out0 && v$B_3016_out0;
assign v$G1_13023_out0 = v$A_7512_out0 && v$B_3017_out0;
assign v$G1_13024_out0 = v$A_7513_out0 && v$B_3018_out0;
assign v$G1_13025_out0 = v$A_7514_out0 && v$B_3019_out0;
assign v$G1_13026_out0 = v$A_7515_out0 && v$B_3020_out0;
assign v$G1_13030_out0 = v$A_7519_out0 && v$B_3024_out0;
assign v$G1_13034_out0 = v$A_7523_out0 && v$B_3028_out0;
assign v$G1_13039_out0 = v$A_7528_out0 && v$B_3033_out0;
assign v$END_18877_out0 = v$A1A_12226_out1;
assign v$END_18880_out0 = v$A1A_12229_out1;
assign v$MUX2_2688_out0 = v$EN_1493_out0 ? v$MUX1_2543_out0 : v$IN_5233_out0;
assign v$MUX2_2690_out0 = v$EN_1495_out0 ? v$MUX1_2548_out0 : v$IN_5235_out0;
assign v$MUX2_2698_out0 = v$EN_1503_out0 ? v$MUX1_2574_out0 : v$IN_5243_out0;
assign v$MUX2_2700_out0 = v$EN_1505_out0 ? v$MUX1_2579_out0 : v$IN_5245_out0;
assign v$G2_5531_out0 = ((v$A_7444_out0 && !v$B_2949_out0) || (!v$A_7444_out0) && v$B_2949_out0);
assign v$G2_5532_out0 = ((v$A_7445_out0 && !v$B_2950_out0) || (!v$A_7445_out0) && v$B_2950_out0);
assign v$G2_5533_out0 = ((v$A_7446_out0 && !v$B_2951_out0) || (!v$A_7446_out0) && v$B_2951_out0);
assign v$G2_5535_out0 = ((v$A_7448_out0 && !v$B_2953_out0) || (!v$A_7448_out0) && v$B_2953_out0);
assign v$G2_5536_out0 = ((v$A_7449_out0 && !v$B_2954_out0) || (!v$A_7449_out0) && v$B_2954_out0);
assign v$G2_5537_out0 = ((v$A_7450_out0 && !v$B_2955_out0) || (!v$A_7450_out0) && v$B_2955_out0);
assign v$G2_5539_out0 = ((v$A_7452_out0 && !v$B_2957_out0) || (!v$A_7452_out0) && v$B_2957_out0);
assign v$G2_5540_out0 = ((v$A_7453_out0 && !v$B_2958_out0) || (!v$A_7453_out0) && v$B_2958_out0);
assign v$G2_5541_out0 = ((v$A_7454_out0 && !v$B_2959_out0) || (!v$A_7454_out0) && v$B_2959_out0);
assign v$G2_5542_out0 = ((v$A_7455_out0 && !v$B_2960_out0) || (!v$A_7455_out0) && v$B_2960_out0);
assign v$G2_5544_out0 = ((v$A_7457_out0 && !v$B_2962_out0) || (!v$A_7457_out0) && v$B_2962_out0);
assign v$G2_5545_out0 = ((v$A_7458_out0 && !v$B_2963_out0) || (!v$A_7458_out0) && v$B_2963_out0);
assign v$G2_5546_out0 = ((v$A_7459_out0 && !v$B_2964_out0) || (!v$A_7459_out0) && v$B_2964_out0);
assign v$G2_5547_out0 = ((v$A_7460_out0 && !v$B_2965_out0) || (!v$A_7460_out0) && v$B_2965_out0);
assign v$G2_5548_out0 = ((v$A_7461_out0 && !v$B_2966_out0) || (!v$A_7461_out0) && v$B_2966_out0);
assign v$G2_5549_out0 = ((v$A_7462_out0 && !v$B_2967_out0) || (!v$A_7462_out0) && v$B_2967_out0);
assign v$G2_5603_out0 = ((v$A_7516_out0 && !v$B_3021_out0) || (!v$A_7516_out0) && v$B_3021_out0);
assign v$G2_5604_out0 = ((v$A_7517_out0 && !v$B_3022_out0) || (!v$A_7517_out0) && v$B_3022_out0);
assign v$G2_5605_out0 = ((v$A_7518_out0 && !v$B_3023_out0) || (!v$A_7518_out0) && v$B_3023_out0);
assign v$G2_5607_out0 = ((v$A_7520_out0 && !v$B_3025_out0) || (!v$A_7520_out0) && v$B_3025_out0);
assign v$G2_5608_out0 = ((v$A_7521_out0 && !v$B_3026_out0) || (!v$A_7521_out0) && v$B_3026_out0);
assign v$G2_5609_out0 = ((v$A_7522_out0 && !v$B_3027_out0) || (!v$A_7522_out0) && v$B_3027_out0);
assign v$G2_5611_out0 = ((v$A_7524_out0 && !v$B_3029_out0) || (!v$A_7524_out0) && v$B_3029_out0);
assign v$G2_5612_out0 = ((v$A_7525_out0 && !v$B_3030_out0) || (!v$A_7525_out0) && v$B_3030_out0);
assign v$G2_5613_out0 = ((v$A_7526_out0 && !v$B_3031_out0) || (!v$A_7526_out0) && v$B_3031_out0);
assign v$G2_5614_out0 = ((v$A_7527_out0 && !v$B_3032_out0) || (!v$A_7527_out0) && v$B_3032_out0);
assign v$G2_5616_out0 = ((v$A_7529_out0 && !v$B_3034_out0) || (!v$A_7529_out0) && v$B_3034_out0);
assign v$G2_5617_out0 = ((v$A_7530_out0 && !v$B_3035_out0) || (!v$A_7530_out0) && v$B_3035_out0);
assign v$G2_5618_out0 = ((v$A_7531_out0 && !v$B_3036_out0) || (!v$A_7531_out0) && v$B_3036_out0);
assign v$G2_5619_out0 = ((v$A_7532_out0 && !v$B_3037_out0) || (!v$A_7532_out0) && v$B_3037_out0);
assign v$G2_5620_out0 = ((v$A_7533_out0 && !v$B_3038_out0) || (!v$A_7533_out0) && v$B_3038_out0);
assign v$G2_5621_out0 = ((v$A_7534_out0 && !v$B_3039_out0) || (!v$A_7534_out0) && v$B_3039_out0);
assign v$G_10530_out0 = v$G1_12950_out0;
assign v$G_10531_out0 = v$G1_12951_out0;
assign v$G_10532_out0 = v$G1_12952_out0;
assign v$G_10533_out0 = v$G1_12953_out0;
assign v$G_10534_out0 = v$G1_12954_out0;
assign v$G_10538_out0 = v$G1_12958_out0;
assign v$G_10542_out0 = v$G1_12962_out0;
assign v$G_10547_out0 = v$G1_12967_out0;
assign v$G_10602_out0 = v$G1_13022_out0;
assign v$G_10603_out0 = v$G1_13023_out0;
assign v$G_10604_out0 = v$G1_13024_out0;
assign v$G_10605_out0 = v$G1_13025_out0;
assign v$G_10606_out0 = v$G1_13026_out0;
assign v$G_10610_out0 = v$G1_13030_out0;
assign v$G_10614_out0 = v$G1_13034_out0;
assign v$G_10619_out0 = v$G1_13039_out0;
assign v$G1_12955_out0 = v$A_7444_out0 && v$B_2949_out0;
assign v$G1_12956_out0 = v$A_7445_out0 && v$B_2950_out0;
assign v$G1_12957_out0 = v$A_7446_out0 && v$B_2951_out0;
assign v$G1_12959_out0 = v$A_7448_out0 && v$B_2953_out0;
assign v$G1_12960_out0 = v$A_7449_out0 && v$B_2954_out0;
assign v$G1_12961_out0 = v$A_7450_out0 && v$B_2955_out0;
assign v$G1_12963_out0 = v$A_7452_out0 && v$B_2957_out0;
assign v$G1_12964_out0 = v$A_7453_out0 && v$B_2958_out0;
assign v$G1_12965_out0 = v$A_7454_out0 && v$B_2959_out0;
assign v$G1_12966_out0 = v$A_7455_out0 && v$B_2960_out0;
assign v$G1_12968_out0 = v$A_7457_out0 && v$B_2962_out0;
assign v$G1_12969_out0 = v$A_7458_out0 && v$B_2963_out0;
assign v$G1_12970_out0 = v$A_7459_out0 && v$B_2964_out0;
assign v$G1_12971_out0 = v$A_7460_out0 && v$B_2965_out0;
assign v$G1_12972_out0 = v$A_7461_out0 && v$B_2966_out0;
assign v$G1_12973_out0 = v$A_7462_out0 && v$B_2967_out0;
assign v$G1_13027_out0 = v$A_7516_out0 && v$B_3021_out0;
assign v$G1_13028_out0 = v$A_7517_out0 && v$B_3022_out0;
assign v$G1_13029_out0 = v$A_7518_out0 && v$B_3023_out0;
assign v$G1_13031_out0 = v$A_7520_out0 && v$B_3025_out0;
assign v$G1_13032_out0 = v$A_7521_out0 && v$B_3026_out0;
assign v$G1_13033_out0 = v$A_7522_out0 && v$B_3027_out0;
assign v$G1_13035_out0 = v$A_7524_out0 && v$B_3029_out0;
assign v$G1_13036_out0 = v$A_7525_out0 && v$B_3030_out0;
assign v$G1_13037_out0 = v$A_7526_out0 && v$B_3031_out0;
assign v$G1_13038_out0 = v$A_7527_out0 && v$B_3032_out0;
assign v$G1_13040_out0 = v$A_7529_out0 && v$B_3034_out0;
assign v$G1_13041_out0 = v$A_7530_out0 && v$B_3035_out0;
assign v$G1_13042_out0 = v$A_7531_out0 && v$B_3036_out0;
assign v$G1_13043_out0 = v$A_7532_out0 && v$B_3037_out0;
assign v$G1_13044_out0 = v$A_7533_out0 && v$B_3038_out0;
assign v$G1_13045_out0 = v$A_7534_out0 && v$B_3039_out0;
assign v$P_14501_out0 = v$G2_5526_out0;
assign v$P_14502_out0 = v$G2_5527_out0;
assign v$P_14503_out0 = v$G2_5528_out0;
assign v$P_14504_out0 = v$G2_5529_out0;
assign v$P_14505_out0 = v$G2_5530_out0;
assign v$P_14509_out0 = v$G2_5534_out0;
assign v$P_14513_out0 = v$G2_5538_out0;
assign v$P_14518_out0 = v$G2_5543_out0;
assign v$P_14573_out0 = v$G2_5598_out0;
assign v$P_14574_out0 = v$G2_5599_out0;
assign v$P_14575_out0 = v$G2_5600_out0;
assign v$P_14576_out0 = v$G2_5601_out0;
assign v$P_14577_out0 = v$G2_5602_out0;
assign v$P_14581_out0 = v$G2_5606_out0;
assign v$P_14585_out0 = v$G2_5610_out0;
assign v$P_14590_out0 = v$G2_5615_out0;
assign v$P12_245_out0 = v$P_14509_out0;
assign v$P12_248_out0 = v$P_14581_out0;
assign v$P21_4983_out0 = v$P_14503_out0;
assign v$P21_4986_out0 = v$P_14575_out0;
assign v$P0_5025_out0 = v$P_14513_out0;
assign v$P0_5028_out0 = v$P_14585_out0;
assign v$P15_7185_out0 = v$P_14505_out0;
assign v$P15_7188_out0 = v$P_14577_out0;
assign v$G12_7329_out0 = v$G_10538_out0;
assign v$G12_7332_out0 = v$G_10610_out0;
assign v$P6_8420_out0 = v$P_14501_out0;
assign v$P6_8423_out0 = v$P_14573_out0;
assign v$G9_9257_out0 = v$G_10533_out0;
assign v$G9_9260_out0 = v$G_10605_out0;
assign v$G_10535_out0 = v$G1_12955_out0;
assign v$G_10536_out0 = v$G1_12956_out0;
assign v$G_10537_out0 = v$G1_12957_out0;
assign v$G_10539_out0 = v$G1_12959_out0;
assign v$G_10540_out0 = v$G1_12960_out0;
assign v$G_10541_out0 = v$G1_12961_out0;
assign v$G_10543_out0 = v$G1_12963_out0;
assign v$G_10544_out0 = v$G1_12964_out0;
assign v$G_10545_out0 = v$G1_12965_out0;
assign v$G_10546_out0 = v$G1_12966_out0;
assign v$G_10548_out0 = v$G1_12968_out0;
assign v$G_10549_out0 = v$G1_12969_out0;
assign v$G_10550_out0 = v$G1_12970_out0;
assign v$G_10551_out0 = v$G1_12971_out0;
assign v$G_10552_out0 = v$G1_12972_out0;
assign v$G_10553_out0 = v$G1_12973_out0;
assign v$G_10607_out0 = v$G1_13027_out0;
assign v$G_10608_out0 = v$G1_13028_out0;
assign v$G_10609_out0 = v$G1_13029_out0;
assign v$G_10611_out0 = v$G1_13031_out0;
assign v$G_10612_out0 = v$G1_13032_out0;
assign v$G_10613_out0 = v$G1_13033_out0;
assign v$G_10615_out0 = v$G1_13035_out0;
assign v$G_10616_out0 = v$G1_13036_out0;
assign v$G_10617_out0 = v$G1_13037_out0;
assign v$G_10618_out0 = v$G1_13038_out0;
assign v$G_10620_out0 = v$G1_13040_out0;
assign v$G_10621_out0 = v$G1_13041_out0;
assign v$G_10622_out0 = v$G1_13042_out0;
assign v$G_10623_out0 = v$G1_13043_out0;
assign v$G_10624_out0 = v$G1_13044_out0;
assign v$G_10625_out0 = v$G1_13045_out0;
assign v$G15_11543_out0 = v$G_10534_out0;
assign v$G15_11546_out0 = v$G_10606_out0;
assign v$G3_11604_out0 = v$G_10531_out0;
assign v$G3_11607_out0 = v$G_10603_out0;
assign v$P18_12292_out0 = v$P_14518_out0;
assign v$P18_12295_out0 = v$P_14590_out0;
assign v$G18_13510_out0 = v$G_10547_out0;
assign v$G18_13513_out0 = v$G_10619_out0;
assign v$P_14506_out0 = v$G2_5531_out0;
assign v$P_14507_out0 = v$G2_5532_out0;
assign v$P_14508_out0 = v$G2_5533_out0;
assign v$P_14510_out0 = v$G2_5535_out0;
assign v$P_14511_out0 = v$G2_5536_out0;
assign v$P_14512_out0 = v$G2_5537_out0;
assign v$P_14514_out0 = v$G2_5539_out0;
assign v$P_14515_out0 = v$G2_5540_out0;
assign v$P_14516_out0 = v$G2_5541_out0;
assign v$P_14517_out0 = v$G2_5542_out0;
assign v$P_14519_out0 = v$G2_5544_out0;
assign v$P_14520_out0 = v$G2_5545_out0;
assign v$P_14521_out0 = v$G2_5546_out0;
assign v$P_14522_out0 = v$G2_5547_out0;
assign v$P_14523_out0 = v$G2_5548_out0;
assign v$P_14524_out0 = v$G2_5549_out0;
assign v$P_14578_out0 = v$G2_5603_out0;
assign v$P_14579_out0 = v$G2_5604_out0;
assign v$P_14580_out0 = v$G2_5605_out0;
assign v$P_14582_out0 = v$G2_5607_out0;
assign v$P_14583_out0 = v$G2_5608_out0;
assign v$P_14584_out0 = v$G2_5609_out0;
assign v$P_14586_out0 = v$G2_5611_out0;
assign v$P_14587_out0 = v$G2_5612_out0;
assign v$P_14588_out0 = v$G2_5613_out0;
assign v$P_14589_out0 = v$G2_5614_out0;
assign v$P_14591_out0 = v$G2_5616_out0;
assign v$P_14592_out0 = v$G2_5617_out0;
assign v$P_14593_out0 = v$G2_5618_out0;
assign v$P_14594_out0 = v$G2_5619_out0;
assign v$P_14595_out0 = v$G2_5620_out0;
assign v$P_14596_out0 = v$G2_5621_out0;
assign v$G21_14628_out0 = v$G_10532_out0;
assign v$G21_14631_out0 = v$G_10604_out0;
assign v$OUT_15515_out0 = v$MUX2_2688_out0;
assign v$OUT_15520_out0 = v$MUX2_2690_out0;
assign v$OUT_15546_out0 = v$MUX2_2698_out0;
assign v$OUT_15551_out0 = v$MUX2_2700_out0;
assign v$P3_15923_out0 = v$P_14502_out0;
assign v$P3_15926_out0 = v$P_14574_out0;
assign v$G0_16550_out0 = v$G_10542_out0;
assign v$G0_16553_out0 = v$G_10614_out0;
assign v$G6_16972_out0 = v$G_10530_out0;
assign v$G6_16975_out0 = v$G_10602_out0;
assign v$P9_19055_out0 = v$P_14504_out0;
assign v$P9_19058_out0 = v$P_14576_out0;
assign v$P5_230_out0 = v$P_14523_out0;
assign v$P5_233_out0 = v$P_14595_out0;
assign v$P10_362_out0 = v$P_14519_out0;
assign v$P10_365_out0 = v$P_14591_out0;
assign v$G$CD_1109_out0 = v$G6_16972_out0;
assign v$G$CD_1110_out0 = v$G3_11604_out0;
assign v$G$CD_1111_out0 = v$G12_7329_out0;
assign v$G$CD_1112_out0 = v$G9_9257_out0;
assign v$G$CD_1115_out0 = v$G18_13510_out0;
assign v$G$CD_1126_out0 = v$G15_11543_out0;
assign v$G$CD_1127_out0 = v$G21_14628_out0;
assign v$G$CD_1232_out0 = v$G6_16975_out0;
assign v$G$CD_1233_out0 = v$G3_11607_out0;
assign v$G$CD_1234_out0 = v$G12_7332_out0;
assign v$G$CD_1235_out0 = v$G9_9260_out0;
assign v$G$CD_1238_out0 = v$G18_13513_out0;
assign v$G$CD_1249_out0 = v$G15_11546_out0;
assign v$G$CD_1250_out0 = v$G21_14631_out0;
assign v$G7_1851_out0 = v$G_10535_out0;
assign v$G7_1854_out0 = v$G_10607_out0;
assign v$P8_1863_out0 = v$P_14510_out0;
assign v$P8_1866_out0 = v$P_14582_out0;
assign v$G10_1995_out0 = v$G_10548_out0;
assign v$G10_1998_out0 = v$G_10620_out0;
assign v$G19_2046_out0 = v$G_10545_out0;
assign v$G19_2049_out0 = v$G_10617_out0;
assign v$P$AB_2250_out0 = v$P0_5025_out0;
assign v$P$AB_2253_out0 = v$P18_12292_out0;
assign v$P$AB_2254_out0 = v$P21_4983_out0;
assign v$P$AB_2266_out0 = v$P12_245_out0;
assign v$P$AB_2268_out0 = v$P15_7185_out0;
assign v$P$AB_2271_out0 = v$P6_8420_out0;
assign v$P$AB_2277_out0 = v$P3_15923_out0;
assign v$P$AB_2282_out0 = v$P9_19055_out0;
assign v$P$AB_2373_out0 = v$P0_5028_out0;
assign v$P$AB_2376_out0 = v$P18_12295_out0;
assign v$P$AB_2377_out0 = v$P21_4986_out0;
assign v$P$AB_2389_out0 = v$P12_248_out0;
assign v$P$AB_2391_out0 = v$P15_7188_out0;
assign v$P$AB_2394_out0 = v$P6_8423_out0;
assign v$P$AB_2400_out0 = v$P3_15926_out0;
assign v$P$AB_2405_out0 = v$P9_19058_out0;
assign v$P2_2426_out0 = v$P_14521_out0;
assign v$P2_2429_out0 = v$P_14593_out0;
assign v$G8_2772_out0 = v$G_10539_out0;
assign v$G8_2775_out0 = v$G_10611_out0;
assign v$G13_3054_out0 = v$G_10543_out0;
assign v$G13_3057_out0 = v$G_10615_out0;
assign v$P1_3170_out0 = v$P_14507_out0;
assign v$P1_3173_out0 = v$P_14579_out0;
assign v$P13_3247_out0 = v$P_14514_out0;
assign v$P13_3250_out0 = v$P_14586_out0;
assign v$P14_3371_out0 = v$P_14508_out0;
assign v$P14_3374_out0 = v$P_14580_out0;
assign v$P22_4947_out0 = v$P_14517_out0;
assign v$P22_4950_out0 = v$P_14589_out0;
assign v$G1_5271_out0 = v$G_10536_out0;
assign v$G1_5274_out0 = v$G_10608_out0;
assign v$G4_6021_out0 = v$G_10544_out0;
assign v$G4_6024_out0 = v$G_10616_out0;
assign v$P23_6628_out0 = v$P_14512_out0;
assign v$P23_6631_out0 = v$P_14584_out0;
assign v$P16_7245_out0 = v$P_14524_out0;
assign v$P16_7248_out0 = v$P_14596_out0;
assign v$G20_8535_out0 = v$G_10549_out0;
assign v$G20_8538_out0 = v$G_10621_out0;
assign v$G$AB_9550_out0 = v$G0_16550_out0;
assign v$G$AB_9553_out0 = v$G18_13510_out0;
assign v$G$AB_9554_out0 = v$G21_14628_out0;
assign v$G$AB_9566_out0 = v$G12_7329_out0;
assign v$G$AB_9568_out0 = v$G15_11543_out0;
assign v$G$AB_9571_out0 = v$G6_16972_out0;
assign v$G$AB_9577_out0 = v$G3_11604_out0;
assign v$G$AB_9582_out0 = v$G9_9257_out0;
assign v$G$AB_9673_out0 = v$G0_16553_out0;
assign v$G$AB_9676_out0 = v$G18_13513_out0;
assign v$G$AB_9677_out0 = v$G21_14631_out0;
assign v$G$AB_9689_out0 = v$G12_7332_out0;
assign v$G$AB_9691_out0 = v$G15_11546_out0;
assign v$G$AB_9694_out0 = v$G6_16975_out0;
assign v$G$AB_9700_out0 = v$G3_11607_out0;
assign v$G$AB_9705_out0 = v$G9_9260_out0;
assign v$G17_9716_out0 = v$G_10540_out0;
assign v$G17_9719_out0 = v$G_10612_out0;
assign v$P11_9994_out0 = v$P_14522_out0;
assign v$P11_9997_out0 = v$P_14594_out0;
assign v$P$CD_10998_out0 = v$P6_8420_out0;
assign v$P$CD_10999_out0 = v$P3_15923_out0;
assign v$P$CD_11000_out0 = v$P12_245_out0;
assign v$P$CD_11001_out0 = v$P9_19055_out0;
assign v$P$CD_11004_out0 = v$P18_12292_out0;
assign v$P$CD_11015_out0 = v$P15_7185_out0;
assign v$P$CD_11016_out0 = v$P21_4983_out0;
assign v$P$CD_11121_out0 = v$P6_8423_out0;
assign v$P$CD_11122_out0 = v$P3_15926_out0;
assign v$P$CD_11123_out0 = v$P12_248_out0;
assign v$P$CD_11124_out0 = v$P9_19058_out0;
assign v$P$CD_11127_out0 = v$P18_12295_out0;
assign v$P$CD_11138_out0 = v$P15_7188_out0;
assign v$P$CD_11139_out0 = v$P21_4986_out0;
assign v$P20_11154_out0 = v$P_14520_out0;
assign v$P20_11157_out0 = v$P_14592_out0;
assign v$G5_11172_out0 = v$G_10552_out0;
assign v$G5_11175_out0 = v$G_10624_out0;
assign v$G11_11577_out0 = v$G_10551_out0;
assign v$G11_11580_out0 = v$G_10623_out0;
assign v$MUX1_12191_out0 = v$G2_18054_out0 ? v$C1_4623_out0 : v$OUT_15515_out0;
assign v$MUX1_12192_out0 = v$G2_18055_out0 ? v$C1_4624_out0 : v$OUT_15520_out0;
assign v$MUX1_12195_out0 = v$G2_18058_out0 ? v$C1_4627_out0 : v$OUT_15546_out0;
assign v$MUX1_12196_out0 = v$G2_18059_out0 ? v$C1_4628_out0 : v$OUT_15551_out0;
assign v$P17_12330_out0 = v$P_14511_out0;
assign v$P17_12333_out0 = v$P_14583_out0;
assign v$P7_12340_out0 = v$P_14506_out0;
assign v$P7_12343_out0 = v$P_14578_out0;
assign v$G22_13106_out0 = v$G_10546_out0;
assign v$G22_13109_out0 = v$G_10618_out0;
assign v$P4_14216_out0 = v$P_14515_out0;
assign v$P4_14219_out0 = v$P_14587_out0;
assign v$G23_14922_out0 = v$G_10541_out0;
assign v$G23_14925_out0 = v$G_10613_out0;
assign v$GATE2_16357_out0 = v$CIN_16719_out0 && v$P0_5025_out0;
assign v$GATE2_16360_out0 = v$CIN_16722_out0 && v$P0_5028_out0;
assign v$G2_16570_out0 = v$G_10550_out0;
assign v$G2_16573_out0 = v$G_10622_out0;
assign v$P19_16934_out0 = v$P_14516_out0;
assign v$P19_16937_out0 = v$P_14588_out0;
assign v$G16_17073_out0 = v$G_10553_out0;
assign v$G16_17076_out0 = v$G_10625_out0;
assign v$G14_18595_out0 = v$G_10537_out0;
assign v$G14_18598_out0 = v$G_10609_out0;
assign v$GATE1_722_out0 = v$GATE2_16357_out0 || v$G0_16550_out0;
assign v$GATE1_725_out0 = v$GATE2_16360_out0 || v$G0_16553_out0;
assign v$G$CD_1100_out0 = v$G14_18595_out0;
assign v$G$CD_1101_out0 = v$G8_2772_out0;
assign v$G$CD_1103_out0 = v$G1_5271_out0;
assign v$G$CD_1106_out0 = v$G19_2046_out0;
assign v$G$CD_1107_out0 = v$G22_13106_out0;
assign v$G$CD_1114_out0 = v$G23_14922_out0;
assign v$G$CD_1116_out0 = v$G2_16570_out0;
assign v$G$CD_1117_out0 = v$G5_11172_out0;
assign v$G$CD_1119_out0 = v$G13_3054_out0;
assign v$G$CD_1120_out0 = v$G17_9716_out0;
assign v$G$CD_1121_out0 = v$G16_17073_out0;
assign v$G$CD_1124_out0 = v$G7_1851_out0;
assign v$G$CD_1130_out0 = v$G4_6021_out0;
assign v$G$CD_1134_out0 = v$G20_8535_out0;
assign v$G$CD_1135_out0 = v$G10_1995_out0;
assign v$G$CD_1139_out0 = v$G11_11577_out0;
assign v$G$CD_1223_out0 = v$G14_18598_out0;
assign v$G$CD_1224_out0 = v$G8_2775_out0;
assign v$G$CD_1226_out0 = v$G1_5274_out0;
assign v$G$CD_1229_out0 = v$G19_2049_out0;
assign v$G$CD_1230_out0 = v$G22_13109_out0;
assign v$G$CD_1237_out0 = v$G23_14925_out0;
assign v$G$CD_1239_out0 = v$G2_16573_out0;
assign v$G$CD_1240_out0 = v$G5_11175_out0;
assign v$G$CD_1242_out0 = v$G13_3057_out0;
assign v$G$CD_1243_out0 = v$G17_9719_out0;
assign v$G$CD_1244_out0 = v$G16_17076_out0;
assign v$G$CD_1247_out0 = v$G7_1854_out0;
assign v$G$CD_1253_out0 = v$G4_6024_out0;
assign v$G$CD_1257_out0 = v$G20_8538_out0;
assign v$G$CD_1258_out0 = v$G10_1998_out0;
assign v$G$CD_1262_out0 = v$G11_11580_out0;
assign v$OUT_10436_out0 = v$MUX1_12191_out0;
assign v$OUT_10437_out0 = v$MUX1_12192_out0;
assign v$OUT_10440_out0 = v$MUX1_12195_out0;
assign v$OUT_10441_out0 = v$MUX1_12196_out0;
assign v$P$CD_10989_out0 = v$P14_3371_out0;
assign v$P$CD_10990_out0 = v$P8_1863_out0;
assign v$P$CD_10992_out0 = v$P1_3170_out0;
assign v$P$CD_10995_out0 = v$P19_16934_out0;
assign v$P$CD_10996_out0 = v$P22_4947_out0;
assign v$P$CD_11003_out0 = v$P23_6628_out0;
assign v$P$CD_11005_out0 = v$P2_2426_out0;
assign v$P$CD_11006_out0 = v$P5_230_out0;
assign v$P$CD_11008_out0 = v$P13_3247_out0;
assign v$P$CD_11009_out0 = v$P17_12330_out0;
assign v$P$CD_11010_out0 = v$P16_7245_out0;
assign v$P$CD_11013_out0 = v$P7_12340_out0;
assign v$P$CD_11019_out0 = v$P4_14216_out0;
assign v$P$CD_11023_out0 = v$P20_11154_out0;
assign v$P$CD_11024_out0 = v$P10_362_out0;
assign v$P$CD_11028_out0 = v$P11_9994_out0;
assign v$P$CD_11112_out0 = v$P14_3374_out0;
assign v$P$CD_11113_out0 = v$P8_1866_out0;
assign v$P$CD_11115_out0 = v$P1_3173_out0;
assign v$P$CD_11118_out0 = v$P19_16937_out0;
assign v$P$CD_11119_out0 = v$P22_4950_out0;
assign v$P$CD_11126_out0 = v$P23_6631_out0;
assign v$P$CD_11128_out0 = v$P2_2429_out0;
assign v$P$CD_11129_out0 = v$P5_233_out0;
assign v$P$CD_11131_out0 = v$P13_3250_out0;
assign v$P$CD_11132_out0 = v$P17_12333_out0;
assign v$P$CD_11133_out0 = v$P16_7248_out0;
assign v$P$CD_11136_out0 = v$P7_12343_out0;
assign v$P$CD_11142_out0 = v$P4_14219_out0;
assign v$P$CD_11146_out0 = v$P20_11157_out0;
assign v$P$CD_11147_out0 = v$P10_365_out0;
assign v$P$CD_11151_out0 = v$P11_9997_out0;
assign v$G8_12011_out0 = v$CINA_8856_out0 && v$P$AB_2250_out0;
assign v$G8_12014_out0 = v$CINA_8859_out0 && v$P$AB_2253_out0;
assign v$G8_12015_out0 = v$CINA_8860_out0 && v$P$AB_2254_out0;
assign v$G8_12027_out0 = v$CINA_8872_out0 && v$P$AB_2266_out0;
assign v$G8_12029_out0 = v$CINA_8874_out0 && v$P$AB_2268_out0;
assign v$G8_12032_out0 = v$CINA_8877_out0 && v$P$AB_2271_out0;
assign v$G8_12038_out0 = v$CINA_8883_out0 && v$P$AB_2277_out0;
assign v$G8_12043_out0 = v$CINA_8888_out0 && v$P$AB_2282_out0;
assign v$G8_12134_out0 = v$CINA_8979_out0 && v$P$AB_2373_out0;
assign v$G8_12137_out0 = v$CINA_8982_out0 && v$P$AB_2376_out0;
assign v$G8_12138_out0 = v$CINA_8983_out0 && v$P$AB_2377_out0;
assign v$G8_12150_out0 = v$CINA_8995_out0 && v$P$AB_2389_out0;
assign v$G8_12152_out0 = v$CINA_8997_out0 && v$P$AB_2391_out0;
assign v$G8_12155_out0 = v$CINA_9000_out0 && v$P$AB_2394_out0;
assign v$G8_12161_out0 = v$CINA_9006_out0 && v$P$AB_2400_out0;
assign v$G8_12166_out0 = v$CINA_9011_out0 && v$P$AB_2405_out0;
assign v$G5_4775_out0 = v$G$AB_9550_out0 && v$P$CD_10992_out0;
assign v$G5_4778_out0 = v$G$AB_9553_out0 && v$P$CD_10995_out0;
assign v$G5_4779_out0 = v$G$AB_9554_out0 && v$P$CD_10996_out0;
assign v$G5_4791_out0 = v$G$AB_9566_out0 && v$P$CD_11008_out0;
assign v$G5_4793_out0 = v$G$AB_9568_out0 && v$P$CD_11010_out0;
assign v$G5_4796_out0 = v$G$AB_9571_out0 && v$P$CD_11013_out0;
assign v$G5_4802_out0 = v$G$AB_9577_out0 && v$P$CD_11019_out0;
assign v$G5_4807_out0 = v$G$AB_9582_out0 && v$P$CD_11024_out0;
assign v$G5_4898_out0 = v$G$AB_9673_out0 && v$P$CD_11115_out0;
assign v$G5_4901_out0 = v$G$AB_9676_out0 && v$P$CD_11118_out0;
assign v$G5_4902_out0 = v$G$AB_9677_out0 && v$P$CD_11119_out0;
assign v$G5_4914_out0 = v$G$AB_9689_out0 && v$P$CD_11131_out0;
assign v$G5_4916_out0 = v$G$AB_9691_out0 && v$P$CD_11133_out0;
assign v$G5_4919_out0 = v$G$AB_9694_out0 && v$P$CD_11136_out0;
assign v$G5_4925_out0 = v$G$AB_9700_out0 && v$P$CD_11142_out0;
assign v$G5_4930_out0 = v$G$AB_9705_out0 && v$P$CD_11147_out0;
assign v$G1_5849_out0 = v$P$AB_2250_out0 && v$P$CD_10992_out0;
assign v$G1_5852_out0 = v$P$AB_2253_out0 && v$P$CD_10995_out0;
assign v$G1_5853_out0 = v$P$AB_2254_out0 && v$P$CD_10996_out0;
assign v$G1_5865_out0 = v$P$AB_2266_out0 && v$P$CD_11008_out0;
assign v$G1_5867_out0 = v$P$AB_2268_out0 && v$P$CD_11010_out0;
assign v$G1_5870_out0 = v$P$AB_2271_out0 && v$P$CD_11013_out0;
assign v$G1_5876_out0 = v$P$AB_2277_out0 && v$P$CD_11019_out0;
assign v$G1_5881_out0 = v$P$AB_2282_out0 && v$P$CD_11024_out0;
assign v$G1_5972_out0 = v$P$AB_2373_out0 && v$P$CD_11115_out0;
assign v$G1_5975_out0 = v$P$AB_2376_out0 && v$P$CD_11118_out0;
assign v$G1_5976_out0 = v$P$AB_2377_out0 && v$P$CD_11119_out0;
assign v$G1_5988_out0 = v$P$AB_2389_out0 && v$P$CD_11131_out0;
assign v$G1_5990_out0 = v$P$AB_2391_out0 && v$P$CD_11133_out0;
assign v$G1_5993_out0 = v$P$AB_2394_out0 && v$P$CD_11136_out0;
assign v$G1_5999_out0 = v$P$AB_2400_out0 && v$P$CD_11142_out0;
assign v$G1_6004_out0 = v$P$AB_2405_out0 && v$P$CD_11147_out0;
assign v$MUX4_6167_out0 = v$NEED$SHIFT$OP1_5034_out0 ? v$OUT_10437_out0 : v$OP1$MANTISA_12378_out0;
assign v$MUX4_6168_out0 = v$NEED$SHIFT$OP1_5035_out0 ? v$OUT_10441_out0 : v$OP1$MANTISA_12379_out0;
assign v$G7_10103_out0 = v$G8_12011_out0 && v$P$CD_10992_out0;
assign v$G7_10106_out0 = v$G8_12014_out0 && v$P$CD_10995_out0;
assign v$G7_10107_out0 = v$G8_12015_out0 && v$P$CD_10996_out0;
assign v$G7_10119_out0 = v$G8_12027_out0 && v$P$CD_11008_out0;
assign v$G7_10121_out0 = v$G8_12029_out0 && v$P$CD_11010_out0;
assign v$G7_10124_out0 = v$G8_12032_out0 && v$P$CD_11013_out0;
assign v$G7_10130_out0 = v$G8_12038_out0 && v$P$CD_11019_out0;
assign v$G7_10135_out0 = v$G8_12043_out0 && v$P$CD_11024_out0;
assign v$G7_10226_out0 = v$G8_12134_out0 && v$P$CD_11115_out0;
assign v$G7_10229_out0 = v$G8_12137_out0 && v$P$CD_11118_out0;
assign v$G7_10230_out0 = v$G8_12138_out0 && v$P$CD_11119_out0;
assign v$G7_10242_out0 = v$G8_12150_out0 && v$P$CD_11131_out0;
assign v$G7_10244_out0 = v$G8_12152_out0 && v$P$CD_11133_out0;
assign v$G7_10247_out0 = v$G8_12155_out0 && v$P$CD_11136_out0;
assign v$G7_10253_out0 = v$G8_12161_out0 && v$P$CD_11142_out0;
assign v$G7_10258_out0 = v$G8_12166_out0 && v$P$CD_11147_out0;
assign v$C0_11190_out0 = v$GATE1_722_out0;
assign v$C0_11193_out0 = v$GATE1_725_out0;
assign v$MUX1_14796_out0 = v$NEED$SHIFT$OP1_5034_out0 ? v$OP2$MANTISA_3710_out0 : v$OUT_10436_out0;
assign v$MUX1_14797_out0 = v$NEED$SHIFT$OP1_5035_out0 ? v$OP2$MANTISA_3711_out0 : v$OUT_10440_out0;
assign v$P$AD_836_out0 = v$G1_5849_out0;
assign v$P$AD_839_out0 = v$G1_5852_out0;
assign v$P$AD_840_out0 = v$G1_5853_out0;
assign v$P$AD_852_out0 = v$G1_5865_out0;
assign v$P$AD_854_out0 = v$G1_5867_out0;
assign v$P$AD_857_out0 = v$G1_5870_out0;
assign v$P$AD_863_out0 = v$G1_5876_out0;
assign v$P$AD_868_out0 = v$G1_5881_out0;
assign v$P$AD_959_out0 = v$G1_5972_out0;
assign v$P$AD_962_out0 = v$G1_5975_out0;
assign v$P$AD_963_out0 = v$G1_5976_out0;
assign v$P$AD_975_out0 = v$G1_5988_out0;
assign v$P$AD_977_out0 = v$G1_5990_out0;
assign v$P$AD_980_out0 = v$G1_5993_out0;
assign v$P$AD_986_out0 = v$G1_5999_out0;
assign v$P$AD_991_out0 = v$G1_6004_out0;
assign {v$A2A_1790_out1,v$A2A_1790_out0 } = v$A1_1871_out0 + v$B1_8428_out0 + v$C0_11190_out0;
assign {v$A2A_1793_out1,v$A2A_1793_out0 } = v$A1_1874_out0 + v$B1_8431_out0 + v$C0_11193_out0;
assign v$XOR2_8172_out0 = v$MUX1_14796_out0 ^ v$MUX3_3953_out0;
assign v$XOR2_8173_out0 = v$MUX1_14797_out0 ^ v$MUX3_3954_out0;
assign v$C0_9747_out0 = v$C0_11190_out0;
assign v$C0_9750_out0 = v$C0_11193_out0;
assign v$G4_11696_out0 = v$G5_4775_out0 || v$G$CD_1103_out0;
assign v$G4_11699_out0 = v$G5_4778_out0 || v$G$CD_1106_out0;
assign v$G4_11700_out0 = v$G5_4779_out0 || v$G$CD_1107_out0;
assign v$G4_11712_out0 = v$G5_4791_out0 || v$G$CD_1119_out0;
assign v$G4_11714_out0 = v$G5_4793_out0 || v$G$CD_1121_out0;
assign v$G4_11717_out0 = v$G5_4796_out0 || v$G$CD_1124_out0;
assign v$G4_11723_out0 = v$G5_4802_out0 || v$G$CD_1130_out0;
assign v$G4_11728_out0 = v$G5_4807_out0 || v$G$CD_1135_out0;
assign v$G4_11819_out0 = v$G5_4898_out0 || v$G$CD_1226_out0;
assign v$G4_11822_out0 = v$G5_4901_out0 || v$G$CD_1229_out0;
assign v$G4_11823_out0 = v$G5_4902_out0 || v$G$CD_1230_out0;
assign v$G4_11835_out0 = v$G5_4914_out0 || v$G$CD_1242_out0;
assign v$G4_11837_out0 = v$G5_4916_out0 || v$G$CD_1244_out0;
assign v$G4_11840_out0 = v$G5_4919_out0 || v$G$CD_1247_out0;
assign v$G4_11846_out0 = v$G5_4925_out0 || v$G$CD_1253_out0;
assign v$G4_11851_out0 = v$G5_4930_out0 || v$G$CD_1258_out0;
assign v$A1_14171_out0 = v$MUX4_6167_out0;
assign v$A1_14174_out0 = v$MUX4_6168_out0;
assign v$G6_538_out0 = v$G4_11696_out0 || v$G7_10103_out0;
assign v$G6_541_out0 = v$G4_11699_out0 || v$G7_10106_out0;
assign v$G6_542_out0 = v$G4_11700_out0 || v$G7_10107_out0;
assign v$G6_554_out0 = v$G4_11712_out0 || v$G7_10119_out0;
assign v$G6_556_out0 = v$G4_11714_out0 || v$G7_10121_out0;
assign v$G6_559_out0 = v$G4_11717_out0 || v$G7_10124_out0;
assign v$G6_565_out0 = v$G4_11723_out0 || v$G7_10130_out0;
assign v$G6_570_out0 = v$G4_11728_out0 || v$G7_10135_out0;
assign v$G6_661_out0 = v$G4_11819_out0 || v$G7_10226_out0;
assign v$G6_664_out0 = v$G4_11822_out0 || v$G7_10229_out0;
assign v$G6_665_out0 = v$G4_11823_out0 || v$G7_10230_out0;
assign v$G6_677_out0 = v$G4_11835_out0 || v$G7_10242_out0;
assign v$G6_679_out0 = v$G4_11837_out0 || v$G7_10244_out0;
assign v$G6_682_out0 = v$G4_11840_out0 || v$G7_10247_out0;
assign v$G6_688_out0 = v$G4_11846_out0 || v$G7_10253_out0;
assign v$G6_693_out0 = v$G4_11851_out0 || v$G7_10258_out0;
assign v$END1_1699_out0 = v$A2A_1790_out1;
assign v$END1_1702_out0 = v$A2A_1793_out1;
assign v$P$AB_2247_out0 = v$P$AD_852_out0;
assign v$P$AB_2248_out0 = v$P$AD_857_out0;
assign v$P$AB_2261_out0 = v$P$AD_840_out0;
assign v$P$AB_2263_out0 = v$P$AD_836_out0;
assign v$P$AB_2264_out0 = v$P$AD_863_out0;
assign v$P$AB_2267_out0 = v$P$AD_854_out0;
assign v$P$AB_2281_out0 = v$P$AD_839_out0;
assign v$P$AB_2286_out0 = v$P$AD_868_out0;
assign v$P$AB_2370_out0 = v$P$AD_975_out0;
assign v$P$AB_2371_out0 = v$P$AD_980_out0;
assign v$P$AB_2384_out0 = v$P$AD_963_out0;
assign v$P$AB_2386_out0 = v$P$AD_959_out0;
assign v$P$AB_2387_out0 = v$P$AD_986_out0;
assign v$P$AB_2390_out0 = v$P$AD_977_out0;
assign v$P$AB_2404_out0 = v$P$AD_962_out0;
assign v$P$AB_2409_out0 = v$P$AD_991_out0;
assign v$_7861_out0 = v$A1_14171_out0[11:0];
assign v$_7861_out1 = v$A1_14171_out0[23:12];
assign v$_7864_out0 = v$A1_14174_out0[11:0];
assign v$_7864_out1 = v$A1_14174_out0[23:12];
assign v$B2_8721_out0 = v$XOR2_8172_out0;
assign v$B2_8724_out0 = v$XOR2_8173_out0;
assign v$P$CD_10993_out0 = v$P$AD_863_out0;
assign v$P$CD_10997_out0 = v$P$AD_840_out0;
assign v$P$CD_11018_out0 = v$P$AD_854_out0;
assign v$P$CD_11021_out0 = v$P$AD_852_out0;
assign v$P$CD_11022_out0 = v$P$AD_868_out0;
assign v$P$CD_11026_out0 = v$P$AD_839_out0;
assign v$P$CD_11027_out0 = v$P$AD_857_out0;
assign v$P$CD_11116_out0 = v$P$AD_986_out0;
assign v$P$CD_11120_out0 = v$P$AD_963_out0;
assign v$P$CD_11141_out0 = v$P$AD_977_out0;
assign v$P$CD_11144_out0 = v$P$AD_975_out0;
assign v$P$CD_11145_out0 = v$P$AD_991_out0;
assign v$P$CD_11149_out0 = v$P$AD_962_out0;
assign v$P$CD_11150_out0 = v$P$AD_980_out0;
assign v$_14023_out0 = { v$A1A_12226_out0,v$A2A_1790_out0 };
assign v$_14026_out0 = { v$A1A_12229_out0,v$A2A_1793_out0 };
assign v$G$AD_17770_out0 = v$G4_11696_out0;
assign v$G$AD_17773_out0 = v$G4_11699_out0;
assign v$G$AD_17774_out0 = v$G4_11700_out0;
assign v$G$AD_17786_out0 = v$G4_11712_out0;
assign v$G$AD_17788_out0 = v$G4_11714_out0;
assign v$G$AD_17791_out0 = v$G4_11717_out0;
assign v$G$AD_17797_out0 = v$G4_11723_out0;
assign v$G$AD_17802_out0 = v$G4_11728_out0;
assign v$G$AD_17893_out0 = v$G4_11819_out0;
assign v$G$AD_17896_out0 = v$G4_11822_out0;
assign v$G$AD_17897_out0 = v$G4_11823_out0;
assign v$G$AD_17909_out0 = v$G4_11835_out0;
assign v$G$AD_17911_out0 = v$G4_11837_out0;
assign v$G$AD_17914_out0 = v$G4_11840_out0;
assign v$G$AD_17920_out0 = v$G4_11846_out0;
assign v$G$AD_17925_out0 = v$G4_11851_out0;
assign v$G$CD_1104_out0 = v$G$AD_17797_out0;
assign v$G$CD_1108_out0 = v$G$AD_17774_out0;
assign v$G$CD_1129_out0 = v$G$AD_17788_out0;
assign v$G$CD_1132_out0 = v$G$AD_17786_out0;
assign v$G$CD_1133_out0 = v$G$AD_17802_out0;
assign v$G$CD_1137_out0 = v$G$AD_17773_out0;
assign v$G$CD_1138_out0 = v$G$AD_17791_out0;
assign v$G$CD_1227_out0 = v$G$AD_17920_out0;
assign v$G$CD_1231_out0 = v$G$AD_17897_out0;
assign v$G$CD_1252_out0 = v$G$AD_17911_out0;
assign v$G$CD_1255_out0 = v$G$AD_17909_out0;
assign v$G$CD_1256_out0 = v$G$AD_17925_out0;
assign v$G$CD_1260_out0 = v$G$AD_17896_out0;
assign v$G$CD_1261_out0 = v$G$AD_17914_out0;
assign v$_4141_out0 = v$B2_8721_out0[11:0];
assign v$_4141_out1 = v$B2_8721_out0[23:12];
assign v$_4144_out0 = v$B2_8724_out0[11:0];
assign v$_4144_out1 = v$B2_8724_out0[23:12];
assign v$G1_5846_out0 = v$P$AB_2247_out0 && v$P$CD_10989_out0;
assign v$G1_5847_out0 = v$P$AB_2248_out0 && v$P$CD_10990_out0;
assign v$G1_5860_out0 = v$P$AB_2261_out0 && v$P$CD_11003_out0;
assign v$G1_5862_out0 = v$P$AB_2263_out0 && v$P$CD_11005_out0;
assign v$G1_5863_out0 = v$P$AB_2264_out0 && v$P$CD_11006_out0;
assign v$G1_5866_out0 = v$P$AB_2267_out0 && v$P$CD_11009_out0;
assign v$G1_5880_out0 = v$P$AB_2281_out0 && v$P$CD_11023_out0;
assign v$G1_5885_out0 = v$P$AB_2286_out0 && v$P$CD_11028_out0;
assign v$G1_5969_out0 = v$P$AB_2370_out0 && v$P$CD_11112_out0;
assign v$G1_5970_out0 = v$P$AB_2371_out0 && v$P$CD_11113_out0;
assign v$G1_5983_out0 = v$P$AB_2384_out0 && v$P$CD_11126_out0;
assign v$G1_5985_out0 = v$P$AB_2386_out0 && v$P$CD_11128_out0;
assign v$G1_5986_out0 = v$P$AB_2387_out0 && v$P$CD_11129_out0;
assign v$G1_5989_out0 = v$P$AB_2390_out0 && v$P$CD_11132_out0;
assign v$G1_6003_out0 = v$P$AB_2404_out0 && v$P$CD_11146_out0;
assign v$G1_6008_out0 = v$P$AB_2409_out0 && v$P$CD_11151_out0;
assign v$COUTD_7016_out0 = v$G6_538_out0;
assign v$COUTD_7019_out0 = v$G6_541_out0;
assign v$COUTD_7020_out0 = v$G6_542_out0;
assign v$COUTD_7032_out0 = v$G6_554_out0;
assign v$COUTD_7034_out0 = v$G6_556_out0;
assign v$COUTD_7037_out0 = v$G6_559_out0;
assign v$COUTD_7043_out0 = v$G6_565_out0;
assign v$COUTD_7048_out0 = v$G6_570_out0;
assign v$COUTD_7139_out0 = v$G6_661_out0;
assign v$COUTD_7142_out0 = v$G6_664_out0;
assign v$COUTD_7143_out0 = v$G6_665_out0;
assign v$COUTD_7155_out0 = v$G6_677_out0;
assign v$COUTD_7157_out0 = v$G6_679_out0;
assign v$COUTD_7160_out0 = v$G6_682_out0;
assign v$COUTD_7166_out0 = v$G6_688_out0;
assign v$COUTD_7171_out0 = v$G6_693_out0;
assign v$G$AB_9547_out0 = v$G$AD_17786_out0;
assign v$G$AB_9548_out0 = v$G$AD_17791_out0;
assign v$G$AB_9561_out0 = v$G$AD_17774_out0;
assign v$G$AB_9563_out0 = v$G$AD_17770_out0;
assign v$G$AB_9564_out0 = v$G$AD_17797_out0;
assign v$G$AB_9567_out0 = v$G$AD_17788_out0;
assign v$G$AB_9581_out0 = v$G$AD_17773_out0;
assign v$G$AB_9586_out0 = v$G$AD_17802_out0;
assign v$G$AB_9670_out0 = v$G$AD_17909_out0;
assign v$G$AB_9671_out0 = v$G$AD_17914_out0;
assign v$G$AB_9684_out0 = v$G$AD_17897_out0;
assign v$G$AB_9686_out0 = v$G$AD_17893_out0;
assign v$G$AB_9687_out0 = v$G$AD_17920_out0;
assign v$G$AB_9690_out0 = v$G$AD_17911_out0;
assign v$G$AB_9704_out0 = v$G$AD_17896_out0;
assign v$G$AB_9709_out0 = v$G$AD_17925_out0;
assign v$_16724_out0 = v$_7861_out0[5:0];
assign v$_16724_out1 = v$_7861_out0[11:6];
assign v$_16727_out0 = v$_7864_out0[5:0];
assign v$_16727_out1 = v$_7864_out0[11:6];
assign v$_17623_out0 = v$_7861_out1[5:0];
assign v$_17623_out1 = v$_7861_out1[11:6];
assign v$_17626_out0 = v$_7864_out1[5:0];
assign v$_17626_out1 = v$_7864_out1[11:6];
assign v$P$AD_833_out0 = v$G1_5846_out0;
assign v$P$AD_834_out0 = v$G1_5847_out0;
assign v$P$AD_847_out0 = v$G1_5860_out0;
assign v$P$AD_849_out0 = v$G1_5862_out0;
assign v$P$AD_850_out0 = v$G1_5863_out0;
assign v$P$AD_853_out0 = v$G1_5866_out0;
assign v$P$AD_867_out0 = v$G1_5880_out0;
assign v$P$AD_872_out0 = v$G1_5885_out0;
assign v$P$AD_956_out0 = v$G1_5969_out0;
assign v$P$AD_957_out0 = v$G1_5970_out0;
assign v$P$AD_970_out0 = v$G1_5983_out0;
assign v$P$AD_972_out0 = v$G1_5985_out0;
assign v$P$AD_973_out0 = v$G1_5986_out0;
assign v$P$AD_976_out0 = v$G1_5989_out0;
assign v$P$AD_990_out0 = v$G1_6003_out0;
assign v$P$AD_995_out0 = v$G1_6008_out0;
assign v$_1370_out0 = v$_4141_out1[5:0];
assign v$_1370_out1 = v$_4141_out1[11:6];
assign v$_1373_out0 = v$_4144_out1[5:0];
assign v$_1373_out1 = v$_4144_out1[11:6];
assign v$_1678_out0 = v$_4141_out0[5:0];
assign v$_1678_out1 = v$_4141_out0[11:6];
assign v$_1681_out0 = v$_4144_out0[5:0];
assign v$_1681_out1 = v$_4144_out0[11:6];
assign v$_2025_out0 = v$_17623_out1[2:0];
assign v$_2025_out1 = v$_17623_out1[5:3];
assign v$_2028_out0 = v$_17626_out1[2:0];
assign v$_2028_out1 = v$_17626_out1[5:3];
assign v$G5_4772_out0 = v$G$AB_9547_out0 && v$P$CD_10989_out0;
assign v$G5_4773_out0 = v$G$AB_9548_out0 && v$P$CD_10990_out0;
assign v$G5_4786_out0 = v$G$AB_9561_out0 && v$P$CD_11003_out0;
assign v$G5_4788_out0 = v$G$AB_9563_out0 && v$P$CD_11005_out0;
assign v$G5_4789_out0 = v$G$AB_9564_out0 && v$P$CD_11006_out0;
assign v$G5_4792_out0 = v$G$AB_9567_out0 && v$P$CD_11009_out0;
assign v$G5_4806_out0 = v$G$AB_9581_out0 && v$P$CD_11023_out0;
assign v$G5_4811_out0 = v$G$AB_9586_out0 && v$P$CD_11028_out0;
assign v$G5_4895_out0 = v$G$AB_9670_out0 && v$P$CD_11112_out0;
assign v$G5_4896_out0 = v$G$AB_9671_out0 && v$P$CD_11113_out0;
assign v$G5_4909_out0 = v$G$AB_9684_out0 && v$P$CD_11126_out0;
assign v$G5_4911_out0 = v$G$AB_9686_out0 && v$P$CD_11128_out0;
assign v$G5_4912_out0 = v$G$AB_9687_out0 && v$P$CD_11129_out0;
assign v$G5_4915_out0 = v$G$AB_9690_out0 && v$P$CD_11132_out0;
assign v$G5_4929_out0 = v$G$AB_9704_out0 && v$P$CD_11146_out0;
assign v$G5_4934_out0 = v$G$AB_9709_out0 && v$P$CD_11151_out0;
assign v$CINA_8853_out0 = v$COUTD_7032_out0;
assign v$CINA_8854_out0 = v$COUTD_7037_out0;
assign v$CINA_8867_out0 = v$COUTD_7020_out0;
assign v$CINA_8869_out0 = v$COUTD_7016_out0;
assign v$CINA_8870_out0 = v$COUTD_7043_out0;
assign v$CINA_8873_out0 = v$COUTD_7034_out0;
assign v$CINA_8887_out0 = v$COUTD_7019_out0;
assign v$CINA_8892_out0 = v$COUTD_7048_out0;
assign v$CINA_8976_out0 = v$COUTD_7155_out0;
assign v$CINA_8977_out0 = v$COUTD_7160_out0;
assign v$CINA_8990_out0 = v$COUTD_7143_out0;
assign v$CINA_8992_out0 = v$COUTD_7139_out0;
assign v$CINA_8993_out0 = v$COUTD_7166_out0;
assign v$CINA_8996_out0 = v$COUTD_7157_out0;
assign v$CINA_9010_out0 = v$COUTD_7142_out0;
assign v$CINA_9015_out0 = v$COUTD_7171_out0;
assign v$_10475_out0 = v$_17623_out0[2:0];
assign v$_10475_out1 = v$_17623_out0[5:3];
assign v$_10478_out0 = v$_17626_out0[2:0];
assign v$_10478_out1 = v$_17626_out0[5:3];
assign v$_14356_out0 = v$_16724_out0[2:0];
assign v$_14356_out1 = v$_16724_out0[5:3];
assign v$_14359_out0 = v$_16727_out0[2:0];
assign v$_14359_out1 = v$_16727_out0[5:3];
assign v$C1_17403_out0 = v$COUTD_7016_out0;
assign v$C1_17406_out0 = v$COUTD_7139_out0;
assign v$_19028_out0 = v$_16724_out1[2:0];
assign v$_19028_out1 = v$_16724_out1[5:3];
assign v$_19031_out0 = v$_16727_out1[2:0];
assign v$_19031_out1 = v$_16727_out1[5:3];
assign v$_1463_out0 = v$_19028_out0[0:0];
assign v$_1463_out1 = v$_19028_out0[2:2];
assign v$_1466_out0 = v$_19031_out0[0:0];
assign v$_1466_out1 = v$_19031_out0[2:2];
assign v$_1516_out0 = v$_14356_out1[0:0];
assign v$_1516_out1 = v$_14356_out1[2:2];
assign v$_1519_out0 = v$_14359_out1[0:0];
assign v$_1519_out1 = v$_14359_out1[2:2];
assign v$_2015_out0 = v$_2025_out1[0:0];
assign v$_2015_out1 = v$_2025_out1[2:2];
assign v$_2018_out0 = v$_2028_out1[0:0];
assign v$_2018_out1 = v$_2028_out1[2:2];
assign v$P$AB_2246_out0 = v$P$AD_834_out0;
assign v$P$AB_2251_out0 = v$P$AD_849_out0;
assign v$P$AB_2257_out0 = v$P$AD_849_out0;
assign v$P$AB_2260_out0 = v$P$AD_867_out0;
assign v$P$AB_2265_out0 = v$P$AD_833_out0;
assign v$P$AB_2278_out0 = v$P$AD_849_out0;
assign v$P$AB_2369_out0 = v$P$AD_957_out0;
assign v$P$AB_2374_out0 = v$P$AD_972_out0;
assign v$P$AB_2380_out0 = v$P$AD_972_out0;
assign v$P$AB_2383_out0 = v$P$AD_990_out0;
assign v$P$AB_2388_out0 = v$P$AD_956_out0;
assign v$P$AB_2401_out0 = v$P$AD_972_out0;
assign v$_7356_out0 = v$_14356_out0[0:0];
assign v$_7356_out1 = v$_14356_out0[2:2];
assign v$_7359_out0 = v$_14359_out0[0:0];
assign v$_7359_out1 = v$_14359_out0[2:2];
assign v$_10357_out0 = v$_1370_out1[2:0];
assign v$_10357_out1 = v$_1370_out1[5:3];
assign v$_10360_out0 = v$_1373_out1[2:0];
assign v$_10360_out1 = v$_1373_out1[5:3];
assign v$_10899_out0 = v$_10475_out0[0:0];
assign v$_10899_out1 = v$_10475_out0[2:2];
assign v$_10902_out0 = v$_10478_out0[0:0];
assign v$_10902_out1 = v$_10478_out0[2:2];
assign v$P$CD_10988_out0 = v$P$AD_872_out0;
assign v$P$CD_10994_out0 = v$P$AD_834_out0;
assign v$P$CD_11002_out0 = v$P$AD_847_out0;
assign v$P$CD_11007_out0 = v$P$AD_853_out0;
assign v$P$CD_11011_out0 = v$P$AD_867_out0;
assign v$P$CD_11012_out0 = v$P$AD_833_out0;
assign v$P$CD_11020_out0 = v$P$AD_850_out0;
assign v$P$CD_11111_out0 = v$P$AD_995_out0;
assign v$P$CD_11117_out0 = v$P$AD_957_out0;
assign v$P$CD_11125_out0 = v$P$AD_970_out0;
assign v$P$CD_11130_out0 = v$P$AD_976_out0;
assign v$P$CD_11134_out0 = v$P$AD_990_out0;
assign v$P$CD_11135_out0 = v$P$AD_956_out0;
assign v$P$CD_11143_out0 = v$P$AD_973_out0;
assign v$_11414_out0 = v$_19028_out1[0:0];
assign v$_11414_out1 = v$_19028_out1[2:2];
assign v$_11417_out0 = v$_19031_out1[0:0];
assign v$_11417_out1 = v$_19031_out1[2:2];
assign v$_11597_out0 = v$_2025_out0[0:0];
assign v$_11597_out1 = v$_2025_out0[2:2];
assign v$_11600_out0 = v$_2028_out0[0:0];
assign v$_11600_out1 = v$_2028_out0[2:2];
assign v$G4_11693_out0 = v$G5_4772_out0 || v$G$CD_1100_out0;
assign v$G4_11694_out0 = v$G5_4773_out0 || v$G$CD_1101_out0;
assign v$G4_11707_out0 = v$G5_4786_out0 || v$G$CD_1114_out0;
assign v$G4_11709_out0 = v$G5_4788_out0 || v$G$CD_1116_out0;
assign v$G4_11710_out0 = v$G5_4789_out0 || v$G$CD_1117_out0;
assign v$G4_11713_out0 = v$G5_4792_out0 || v$G$CD_1120_out0;
assign v$G4_11727_out0 = v$G5_4806_out0 || v$G$CD_1134_out0;
assign v$G4_11732_out0 = v$G5_4811_out0 || v$G$CD_1139_out0;
assign v$G4_11816_out0 = v$G5_4895_out0 || v$G$CD_1223_out0;
assign v$G4_11817_out0 = v$G5_4896_out0 || v$G$CD_1224_out0;
assign v$G4_11830_out0 = v$G5_4909_out0 || v$G$CD_1237_out0;
assign v$G4_11832_out0 = v$G5_4911_out0 || v$G$CD_1239_out0;
assign v$G4_11833_out0 = v$G5_4912_out0 || v$G$CD_1240_out0;
assign v$G4_11836_out0 = v$G5_4915_out0 || v$G$CD_1243_out0;
assign v$G4_11850_out0 = v$G5_4929_out0 || v$G$CD_1257_out0;
assign v$G4_11855_out0 = v$G5_4934_out0 || v$G$CD_1262_out0;
assign v$G8_12008_out0 = v$CINA_8853_out0 && v$P$AB_2247_out0;
assign v$G8_12009_out0 = v$CINA_8854_out0 && v$P$AB_2248_out0;
assign v$G8_12022_out0 = v$CINA_8867_out0 && v$P$AB_2261_out0;
assign v$G8_12024_out0 = v$CINA_8869_out0 && v$P$AB_2263_out0;
assign v$G8_12025_out0 = v$CINA_8870_out0 && v$P$AB_2264_out0;
assign v$G8_12028_out0 = v$CINA_8873_out0 && v$P$AB_2267_out0;
assign v$G8_12042_out0 = v$CINA_8887_out0 && v$P$AB_2281_out0;
assign v$G8_12047_out0 = v$CINA_8892_out0 && v$P$AB_2286_out0;
assign v$G8_12131_out0 = v$CINA_8976_out0 && v$P$AB_2370_out0;
assign v$G8_12132_out0 = v$CINA_8977_out0 && v$P$AB_2371_out0;
assign v$G8_12145_out0 = v$CINA_8990_out0 && v$P$AB_2384_out0;
assign v$G8_12147_out0 = v$CINA_8992_out0 && v$P$AB_2386_out0;
assign v$G8_12148_out0 = v$CINA_8993_out0 && v$P$AB_2387_out0;
assign v$G8_12151_out0 = v$CINA_8996_out0 && v$P$AB_2390_out0;
assign v$G8_12165_out0 = v$CINA_9010_out0 && v$P$AB_2404_out0;
assign v$G8_12170_out0 = v$CINA_9015_out0 && v$P$AB_2409_out0;
assign v$C1_12423_out0 = v$C1_17403_out0;
assign v$C1_12426_out0 = v$C1_17406_out0;
assign {v$A3A_12527_out1,v$A3A_12527_out0 } = v$A2_18870_out0 + v$B2_3328_out0 + v$C1_17403_out0;
assign {v$A3A_12530_out1,v$A3A_12530_out0 } = v$A2_18873_out0 + v$B2_3331_out0 + v$C1_17406_out0;
assign v$_13562_out0 = v$_1678_out1[2:0];
assign v$_13562_out1 = v$_1678_out1[5:3];
assign v$_13565_out0 = v$_1681_out1[2:0];
assign v$_13565_out1 = v$_1681_out1[5:3];
assign v$_14325_out0 = v$_1678_out0[2:0];
assign v$_14325_out1 = v$_1678_out0[5:3];
assign v$_14328_out0 = v$_1681_out0[2:0];
assign v$_14328_out1 = v$_1681_out0[5:3];
assign v$_16743_out0 = v$_10475_out1[0:0];
assign v$_16743_out1 = v$_10475_out1[2:2];
assign v$_16746_out0 = v$_10478_out1[0:0];
assign v$_16746_out1 = v$_10478_out1[2:2];
assign v$_18341_out0 = v$_1370_out0[2:0];
assign v$_18341_out1 = v$_1370_out0[5:3];
assign v$_18344_out0 = v$_1373_out0[2:0];
assign v$_18344_out1 = v$_1373_out0[5:3];
assign v$A6_321_out0 = v$_1463_out0;
assign v$A6_324_out0 = v$_1466_out0;
assign v$A21_2793_out0 = v$_2015_out0;
assign v$A21_2796_out0 = v$_2018_out0;
assign v$_3130_out0 = v$_14325_out0[0:0];
assign v$_3130_out1 = v$_14325_out0[2:2];
assign v$_3133_out0 = v$_14328_out0[0:0];
assign v$_3133_out1 = v$_14328_out0[2:2];
assign v$A12_3356_out0 = v$_10899_out0;
assign v$A12_3359_out0 = v$_10902_out0;
assign v$A9_3644_out0 = v$_11414_out0;
assign v$A9_3647_out0 = v$_11417_out0;
assign v$A0_4469_out0 = v$_7356_out0;
assign v$A0_4472_out0 = v$_7359_out0;
assign v$END2_5451_out0 = v$A3A_12527_out1;
assign v$END2_5454_out0 = v$A3A_12530_out1;
assign v$G1_5845_out0 = v$P$AB_2246_out0 && v$P$CD_10988_out0;
assign v$G1_5850_out0 = v$P$AB_2251_out0 && v$P$CD_10993_out0;
assign v$G1_5856_out0 = v$P$AB_2257_out0 && v$P$CD_10999_out0;
assign v$G1_5859_out0 = v$P$AB_2260_out0 && v$P$CD_11002_out0;
assign v$G1_5864_out0 = v$P$AB_2265_out0 && v$P$CD_11007_out0;
assign v$G1_5877_out0 = v$P$AB_2278_out0 && v$P$CD_11020_out0;
assign v$G1_5968_out0 = v$P$AB_2369_out0 && v$P$CD_11111_out0;
assign v$G1_5973_out0 = v$P$AB_2374_out0 && v$P$CD_11116_out0;
assign v$G1_5979_out0 = v$P$AB_2380_out0 && v$P$CD_11122_out0;
assign v$G1_5982_out0 = v$P$AB_2383_out0 && v$P$CD_11125_out0;
assign v$G1_5987_out0 = v$P$AB_2388_out0 && v$P$CD_11130_out0;
assign v$G1_6000_out0 = v$P$AB_2401_out0 && v$P$CD_11143_out0;
assign v$_6229_out0 = v$_16743_out1[0:0];
assign v$_6229_out1 = v$_16743_out1[1:1];
assign v$_6232_out0 = v$_16746_out1[0:0];
assign v$_6232_out1 = v$_16746_out1[1:1];
assign v$_7677_out0 = v$_1516_out1[0:0];
assign v$_7677_out1 = v$_1516_out1[1:1];
assign v$_7680_out0 = v$_1519_out1[0:0];
assign v$_7680_out1 = v$_1519_out1[1:1];
assign v$_8089_out0 = v$_18341_out0[0:0];
assign v$_8089_out1 = v$_18341_out0[2:2];
assign v$_8092_out0 = v$_18344_out0[0:0];
assign v$_8092_out1 = v$_18344_out0[2:2];
assign v$_9237_out0 = { v$C0_9747_out0,v$C1_12423_out0 };
assign v$_9240_out0 = { v$C0_9750_out0,v$C1_12426_out0 };
assign v$_9390_out0 = v$_10357_out1[0:0];
assign v$_9390_out1 = v$_10357_out1[2:2];
assign v$_9393_out0 = v$_10360_out1[0:0];
assign v$_9393_out1 = v$_10360_out1[2:2];
assign v$G7_10100_out0 = v$G8_12008_out0 && v$P$CD_10989_out0;
assign v$G7_10101_out0 = v$G8_12009_out0 && v$P$CD_10990_out0;
assign v$G7_10114_out0 = v$G8_12022_out0 && v$P$CD_11003_out0;
assign v$G7_10116_out0 = v$G8_12024_out0 && v$P$CD_11005_out0;
assign v$G7_10117_out0 = v$G8_12025_out0 && v$P$CD_11006_out0;
assign v$G7_10120_out0 = v$G8_12028_out0 && v$P$CD_11009_out0;
assign v$G7_10134_out0 = v$G8_12042_out0 && v$P$CD_11023_out0;
assign v$G7_10139_out0 = v$G8_12047_out0 && v$P$CD_11028_out0;
assign v$G7_10223_out0 = v$G8_12131_out0 && v$P$CD_11112_out0;
assign v$G7_10224_out0 = v$G8_12132_out0 && v$P$CD_11113_out0;
assign v$G7_10237_out0 = v$G8_12145_out0 && v$P$CD_11126_out0;
assign v$G7_10239_out0 = v$G8_12147_out0 && v$P$CD_11128_out0;
assign v$G7_10240_out0 = v$G8_12148_out0 && v$P$CD_11129_out0;
assign v$G7_10243_out0 = v$G8_12151_out0 && v$P$CD_11132_out0;
assign v$G7_10257_out0 = v$G8_12165_out0 && v$P$CD_11146_out0;
assign v$G7_10262_out0 = v$G8_12170_out0 && v$P$CD_11151_out0;
assign v$_10740_out0 = v$_2015_out1[0:0];
assign v$_10740_out1 = v$_2015_out1[1:1];
assign v$_10743_out0 = v$_2018_out1[0:0];
assign v$_10743_out1 = v$_2018_out1[1:1];
assign v$_11265_out0 = v$_13562_out1[0:0];
assign v$_11265_out1 = v$_13562_out1[2:2];
assign v$_11268_out0 = v$_13565_out1[0:0];
assign v$_11268_out1 = v$_13565_out1[2:2];
assign v$_12179_out0 = v$_7356_out1[0:0];
assign v$_12179_out1 = v$_7356_out1[1:1];
assign v$_12182_out0 = v$_7359_out1[0:0];
assign v$_12182_out1 = v$_7359_out1[1:1];
assign v$A3_15210_out0 = v$_1516_out0;
assign v$A3_15213_out0 = v$_1519_out0;
assign v$_15759_out0 = v$_10357_out0[0:0];
assign v$_15759_out1 = v$_10357_out0[2:2];
assign v$_15762_out0 = v$_10360_out0[0:0];
assign v$_15762_out1 = v$_10360_out0[2:2];
assign v$_16340_out0 = v$_1463_out1[0:0];
assign v$_16340_out1 = v$_1463_out1[1:1];
assign v$_16343_out0 = v$_1466_out1[0:0];
assign v$_16343_out1 = v$_1466_out1[1:1];
assign v$_16792_out0 = v$_10899_out1[0:0];
assign v$_16792_out1 = v$_10899_out1[1:1];
assign v$_16795_out0 = v$_10902_out1[0:0];
assign v$_16795_out1 = v$_10902_out1[1:1];
assign v$_16877_out0 = v$_18341_out1[0:0];
assign v$_16877_out1 = v$_18341_out1[2:2];
assign v$_16880_out0 = v$_18344_out1[0:0];
assign v$_16880_out1 = v$_18344_out1[2:2];
assign v$_17323_out0 = v$_11597_out1[0:0];
assign v$_17323_out1 = v$_11597_out1[1:1];
assign v$_17326_out0 = v$_11600_out1[0:0];
assign v$_17326_out1 = v$_11600_out1[1:1];
assign v$_17362_out0 = v$_14325_out1[0:0];
assign v$_17362_out1 = v$_14325_out1[2:2];
assign v$_17365_out0 = v$_14328_out1[0:0];
assign v$_17365_out1 = v$_14328_out1[2:2];
assign v$G$AD_17767_out0 = v$G4_11693_out0;
assign v$G$AD_17768_out0 = v$G4_11694_out0;
assign v$G$AD_17781_out0 = v$G4_11707_out0;
assign v$G$AD_17783_out0 = v$G4_11709_out0;
assign v$G$AD_17784_out0 = v$G4_11710_out0;
assign v$G$AD_17787_out0 = v$G4_11713_out0;
assign v$G$AD_17801_out0 = v$G4_11727_out0;
assign v$G$AD_17806_out0 = v$G4_11732_out0;
assign v$G$AD_17890_out0 = v$G4_11816_out0;
assign v$G$AD_17891_out0 = v$G4_11817_out0;
assign v$G$AD_17904_out0 = v$G4_11830_out0;
assign v$G$AD_17906_out0 = v$G4_11832_out0;
assign v$G$AD_17907_out0 = v$G4_11833_out0;
assign v$G$AD_17910_out0 = v$G4_11836_out0;
assign v$G$AD_17924_out0 = v$G4_11850_out0;
assign v$G$AD_17929_out0 = v$G4_11855_out0;
assign v$A15_17958_out0 = v$_16743_out0;
assign v$A15_17961_out0 = v$_16746_out0;
assign v$A18_18301_out0 = v$_11597_out0;
assign v$A18_18304_out0 = v$_11600_out0;
assign v$_18367_out0 = v$_11414_out1[0:0];
assign v$_18367_out1 = v$_11414_out1[1:1];
assign v$_18370_out0 = v$_11417_out1[0:0];
assign v$_18370_out1 = v$_11417_out1[1:1];
assign v$_18788_out0 = v$_13562_out0[0:0];
assign v$_18788_out1 = v$_13562_out0[2:2];
assign v$_18791_out0 = v$_13565_out0[0:0];
assign v$_18791_out1 = v$_13565_out0[2:2];
assign v$G6_535_out0 = v$G4_11693_out0 || v$G7_10100_out0;
assign v$G6_536_out0 = v$G4_11694_out0 || v$G7_10101_out0;
assign v$G6_549_out0 = v$G4_11707_out0 || v$G7_10114_out0;
assign v$G6_551_out0 = v$G4_11709_out0 || v$G7_10116_out0;
assign v$G6_552_out0 = v$G4_11710_out0 || v$G7_10117_out0;
assign v$G6_555_out0 = v$G4_11713_out0 || v$G7_10120_out0;
assign v$G6_569_out0 = v$G4_11727_out0 || v$G7_10134_out0;
assign v$G6_574_out0 = v$G4_11732_out0 || v$G7_10139_out0;
assign v$G6_658_out0 = v$G4_11816_out0 || v$G7_10223_out0;
assign v$G6_659_out0 = v$G4_11817_out0 || v$G7_10224_out0;
assign v$G6_672_out0 = v$G4_11830_out0 || v$G7_10237_out0;
assign v$G6_674_out0 = v$G4_11832_out0 || v$G7_10239_out0;
assign v$G6_675_out0 = v$G4_11833_out0 || v$G7_10240_out0;
assign v$G6_678_out0 = v$G4_11836_out0 || v$G7_10243_out0;
assign v$G6_692_out0 = v$G4_11850_out0 || v$G7_10257_out0;
assign v$G6_697_out0 = v$G4_11855_out0 || v$G7_10262_out0;
assign v$A14_739_out0 = v$_16792_out1;
assign v$A14_742_out0 = v$_16795_out1;
assign v$P$AD_832_out0 = v$G1_5845_out0;
assign v$P$AD_837_out0 = v$G1_5850_out0;
assign v$P$AD_843_out0 = v$G1_5856_out0;
assign v$P$AD_846_out0 = v$G1_5859_out0;
assign v$P$AD_851_out0 = v$G1_5864_out0;
assign v$P$AD_864_out0 = v$G1_5877_out0;
assign v$P$AD_955_out0 = v$G1_5968_out0;
assign v$P$AD_960_out0 = v$G1_5973_out0;
assign v$P$AD_966_out0 = v$G1_5979_out0;
assign v$P$AD_969_out0 = v$G1_5982_out0;
assign v$P$AD_974_out0 = v$G1_5987_out0;
assign v$P$AD_987_out0 = v$G1_6000_out0;
assign v$G$CD_1099_out0 = v$G$AD_17806_out0;
assign v$G$CD_1105_out0 = v$G$AD_17768_out0;
assign v$G$CD_1113_out0 = v$G$AD_17781_out0;
assign v$G$CD_1118_out0 = v$G$AD_17787_out0;
assign v$G$CD_1122_out0 = v$G$AD_17801_out0;
assign v$G$CD_1123_out0 = v$G$AD_17767_out0;
assign v$G$CD_1131_out0 = v$G$AD_17784_out0;
assign v$G$CD_1222_out0 = v$G$AD_17929_out0;
assign v$G$CD_1228_out0 = v$G$AD_17891_out0;
assign v$G$CD_1236_out0 = v$G$AD_17904_out0;
assign v$G$CD_1241_out0 = v$G$AD_17910_out0;
assign v$G$CD_1245_out0 = v$G$AD_17924_out0;
assign v$G$CD_1246_out0 = v$G$AD_17890_out0;
assign v$G$CD_1254_out0 = v$G$AD_17907_out0;
assign v$A19_1364_out0 = v$_17323_out0;
assign v$A19_1367_out0 = v$_17326_out0;
assign v$A10_1704_out0 = v$_18367_out0;
assign v$A10_1707_out0 = v$_18370_out0;
assign v$A1_1870_out0 = v$_12179_out0;
assign v$A1_1873_out0 = v$_12182_out0;
assign v$B12_2115_out0 = v$_8089_out0;
assign v$B12_2118_out0 = v$_8092_out0;
assign v$B0_3422_out0 = v$_3130_out0;
assign v$B0_3425_out0 = v$_3133_out0;
assign v$B9_4221_out0 = v$_11265_out0;
assign v$B9_4224_out0 = v$_11268_out0;
assign v$A22_4591_out0 = v$_10740_out0;
assign v$A22_4594_out0 = v$_10743_out0;
assign v$A20_4604_out0 = v$_17323_out1;
assign v$A20_4607_out0 = v$_17326_out1;
assign v$A23_5282_out0 = v$_10740_out1;
assign v$A23_5285_out0 = v$_10743_out1;
assign v$A5_6902_out0 = v$_7677_out1;
assign v$A5_6905_out0 = v$_7680_out1;
assign v$_7177_out0 = v$_18788_out1[0:0];
assign v$_7177_out1 = v$_18788_out1[1:1];
assign v$_7180_out0 = v$_18791_out1[0:0];
assign v$_7180_out1 = v$_18791_out1[1:1];
assign v$_7259_out0 = v$_17362_out1[0:0];
assign v$_7259_out1 = v$_17362_out1[1:1];
assign v$_7262_out0 = v$_17365_out1[0:0];
assign v$_7262_out1 = v$_17365_out1[1:1];
assign v$A_7415_out0 = v$A6_321_out0;
assign v$A_7416_out0 = v$A3_15210_out0;
assign v$A_7417_out0 = v$A21_2793_out0;
assign v$A_7418_out0 = v$A9_3644_out0;
assign v$A_7419_out0 = v$A15_17958_out0;
assign v$A_7423_out0 = v$A12_3356_out0;
assign v$A_7427_out0 = v$A0_4469_out0;
assign v$A_7432_out0 = v$A18_18301_out0;
assign v$A_7487_out0 = v$A6_324_out0;
assign v$A_7488_out0 = v$A3_15213_out0;
assign v$A_7489_out0 = v$A21_2796_out0;
assign v$A_7490_out0 = v$A9_3647_out0;
assign v$A_7491_out0 = v$A15_17961_out0;
assign v$A_7495_out0 = v$A12_3359_out0;
assign v$A_7499_out0 = v$A0_4472_out0;
assign v$A_7504_out0 = v$A18_18304_out0;
assign v$G$AB_9546_out0 = v$G$AD_17768_out0;
assign v$G$AB_9551_out0 = v$G$AD_17783_out0;
assign v$G$AB_9557_out0 = v$G$AD_17783_out0;
assign v$G$AB_9560_out0 = v$G$AD_17801_out0;
assign v$G$AB_9565_out0 = v$G$AD_17767_out0;
assign v$G$AB_9578_out0 = v$G$AD_17783_out0;
assign v$G$AB_9669_out0 = v$G$AD_17891_out0;
assign v$G$AB_9674_out0 = v$G$AD_17906_out0;
assign v$G$AB_9680_out0 = v$G$AD_17906_out0;
assign v$G$AB_9683_out0 = v$G$AD_17924_out0;
assign v$G$AB_9688_out0 = v$G$AD_17890_out0;
assign v$G$AB_9701_out0 = v$G$AD_17906_out0;
assign v$_9754_out0 = v$_9390_out1[0:0];
assign v$_9754_out1 = v$_9390_out1[1:1];
assign v$_9757_out0 = v$_9393_out1[0:0];
assign v$_9757_out1 = v$_9393_out1[1:1];
assign v$B3_9846_out0 = v$_17362_out0;
assign v$B3_9849_out0 = v$_17365_out0;
assign v$_9874_out0 = v$_11265_out1[0:0];
assign v$_9874_out1 = v$_11265_out1[1:1];
assign v$_9877_out0 = v$_11268_out1[0:0];
assign v$_9877_out1 = v$_11268_out1[1:1];
assign v$A11_10387_out0 = v$_18367_out1;
assign v$A11_10390_out0 = v$_18370_out1;
assign v$B15_10447_out0 = v$_16877_out0;
assign v$B15_10450_out0 = v$_16880_out0;
assign v$B18_11369_out0 = v$_15759_out0;
assign v$B18_11372_out0 = v$_15762_out0;
assign v$_11532_out0 = v$_3130_out1[0:0];
assign v$_11532_out1 = v$_3130_out1[1:1];
assign v$_11535_out0 = v$_3133_out1[0:0];
assign v$_11535_out1 = v$_3133_out1[1:1];
assign v$_13759_out0 = v$_16877_out1[0:0];
assign v$_13759_out1 = v$_16877_out1[1:1];
assign v$_13762_out0 = v$_16880_out1[0:0];
assign v$_13762_out1 = v$_16880_out1[1:1];
assign v$B6_13884_out0 = v$_18788_out0;
assign v$B6_13887_out0 = v$_18791_out0;
assign v$A16_14192_out0 = v$_6229_out0;
assign v$A16_14195_out0 = v$_6232_out0;
assign v$A13_14446_out0 = v$_16792_out0;
assign v$A13_14449_out0 = v$_16795_out0;
assign v$A7_15892_out0 = v$_16340_out0;
assign v$A7_15895_out0 = v$_16343_out0;
assign v$_17209_out0 = v$_15759_out1[0:0];
assign v$_17209_out1 = v$_15759_out1[1:1];
assign v$_17212_out0 = v$_15762_out1[0:0];
assign v$_17212_out1 = v$_15762_out1[1:1];
assign v$A17_17343_out0 = v$_6229_out1;
assign v$A17_17346_out0 = v$_6232_out1;
assign v$_17966_out0 = v$_8089_out1[0:0];
assign v$_17966_out1 = v$_8089_out1[1:1];
assign v$_17969_out0 = v$_8092_out1[0:0];
assign v$_17969_out1 = v$_8092_out1[1:1];
assign v$A4_18139_out0 = v$_7677_out0;
assign v$A4_18142_out0 = v$_7680_out0;
assign v$B21_18690_out0 = v$_9390_out0;
assign v$B21_18693_out0 = v$_9393_out0;
assign v$A8_18698_out0 = v$_16340_out1;
assign v$A8_18701_out0 = v$_16343_out1;
assign v$A2_18869_out0 = v$_12179_out1;
assign v$A2_18872_out0 = v$_12182_out1;
assign v$B23_1442_out0 = v$_9754_out1;
assign v$B23_1445_out0 = v$_9757_out1;
assign v$P$AB_2252_out0 = v$P$AD_864_out0;
assign v$P$AB_2256_out0 = v$P$AD_864_out0;
assign v$P$AB_2275_out0 = v$P$AD_864_out0;
assign v$P$AB_2283_out0 = v$P$AD_851_out0;
assign v$P$AB_2285_out0 = v$P$AD_864_out0;
assign v$P$AB_2375_out0 = v$P$AD_987_out0;
assign v$P$AB_2379_out0 = v$P$AD_987_out0;
assign v$P$AB_2398_out0 = v$P$AD_987_out0;
assign v$P$AB_2406_out0 = v$P$AD_974_out0;
assign v$P$AB_2408_out0 = v$P$AD_987_out0;
assign v$B_2920_out0 = v$B6_13884_out0;
assign v$B_2921_out0 = v$B3_9846_out0;
assign v$B_2922_out0 = v$B21_18690_out0;
assign v$B_2923_out0 = v$B9_4221_out0;
assign v$B_2924_out0 = v$B15_10447_out0;
assign v$B_2928_out0 = v$B12_2115_out0;
assign v$B_2932_out0 = v$B0_3422_out0;
assign v$B_2937_out0 = v$B18_11369_out0;
assign v$B_2992_out0 = v$B6_13887_out0;
assign v$B_2993_out0 = v$B3_9849_out0;
assign v$B_2994_out0 = v$B21_18693_out0;
assign v$B_2995_out0 = v$B9_4224_out0;
assign v$B_2996_out0 = v$B15_10450_out0;
assign v$B_3000_out0 = v$B12_2118_out0;
assign v$B_3004_out0 = v$B0_3425_out0;
assign v$B_3009_out0 = v$B18_11372_out0;
assign v$B2_3327_out0 = v$_11532_out1;
assign v$B2_3330_out0 = v$_11535_out1;
assign v$B20_4113_out0 = v$_17209_out1;
assign v$B20_4116_out0 = v$_17212_out1;
assign v$B14_4159_out0 = v$_17966_out1;
assign v$B14_4162_out0 = v$_17969_out1;
assign v$G5_4771_out0 = v$G$AB_9546_out0 && v$P$CD_10988_out0;
assign v$G5_4776_out0 = v$G$AB_9551_out0 && v$P$CD_10993_out0;
assign v$G5_4782_out0 = v$G$AB_9557_out0 && v$P$CD_10999_out0;
assign v$G5_4785_out0 = v$G$AB_9560_out0 && v$P$CD_11002_out0;
assign v$G5_4790_out0 = v$G$AB_9565_out0 && v$P$CD_11007_out0;
assign v$G5_4803_out0 = v$G$AB_9578_out0 && v$P$CD_11020_out0;
assign v$G5_4894_out0 = v$G$AB_9669_out0 && v$P$CD_11111_out0;
assign v$G5_4899_out0 = v$G$AB_9674_out0 && v$P$CD_11116_out0;
assign v$G5_4905_out0 = v$G$AB_9680_out0 && v$P$CD_11122_out0;
assign v$G5_4908_out0 = v$G$AB_9683_out0 && v$P$CD_11125_out0;
assign v$G5_4913_out0 = v$G$AB_9688_out0 && v$P$CD_11130_out0;
assign v$G5_4926_out0 = v$G$AB_9701_out0 && v$P$CD_11143_out0;
assign v$COUTD_7013_out0 = v$G6_535_out0;
assign v$COUTD_7014_out0 = v$G6_536_out0;
assign v$COUTD_7027_out0 = v$G6_549_out0;
assign v$COUTD_7029_out0 = v$G6_551_out0;
assign v$COUTD_7030_out0 = v$G6_552_out0;
assign v$COUTD_7033_out0 = v$G6_555_out0;
assign v$COUTD_7047_out0 = v$G6_569_out0;
assign v$COUTD_7052_out0 = v$G6_574_out0;
assign v$COUTD_7136_out0 = v$G6_658_out0;
assign v$COUTD_7137_out0 = v$G6_659_out0;
assign v$COUTD_7150_out0 = v$G6_672_out0;
assign v$COUTD_7152_out0 = v$G6_674_out0;
assign v$COUTD_7153_out0 = v$G6_675_out0;
assign v$COUTD_7156_out0 = v$G6_678_out0;
assign v$COUTD_7170_out0 = v$G6_692_out0;
assign v$COUTD_7175_out0 = v$G6_697_out0;
assign v$A_7420_out0 = v$A7_15892_out0;
assign v$A_7421_out0 = v$A1_1870_out0;
assign v$A_7422_out0 = v$A14_739_out0;
assign v$A_7424_out0 = v$A8_18698_out0;
assign v$A_7425_out0 = v$A17_17343_out0;
assign v$A_7426_out0 = v$A23_5282_out0;
assign v$A_7428_out0 = v$A13_14446_out0;
assign v$A_7429_out0 = v$A4_18139_out0;
assign v$A_7430_out0 = v$A19_1364_out0;
assign v$A_7431_out0 = v$A22_4591_out0;
assign v$A_7433_out0 = v$A10_1704_out0;
assign v$A_7434_out0 = v$A20_4604_out0;
assign v$A_7435_out0 = v$A2_18869_out0;
assign v$A_7436_out0 = v$A11_10387_out0;
assign v$A_7437_out0 = v$A5_6902_out0;
assign v$A_7438_out0 = v$A16_14192_out0;
assign v$A_7492_out0 = v$A7_15895_out0;
assign v$A_7493_out0 = v$A1_1873_out0;
assign v$A_7494_out0 = v$A14_742_out0;
assign v$A_7496_out0 = v$A8_18701_out0;
assign v$A_7497_out0 = v$A17_17346_out0;
assign v$A_7498_out0 = v$A23_5285_out0;
assign v$A_7500_out0 = v$A13_14449_out0;
assign v$A_7501_out0 = v$A4_18142_out0;
assign v$A_7502_out0 = v$A19_1367_out0;
assign v$A_7503_out0 = v$A22_4594_out0;
assign v$A_7505_out0 = v$A10_1707_out0;
assign v$A_7506_out0 = v$A20_4607_out0;
assign v$A_7507_out0 = v$A2_18872_out0;
assign v$A_7508_out0 = v$A11_10390_out0;
assign v$A_7509_out0 = v$A5_6905_out0;
assign v$A_7510_out0 = v$A16_14195_out0;
assign v$B1_8427_out0 = v$_11532_out0;
assign v$B1_8430_out0 = v$_11535_out0;
assign v$B13_9023_out0 = v$_17966_out0;
assign v$B13_9026_out0 = v$_17969_out0;
assign v$B11_9444_out0 = v$_9874_out1;
assign v$B11_9447_out0 = v$_9877_out1;
assign v$B10_10298_out0 = v$_9874_out0;
assign v$B10_10301_out0 = v$_9877_out0;
assign v$P$CD_10991_out0 = v$P$AD_851_out0;
assign v$P$CD_11017_out0 = v$P$AD_832_out0;
assign v$P$CD_11025_out0 = v$P$AD_846_out0;
assign v$P$CD_11114_out0 = v$P$AD_974_out0;
assign v$P$CD_11140_out0 = v$P$AD_955_out0;
assign v$P$CD_11148_out0 = v$P$AD_969_out0;
assign v$B22_11301_out0 = v$_9754_out0;
assign v$B22_11304_out0 = v$_9757_out0;
assign {v$A1A_12225_out1,v$A1A_12225_out0 } = v$A0_4469_out0 + v$B0_3422_out0 + v$C1_4634_out0;
assign {v$A1A_12228_out1,v$A1A_12228_out0 } = v$A0_4472_out0 + v$B0_3425_out0 + v$C1_4637_out0;
assign v$END11_12657_out0 = v$P$AD_843_out0;
assign v$END11_12660_out0 = v$P$AD_966_out0;
assign v$B8_13716_out0 = v$_7177_out1;
assign v$B8_13719_out0 = v$_7180_out1;
assign v$B4_15267_out0 = v$_7259_out0;
assign v$B4_15270_out0 = v$_7262_out0;
assign v$B17_16126_out0 = v$_13759_out1;
assign v$B17_16129_out0 = v$_13762_out1;
assign v$B16_17035_out0 = v$_13759_out0;
assign v$B16_17038_out0 = v$_13762_out0;
assign v$B19_17411_out0 = v$_17209_out0;
assign v$B19_17414_out0 = v$_17212_out0;
assign v$B7_17635_out0 = v$_7177_out0;
assign v$B7_17638_out0 = v$_7180_out0;
assign v$END13_18675_out0 = v$P$AD_837_out0;
assign v$END13_18678_out0 = v$P$AD_960_out0;
assign v$B5_18979_out0 = v$_7259_out1;
assign v$B5_18982_out0 = v$_7262_out1;
assign v$END1_1452_out0 = v$COUTD_7052_out0;
assign v$END1_1455_out0 = v$COUTD_7175_out0;
assign v$C2_2886_out0 = v$COUTD_7029_out0;
assign v$C2_2889_out0 = v$COUTD_7152_out0;
assign v$B_2925_out0 = v$B7_17635_out0;
assign v$B_2926_out0 = v$B1_8427_out0;
assign v$B_2927_out0 = v$B14_4159_out0;
assign v$B_2929_out0 = v$B8_13716_out0;
assign v$B_2930_out0 = v$B17_16126_out0;
assign v$B_2931_out0 = v$B23_1442_out0;
assign v$B_2933_out0 = v$B13_9023_out0;
assign v$B_2934_out0 = v$B4_15267_out0;
assign v$B_2935_out0 = v$B19_17411_out0;
assign v$B_2936_out0 = v$B22_11301_out0;
assign v$B_2938_out0 = v$B10_10298_out0;
assign v$B_2939_out0 = v$B20_4113_out0;
assign v$B_2940_out0 = v$B2_3327_out0;
assign v$B_2941_out0 = v$B11_9444_out0;
assign v$B_2942_out0 = v$B5_18979_out0;
assign v$B_2943_out0 = v$B16_17035_out0;
assign v$B_2997_out0 = v$B7_17638_out0;
assign v$B_2998_out0 = v$B1_8430_out0;
assign v$B_2999_out0 = v$B14_4162_out0;
assign v$B_3001_out0 = v$B8_13719_out0;
assign v$B_3002_out0 = v$B17_16129_out0;
assign v$B_3003_out0 = v$B23_1445_out0;
assign v$B_3005_out0 = v$B13_9026_out0;
assign v$B_3006_out0 = v$B4_15270_out0;
assign v$B_3007_out0 = v$B19_17414_out0;
assign v$B_3008_out0 = v$B22_11304_out0;
assign v$B_3010_out0 = v$B10_10301_out0;
assign v$B_3011_out0 = v$B20_4116_out0;
assign v$B_3012_out0 = v$B2_3330_out0;
assign v$B_3013_out0 = v$B11_9447_out0;
assign v$B_3014_out0 = v$B5_18982_out0;
assign v$B_3015_out0 = v$B16_17038_out0;
assign v$END_3543_out0 = v$COUTD_7030_out0;
assign v$END_3546_out0 = v$COUTD_7153_out0;
assign v$END3_3657_out0 = v$COUTD_7027_out0;
assign v$END3_3660_out0 = v$COUTD_7150_out0;
assign v$G2_5502_out0 = ((v$A_7415_out0 && !v$B_2920_out0) || (!v$A_7415_out0) && v$B_2920_out0);
assign v$G2_5503_out0 = ((v$A_7416_out0 && !v$B_2921_out0) || (!v$A_7416_out0) && v$B_2921_out0);
assign v$G2_5504_out0 = ((v$A_7417_out0 && !v$B_2922_out0) || (!v$A_7417_out0) && v$B_2922_out0);
assign v$G2_5505_out0 = ((v$A_7418_out0 && !v$B_2923_out0) || (!v$A_7418_out0) && v$B_2923_out0);
assign v$G2_5506_out0 = ((v$A_7419_out0 && !v$B_2924_out0) || (!v$A_7419_out0) && v$B_2924_out0);
assign v$G2_5510_out0 = ((v$A_7423_out0 && !v$B_2928_out0) || (!v$A_7423_out0) && v$B_2928_out0);
assign v$G2_5514_out0 = ((v$A_7427_out0 && !v$B_2932_out0) || (!v$A_7427_out0) && v$B_2932_out0);
assign v$G2_5519_out0 = ((v$A_7432_out0 && !v$B_2937_out0) || (!v$A_7432_out0) && v$B_2937_out0);
assign v$G2_5574_out0 = ((v$A_7487_out0 && !v$B_2992_out0) || (!v$A_7487_out0) && v$B_2992_out0);
assign v$G2_5575_out0 = ((v$A_7488_out0 && !v$B_2993_out0) || (!v$A_7488_out0) && v$B_2993_out0);
assign v$G2_5576_out0 = ((v$A_7489_out0 && !v$B_2994_out0) || (!v$A_7489_out0) && v$B_2994_out0);
assign v$G2_5577_out0 = ((v$A_7490_out0 && !v$B_2995_out0) || (!v$A_7490_out0) && v$B_2995_out0);
assign v$G2_5578_out0 = ((v$A_7491_out0 && !v$B_2996_out0) || (!v$A_7491_out0) && v$B_2996_out0);
assign v$G2_5582_out0 = ((v$A_7495_out0 && !v$B_3000_out0) || (!v$A_7495_out0) && v$B_3000_out0);
assign v$G2_5586_out0 = ((v$A_7499_out0 && !v$B_3004_out0) || (!v$A_7499_out0) && v$B_3004_out0);
assign v$G2_5591_out0 = ((v$A_7504_out0 && !v$B_3009_out0) || (!v$A_7504_out0) && v$B_3009_out0);
assign v$G1_5851_out0 = v$P$AB_2252_out0 && v$P$CD_10994_out0;
assign v$G1_5855_out0 = v$P$AB_2256_out0 && v$P$CD_10998_out0;
assign v$G1_5874_out0 = v$P$AB_2275_out0 && v$P$CD_11017_out0;
assign v$G1_5882_out0 = v$P$AB_2283_out0 && v$P$CD_11025_out0;
assign v$G1_5884_out0 = v$P$AB_2285_out0 && v$P$CD_11027_out0;
assign v$G1_5974_out0 = v$P$AB_2375_out0 && v$P$CD_11117_out0;
assign v$G1_5978_out0 = v$P$AB_2379_out0 && v$P$CD_11121_out0;
assign v$G1_5997_out0 = v$P$AB_2398_out0 && v$P$CD_11140_out0;
assign v$G1_6005_out0 = v$P$AB_2406_out0 && v$P$CD_11148_out0;
assign v$G1_6007_out0 = v$P$AB_2408_out0 && v$P$CD_11150_out0;
assign v$END2_8070_out0 = v$COUTD_7033_out0;
assign v$END2_8073_out0 = v$COUTD_7156_out0;
assign v$CINA_8852_out0 = v$COUTD_7014_out0;
assign v$CINA_8857_out0 = v$COUTD_7029_out0;
assign v$CINA_8863_out0 = v$COUTD_7029_out0;
assign v$CINA_8866_out0 = v$COUTD_7047_out0;
assign v$CINA_8871_out0 = v$COUTD_7013_out0;
assign v$CINA_8884_out0 = v$COUTD_7029_out0;
assign v$CINA_8975_out0 = v$COUTD_7137_out0;
assign v$CINA_8980_out0 = v$COUTD_7152_out0;
assign v$CINA_8986_out0 = v$COUTD_7152_out0;
assign v$CINA_8989_out0 = v$COUTD_7170_out0;
assign v$CINA_8994_out0 = v$COUTD_7136_out0;
assign v$CINA_9007_out0 = v$COUTD_7152_out0;
assign v$END45_9385_out0 = v$COUTD_7047_out0;
assign v$END45_9388_out0 = v$COUTD_7170_out0;
assign v$G4_11692_out0 = v$G5_4771_out0 || v$G$CD_1099_out0;
assign v$G4_11697_out0 = v$G5_4776_out0 || v$G$CD_1104_out0;
assign v$G4_11703_out0 = v$G5_4782_out0 || v$G$CD_1110_out0;
assign v$G4_11706_out0 = v$G5_4785_out0 || v$G$CD_1113_out0;
assign v$G4_11711_out0 = v$G5_4790_out0 || v$G$CD_1118_out0;
assign v$G4_11724_out0 = v$G5_4803_out0 || v$G$CD_1131_out0;
assign v$G4_11815_out0 = v$G5_4894_out0 || v$G$CD_1222_out0;
assign v$G4_11820_out0 = v$G5_4899_out0 || v$G$CD_1227_out0;
assign v$G4_11826_out0 = v$G5_4905_out0 || v$G$CD_1233_out0;
assign v$G4_11829_out0 = v$G5_4908_out0 || v$G$CD_1236_out0;
assign v$G4_11834_out0 = v$G5_4913_out0 || v$G$CD_1241_out0;
assign v$G4_11847_out0 = v$G5_4926_out0 || v$G$CD_1254_out0;
assign v$G1_12926_out0 = v$A_7415_out0 && v$B_2920_out0;
assign v$G1_12927_out0 = v$A_7416_out0 && v$B_2921_out0;
assign v$G1_12928_out0 = v$A_7417_out0 && v$B_2922_out0;
assign v$G1_12929_out0 = v$A_7418_out0 && v$B_2923_out0;
assign v$G1_12930_out0 = v$A_7419_out0 && v$B_2924_out0;
assign v$G1_12934_out0 = v$A_7423_out0 && v$B_2928_out0;
assign v$G1_12938_out0 = v$A_7427_out0 && v$B_2932_out0;
assign v$G1_12943_out0 = v$A_7432_out0 && v$B_2937_out0;
assign v$G1_12998_out0 = v$A_7487_out0 && v$B_2992_out0;
assign v$G1_12999_out0 = v$A_7488_out0 && v$B_2993_out0;
assign v$G1_13000_out0 = v$A_7489_out0 && v$B_2994_out0;
assign v$G1_13001_out0 = v$A_7490_out0 && v$B_2995_out0;
assign v$G1_13002_out0 = v$A_7491_out0 && v$B_2996_out0;
assign v$G1_13006_out0 = v$A_7495_out0 && v$B_3000_out0;
assign v$G1_13010_out0 = v$A_7499_out0 && v$B_3004_out0;
assign v$G1_13015_out0 = v$A_7504_out0 && v$B_3009_out0;
assign v$END_18876_out0 = v$A1A_12225_out1;
assign v$END_18879_out0 = v$A1A_12228_out1;
assign v$P$AD_838_out0 = v$G1_5851_out0;
assign v$P$AD_842_out0 = v$G1_5855_out0;
assign v$P$AD_861_out0 = v$G1_5874_out0;
assign v$P$AD_869_out0 = v$G1_5882_out0;
assign v$P$AD_871_out0 = v$G1_5884_out0;
assign v$P$AD_961_out0 = v$G1_5974_out0;
assign v$P$AD_965_out0 = v$G1_5978_out0;
assign v$P$AD_984_out0 = v$G1_5997_out0;
assign v$P$AD_992_out0 = v$G1_6005_out0;
assign v$P$AD_994_out0 = v$G1_6007_out0;
assign v$G2_5507_out0 = ((v$A_7420_out0 && !v$B_2925_out0) || (!v$A_7420_out0) && v$B_2925_out0);
assign v$G2_5508_out0 = ((v$A_7421_out0 && !v$B_2926_out0) || (!v$A_7421_out0) && v$B_2926_out0);
assign v$G2_5509_out0 = ((v$A_7422_out0 && !v$B_2927_out0) || (!v$A_7422_out0) && v$B_2927_out0);
assign v$G2_5511_out0 = ((v$A_7424_out0 && !v$B_2929_out0) || (!v$A_7424_out0) && v$B_2929_out0);
assign v$G2_5512_out0 = ((v$A_7425_out0 && !v$B_2930_out0) || (!v$A_7425_out0) && v$B_2930_out0);
assign v$G2_5513_out0 = ((v$A_7426_out0 && !v$B_2931_out0) || (!v$A_7426_out0) && v$B_2931_out0);
assign v$G2_5515_out0 = ((v$A_7428_out0 && !v$B_2933_out0) || (!v$A_7428_out0) && v$B_2933_out0);
assign v$G2_5516_out0 = ((v$A_7429_out0 && !v$B_2934_out0) || (!v$A_7429_out0) && v$B_2934_out0);
assign v$G2_5517_out0 = ((v$A_7430_out0 && !v$B_2935_out0) || (!v$A_7430_out0) && v$B_2935_out0);
assign v$G2_5518_out0 = ((v$A_7431_out0 && !v$B_2936_out0) || (!v$A_7431_out0) && v$B_2936_out0);
assign v$G2_5520_out0 = ((v$A_7433_out0 && !v$B_2938_out0) || (!v$A_7433_out0) && v$B_2938_out0);
assign v$G2_5521_out0 = ((v$A_7434_out0 && !v$B_2939_out0) || (!v$A_7434_out0) && v$B_2939_out0);
assign v$G2_5522_out0 = ((v$A_7435_out0 && !v$B_2940_out0) || (!v$A_7435_out0) && v$B_2940_out0);
assign v$G2_5523_out0 = ((v$A_7436_out0 && !v$B_2941_out0) || (!v$A_7436_out0) && v$B_2941_out0);
assign v$G2_5524_out0 = ((v$A_7437_out0 && !v$B_2942_out0) || (!v$A_7437_out0) && v$B_2942_out0);
assign v$G2_5525_out0 = ((v$A_7438_out0 && !v$B_2943_out0) || (!v$A_7438_out0) && v$B_2943_out0);
assign v$G2_5579_out0 = ((v$A_7492_out0 && !v$B_2997_out0) || (!v$A_7492_out0) && v$B_2997_out0);
assign v$G2_5580_out0 = ((v$A_7493_out0 && !v$B_2998_out0) || (!v$A_7493_out0) && v$B_2998_out0);
assign v$G2_5581_out0 = ((v$A_7494_out0 && !v$B_2999_out0) || (!v$A_7494_out0) && v$B_2999_out0);
assign v$G2_5583_out0 = ((v$A_7496_out0 && !v$B_3001_out0) || (!v$A_7496_out0) && v$B_3001_out0);
assign v$G2_5584_out0 = ((v$A_7497_out0 && !v$B_3002_out0) || (!v$A_7497_out0) && v$B_3002_out0);
assign v$G2_5585_out0 = ((v$A_7498_out0 && !v$B_3003_out0) || (!v$A_7498_out0) && v$B_3003_out0);
assign v$G2_5587_out0 = ((v$A_7500_out0 && !v$B_3005_out0) || (!v$A_7500_out0) && v$B_3005_out0);
assign v$G2_5588_out0 = ((v$A_7501_out0 && !v$B_3006_out0) || (!v$A_7501_out0) && v$B_3006_out0);
assign v$G2_5589_out0 = ((v$A_7502_out0 && !v$B_3007_out0) || (!v$A_7502_out0) && v$B_3007_out0);
assign v$G2_5590_out0 = ((v$A_7503_out0 && !v$B_3008_out0) || (!v$A_7503_out0) && v$B_3008_out0);
assign v$G2_5592_out0 = ((v$A_7505_out0 && !v$B_3010_out0) || (!v$A_7505_out0) && v$B_3010_out0);
assign v$G2_5593_out0 = ((v$A_7506_out0 && !v$B_3011_out0) || (!v$A_7506_out0) && v$B_3011_out0);
assign v$G2_5594_out0 = ((v$A_7507_out0 && !v$B_3012_out0) || (!v$A_7507_out0) && v$B_3012_out0);
assign v$G2_5595_out0 = ((v$A_7508_out0 && !v$B_3013_out0) || (!v$A_7508_out0) && v$B_3013_out0);
assign v$G2_5596_out0 = ((v$A_7509_out0 && !v$B_3014_out0) || (!v$A_7509_out0) && v$B_3014_out0);
assign v$G2_5597_out0 = ((v$A_7510_out0 && !v$B_3015_out0) || (!v$A_7510_out0) && v$B_3015_out0);
assign v$G_10506_out0 = v$G1_12926_out0;
assign v$G_10507_out0 = v$G1_12927_out0;
assign v$G_10508_out0 = v$G1_12928_out0;
assign v$G_10509_out0 = v$G1_12929_out0;
assign v$G_10510_out0 = v$G1_12930_out0;
assign v$G_10514_out0 = v$G1_12934_out0;
assign v$G_10518_out0 = v$G1_12938_out0;
assign v$G_10523_out0 = v$G1_12943_out0;
assign v$G_10578_out0 = v$G1_12998_out0;
assign v$G_10579_out0 = v$G1_12999_out0;
assign v$G_10580_out0 = v$G1_13000_out0;
assign v$G_10581_out0 = v$G1_13001_out0;
assign v$G_10582_out0 = v$G1_13002_out0;
assign v$G_10586_out0 = v$G1_13006_out0;
assign v$G_10590_out0 = v$G1_13010_out0;
assign v$G_10595_out0 = v$G1_13015_out0;
assign v$G8_12007_out0 = v$CINA_8852_out0 && v$P$AB_2246_out0;
assign v$G8_12012_out0 = v$CINA_8857_out0 && v$P$AB_2251_out0;
assign v$G8_12018_out0 = v$CINA_8863_out0 && v$P$AB_2257_out0;
assign v$G8_12021_out0 = v$CINA_8866_out0 && v$P$AB_2260_out0;
assign v$G8_12026_out0 = v$CINA_8871_out0 && v$P$AB_2265_out0;
assign v$G8_12039_out0 = v$CINA_8884_out0 && v$P$AB_2278_out0;
assign v$G8_12130_out0 = v$CINA_8975_out0 && v$P$AB_2369_out0;
assign v$G8_12135_out0 = v$CINA_8980_out0 && v$P$AB_2374_out0;
assign v$G8_12141_out0 = v$CINA_8986_out0 && v$P$AB_2380_out0;
assign v$G8_12144_out0 = v$CINA_8989_out0 && v$P$AB_2383_out0;
assign v$G8_12149_out0 = v$CINA_8994_out0 && v$P$AB_2388_out0;
assign v$G8_12162_out0 = v$CINA_9007_out0 && v$P$AB_2401_out0;
assign v$G1_12931_out0 = v$A_7420_out0 && v$B_2925_out0;
assign v$G1_12932_out0 = v$A_7421_out0 && v$B_2926_out0;
assign v$G1_12933_out0 = v$A_7422_out0 && v$B_2927_out0;
assign v$G1_12935_out0 = v$A_7424_out0 && v$B_2929_out0;
assign v$G1_12936_out0 = v$A_7425_out0 && v$B_2930_out0;
assign v$G1_12937_out0 = v$A_7426_out0 && v$B_2931_out0;
assign v$G1_12939_out0 = v$A_7428_out0 && v$B_2933_out0;
assign v$G1_12940_out0 = v$A_7429_out0 && v$B_2934_out0;
assign v$G1_12941_out0 = v$A_7430_out0 && v$B_2935_out0;
assign v$G1_12942_out0 = v$A_7431_out0 && v$B_2936_out0;
assign v$G1_12944_out0 = v$A_7433_out0 && v$B_2938_out0;
assign v$G1_12945_out0 = v$A_7434_out0 && v$B_2939_out0;
assign v$G1_12946_out0 = v$A_7435_out0 && v$B_2940_out0;
assign v$G1_12947_out0 = v$A_7436_out0 && v$B_2941_out0;
assign v$G1_12948_out0 = v$A_7437_out0 && v$B_2942_out0;
assign v$G1_12949_out0 = v$A_7438_out0 && v$B_2943_out0;
assign v$G1_13003_out0 = v$A_7492_out0 && v$B_2997_out0;
assign v$G1_13004_out0 = v$A_7493_out0 && v$B_2998_out0;
assign v$G1_13005_out0 = v$A_7494_out0 && v$B_2999_out0;
assign v$G1_13007_out0 = v$A_7496_out0 && v$B_3001_out0;
assign v$G1_13008_out0 = v$A_7497_out0 && v$B_3002_out0;
assign v$G1_13009_out0 = v$A_7498_out0 && v$B_3003_out0;
assign v$G1_13011_out0 = v$A_7500_out0 && v$B_3005_out0;
assign v$G1_13012_out0 = v$A_7501_out0 && v$B_3006_out0;
assign v$G1_13013_out0 = v$A_7502_out0 && v$B_3007_out0;
assign v$G1_13014_out0 = v$A_7503_out0 && v$B_3008_out0;
assign v$G1_13016_out0 = v$A_7505_out0 && v$B_3010_out0;
assign v$G1_13017_out0 = v$A_7506_out0 && v$B_3011_out0;
assign v$G1_13018_out0 = v$A_7507_out0 && v$B_3012_out0;
assign v$G1_13019_out0 = v$A_7508_out0 && v$B_3013_out0;
assign v$G1_13020_out0 = v$A_7509_out0 && v$B_3014_out0;
assign v$G1_13021_out0 = v$A_7510_out0 && v$B_3015_out0;
assign {v$A4A_13733_out1,v$A4A_13733_out0 } = v$A3_15211_out0 + v$B3_9847_out0 + v$C2_2886_out0;
assign {v$A4A_13736_out1,v$A4A_13736_out0 } = v$A3_15214_out0 + v$B3_9850_out0 + v$C2_2889_out0;
assign v$P_14477_out0 = v$G2_5502_out0;
assign v$P_14478_out0 = v$G2_5503_out0;
assign v$P_14479_out0 = v$G2_5504_out0;
assign v$P_14480_out0 = v$G2_5505_out0;
assign v$P_14481_out0 = v$G2_5506_out0;
assign v$P_14485_out0 = v$G2_5510_out0;
assign v$P_14489_out0 = v$G2_5514_out0;
assign v$P_14494_out0 = v$G2_5519_out0;
assign v$P_14549_out0 = v$G2_5574_out0;
assign v$P_14550_out0 = v$G2_5575_out0;
assign v$P_14551_out0 = v$G2_5576_out0;
assign v$P_14552_out0 = v$G2_5577_out0;
assign v$P_14553_out0 = v$G2_5578_out0;
assign v$P_14557_out0 = v$G2_5582_out0;
assign v$P_14561_out0 = v$G2_5586_out0;
assign v$P_14566_out0 = v$G2_5591_out0;
assign v$G$AD_17766_out0 = v$G4_11692_out0;
assign v$G$AD_17771_out0 = v$G4_11697_out0;
assign v$G$AD_17777_out0 = v$G4_11703_out0;
assign v$G$AD_17780_out0 = v$G4_11706_out0;
assign v$G$AD_17785_out0 = v$G4_11711_out0;
assign v$G$AD_17798_out0 = v$G4_11724_out0;
assign v$G$AD_17889_out0 = v$G4_11815_out0;
assign v$G$AD_17894_out0 = v$G4_11820_out0;
assign v$G$AD_17900_out0 = v$G4_11826_out0;
assign v$G$AD_17903_out0 = v$G4_11829_out0;
assign v$G$AD_17908_out0 = v$G4_11834_out0;
assign v$G$AD_17921_out0 = v$G4_11847_out0;
assign v$C2_18779_out0 = v$C2_2886_out0;
assign v$C2_18782_out0 = v$C2_2889_out0;
assign v$P12_244_out0 = v$P_14485_out0;
assign v$P12_247_out0 = v$P_14557_out0;
assign v$G$CD_1102_out0 = v$G$AD_17785_out0;
assign v$G$CD_1128_out0 = v$G$AD_17766_out0;
assign v$G$CD_1136_out0 = v$G$AD_17780_out0;
assign v$G$CD_1225_out0 = v$G$AD_17908_out0;
assign v$G$CD_1251_out0 = v$G$AD_17889_out0;
assign v$G$CD_1259_out0 = v$G$AD_17903_out0;
assign v$END10_1297_out0 = v$G$AD_17777_out0;
assign v$END10_1300_out0 = v$G$AD_17900_out0;
assign v$P$AB_2249_out0 = v$P$AD_861_out0;
assign v$P$AB_2258_out0 = v$P$AD_861_out0;
assign v$P$AB_2259_out0 = v$P$AD_838_out0;
assign v$P$AB_2270_out0 = v$P$AD_861_out0;
assign v$P$AB_2272_out0 = v$P$AD_861_out0;
assign v$P$AB_2279_out0 = v$P$AD_861_out0;
assign v$P$AB_2280_out0 = v$P$AD_838_out0;
assign v$P$AB_2372_out0 = v$P$AD_984_out0;
assign v$P$AB_2381_out0 = v$P$AD_984_out0;
assign v$P$AB_2382_out0 = v$P$AD_961_out0;
assign v$P$AB_2393_out0 = v$P$AD_984_out0;
assign v$P$AB_2395_out0 = v$P$AD_984_out0;
assign v$P$AB_2402_out0 = v$P$AD_984_out0;
assign v$P$AB_2403_out0 = v$P$AD_961_out0;
assign v$P21_4982_out0 = v$P_14479_out0;
assign v$P21_4985_out0 = v$P_14551_out0;
assign v$P0_5024_out0 = v$P_14489_out0;
assign v$P0_5027_out0 = v$P_14561_out0;
assign v$P15_7184_out0 = v$P_14481_out0;
assign v$P15_7187_out0 = v$P_14553_out0;
assign v$G12_7328_out0 = v$G_10514_out0;
assign v$G12_7331_out0 = v$G_10586_out0;
assign v$END15_7698_out0 = v$P$AD_842_out0;
assign v$END15_7701_out0 = v$P$AD_965_out0;
assign v$END17_7967_out0 = v$P$AD_871_out0;
assign v$END17_7970_out0 = v$P$AD_994_out0;
assign v$END3_8259_out0 = v$A4A_13733_out1;
assign v$END3_8262_out0 = v$A4A_13736_out1;
assign v$P6_8419_out0 = v$P_14477_out0;
assign v$P6_8422_out0 = v$P_14549_out0;
assign v$G9_9256_out0 = v$G_10509_out0;
assign v$G9_9259_out0 = v$G_10581_out0;
assign v$G$AB_9552_out0 = v$G$AD_17798_out0;
assign v$G$AB_9556_out0 = v$G$AD_17798_out0;
assign v$G$AB_9575_out0 = v$G$AD_17798_out0;
assign v$G$AB_9583_out0 = v$G$AD_17785_out0;
assign v$G$AB_9585_out0 = v$G$AD_17798_out0;
assign v$G$AB_9675_out0 = v$G$AD_17921_out0;
assign v$G$AB_9679_out0 = v$G$AD_17921_out0;
assign v$G$AB_9698_out0 = v$G$AD_17921_out0;
assign v$G$AB_9706_out0 = v$G$AD_17908_out0;
assign v$G$AB_9708_out0 = v$G$AD_17921_out0;
assign v$G7_10099_out0 = v$G8_12007_out0 && v$P$CD_10988_out0;
assign v$G7_10104_out0 = v$G8_12012_out0 && v$P$CD_10993_out0;
assign v$G7_10110_out0 = v$G8_12018_out0 && v$P$CD_10999_out0;
assign v$G7_10113_out0 = v$G8_12021_out0 && v$P$CD_11002_out0;
assign v$G7_10118_out0 = v$G8_12026_out0 && v$P$CD_11007_out0;
assign v$G7_10131_out0 = v$G8_12039_out0 && v$P$CD_11020_out0;
assign v$G7_10222_out0 = v$G8_12130_out0 && v$P$CD_11111_out0;
assign v$G7_10227_out0 = v$G8_12135_out0 && v$P$CD_11116_out0;
assign v$G7_10233_out0 = v$G8_12141_out0 && v$P$CD_11122_out0;
assign v$G7_10236_out0 = v$G8_12144_out0 && v$P$CD_11125_out0;
assign v$G7_10241_out0 = v$G8_12149_out0 && v$P$CD_11130_out0;
assign v$G7_10254_out0 = v$G8_12162_out0 && v$P$CD_11143_out0;
assign v$G_10511_out0 = v$G1_12931_out0;
assign v$G_10512_out0 = v$G1_12932_out0;
assign v$G_10513_out0 = v$G1_12933_out0;
assign v$G_10515_out0 = v$G1_12935_out0;
assign v$G_10516_out0 = v$G1_12936_out0;
assign v$G_10517_out0 = v$G1_12937_out0;
assign v$G_10519_out0 = v$G1_12939_out0;
assign v$G_10520_out0 = v$G1_12940_out0;
assign v$G_10521_out0 = v$G1_12941_out0;
assign v$G_10522_out0 = v$G1_12942_out0;
assign v$G_10524_out0 = v$G1_12944_out0;
assign v$G_10525_out0 = v$G1_12945_out0;
assign v$G_10526_out0 = v$G1_12946_out0;
assign v$G_10527_out0 = v$G1_12947_out0;
assign v$G_10528_out0 = v$G1_12948_out0;
assign v$G_10529_out0 = v$G1_12949_out0;
assign v$G_10583_out0 = v$G1_13003_out0;
assign v$G_10584_out0 = v$G1_13004_out0;
assign v$G_10585_out0 = v$G1_13005_out0;
assign v$G_10587_out0 = v$G1_13007_out0;
assign v$G_10588_out0 = v$G1_13008_out0;
assign v$G_10589_out0 = v$G1_13009_out0;
assign v$G_10591_out0 = v$G1_13011_out0;
assign v$G_10592_out0 = v$G1_13012_out0;
assign v$G_10593_out0 = v$G1_13013_out0;
assign v$G_10594_out0 = v$G1_13014_out0;
assign v$G_10596_out0 = v$G1_13016_out0;
assign v$G_10597_out0 = v$G1_13017_out0;
assign v$G_10598_out0 = v$G1_13018_out0;
assign v$G_10599_out0 = v$G1_13019_out0;
assign v$G_10600_out0 = v$G1_13020_out0;
assign v$G_10601_out0 = v$G1_13021_out0;
assign v$P$CD_11014_out0 = v$P$AD_869_out0;
assign v$P$CD_11137_out0 = v$P$AD_992_out0;
assign v$END12_11276_out0 = v$G$AD_17771_out0;
assign v$END12_11279_out0 = v$G$AD_17894_out0;
assign v$G15_11542_out0 = v$G_10510_out0;
assign v$G15_11545_out0 = v$G_10582_out0;
assign v$G3_11603_out0 = v$G_10507_out0;
assign v$G3_11606_out0 = v$G_10579_out0;
assign v$END19_12220_out0 = v$P$AD_838_out0;
assign v$END19_12223_out0 = v$P$AD_961_out0;
assign v$P18_12291_out0 = v$P_14494_out0;
assign v$P18_12294_out0 = v$P_14566_out0;
assign v$G18_13509_out0 = v$G_10523_out0;
assign v$G18_13512_out0 = v$G_10595_out0;
assign v$P_14482_out0 = v$G2_5507_out0;
assign v$P_14483_out0 = v$G2_5508_out0;
assign v$P_14484_out0 = v$G2_5509_out0;
assign v$P_14486_out0 = v$G2_5511_out0;
assign v$P_14487_out0 = v$G2_5512_out0;
assign v$P_14488_out0 = v$G2_5513_out0;
assign v$P_14490_out0 = v$G2_5515_out0;
assign v$P_14491_out0 = v$G2_5516_out0;
assign v$P_14492_out0 = v$G2_5517_out0;
assign v$P_14493_out0 = v$G2_5518_out0;
assign v$P_14495_out0 = v$G2_5520_out0;
assign v$P_14496_out0 = v$G2_5521_out0;
assign v$P_14497_out0 = v$G2_5522_out0;
assign v$P_14498_out0 = v$G2_5523_out0;
assign v$P_14499_out0 = v$G2_5524_out0;
assign v$P_14500_out0 = v$G2_5525_out0;
assign v$P_14554_out0 = v$G2_5579_out0;
assign v$P_14555_out0 = v$G2_5580_out0;
assign v$P_14556_out0 = v$G2_5581_out0;
assign v$P_14558_out0 = v$G2_5583_out0;
assign v$P_14559_out0 = v$G2_5584_out0;
assign v$P_14560_out0 = v$G2_5585_out0;
assign v$P_14562_out0 = v$G2_5587_out0;
assign v$P_14563_out0 = v$G2_5588_out0;
assign v$P_14564_out0 = v$G2_5589_out0;
assign v$P_14565_out0 = v$G2_5590_out0;
assign v$P_14567_out0 = v$G2_5592_out0;
assign v$P_14568_out0 = v$G2_5593_out0;
assign v$P_14569_out0 = v$G2_5594_out0;
assign v$P_14570_out0 = v$G2_5595_out0;
assign v$P_14571_out0 = v$G2_5596_out0;
assign v$P_14572_out0 = v$G2_5597_out0;
assign v$G21_14627_out0 = v$G_10508_out0;
assign v$G21_14630_out0 = v$G_10580_out0;
assign v$P3_15922_out0 = v$P_14478_out0;
assign v$P3_15925_out0 = v$P_14550_out0;
assign v$G0_16549_out0 = v$G_10518_out0;
assign v$G0_16552_out0 = v$G_10590_out0;
assign v$G6_16971_out0 = v$G_10506_out0;
assign v$G6_16974_out0 = v$G_10578_out0;
assign v$P9_19054_out0 = v$P_14480_out0;
assign v$P9_19057_out0 = v$P_14552_out0;
assign v$_19276_out0 = { v$A3A_12527_out0,v$A4A_13733_out0 };
assign v$_19279_out0 = { v$A3A_12530_out0,v$A4A_13736_out0 };
assign v$P5_229_out0 = v$P_14499_out0;
assign v$P5_232_out0 = v$P_14571_out0;
assign v$P10_361_out0 = v$P_14495_out0;
assign v$P10_364_out0 = v$P_14567_out0;
assign v$G6_534_out0 = v$G4_11692_out0 || v$G7_10099_out0;
assign v$G6_539_out0 = v$G4_11697_out0 || v$G7_10104_out0;
assign v$G6_545_out0 = v$G4_11703_out0 || v$G7_10110_out0;
assign v$G6_548_out0 = v$G4_11706_out0 || v$G7_10113_out0;
assign v$G6_553_out0 = v$G4_11711_out0 || v$G7_10118_out0;
assign v$G6_566_out0 = v$G4_11724_out0 || v$G7_10131_out0;
assign v$G6_657_out0 = v$G4_11815_out0 || v$G7_10222_out0;
assign v$G6_662_out0 = v$G4_11820_out0 || v$G7_10227_out0;
assign v$G6_668_out0 = v$G4_11826_out0 || v$G7_10233_out0;
assign v$G6_671_out0 = v$G4_11829_out0 || v$G7_10236_out0;
assign v$G6_676_out0 = v$G4_11834_out0 || v$G7_10241_out0;
assign v$G6_689_out0 = v$G4_11847_out0 || v$G7_10254_out0;
assign v$G$CD_1068_out0 = v$G6_16971_out0;
assign v$G$CD_1069_out0 = v$G3_11603_out0;
assign v$G$CD_1070_out0 = v$G12_7328_out0;
assign v$G$CD_1071_out0 = v$G9_9256_out0;
assign v$G$CD_1074_out0 = v$G18_13509_out0;
assign v$G$CD_1085_out0 = v$G15_11542_out0;
assign v$G$CD_1086_out0 = v$G21_14627_out0;
assign v$G$CD_1191_out0 = v$G6_16974_out0;
assign v$G$CD_1192_out0 = v$G3_11606_out0;
assign v$G$CD_1193_out0 = v$G12_7331_out0;
assign v$G$CD_1194_out0 = v$G9_9259_out0;
assign v$G$CD_1197_out0 = v$G18_13512_out0;
assign v$G$CD_1208_out0 = v$G15_11545_out0;
assign v$G$CD_1209_out0 = v$G21_14630_out0;
assign v$G7_1850_out0 = v$G_10511_out0;
assign v$G7_1853_out0 = v$G_10583_out0;
assign v$P8_1862_out0 = v$P_14486_out0;
assign v$P8_1865_out0 = v$P_14558_out0;
assign v$G10_1994_out0 = v$G_10524_out0;
assign v$G10_1997_out0 = v$G_10596_out0;
assign v$G19_2045_out0 = v$G_10521_out0;
assign v$G19_2048_out0 = v$G_10593_out0;
assign v$P$AB_2209_out0 = v$P0_5024_out0;
assign v$P$AB_2212_out0 = v$P18_12291_out0;
assign v$P$AB_2213_out0 = v$P21_4982_out0;
assign v$P$AB_2225_out0 = v$P12_244_out0;
assign v$P$AB_2227_out0 = v$P15_7184_out0;
assign v$P$AB_2230_out0 = v$P6_8419_out0;
assign v$P$AB_2236_out0 = v$P3_15922_out0;
assign v$P$AB_2241_out0 = v$P9_19054_out0;
assign v$P$AB_2332_out0 = v$P0_5027_out0;
assign v$P$AB_2335_out0 = v$P18_12294_out0;
assign v$P$AB_2336_out0 = v$P21_4985_out0;
assign v$P$AB_2348_out0 = v$P12_247_out0;
assign v$P$AB_2350_out0 = v$P15_7187_out0;
assign v$P$AB_2353_out0 = v$P6_8422_out0;
assign v$P$AB_2359_out0 = v$P3_15925_out0;
assign v$P$AB_2364_out0 = v$P9_19057_out0;
assign v$P2_2425_out0 = v$P_14497_out0;
assign v$P2_2428_out0 = v$P_14569_out0;
assign v$G8_2771_out0 = v$G_10515_out0;
assign v$G8_2774_out0 = v$G_10587_out0;
assign v$G13_3053_out0 = v$G_10519_out0;
assign v$G13_3056_out0 = v$G_10591_out0;
assign v$P1_3169_out0 = v$P_14483_out0;
assign v$P1_3172_out0 = v$P_14555_out0;
assign v$P13_3246_out0 = v$P_14490_out0;
assign v$P13_3249_out0 = v$P_14562_out0;
assign v$P14_3370_out0 = v$P_14484_out0;
assign v$P14_3373_out0 = v$P_14556_out0;
assign v$G5_4777_out0 = v$G$AB_9552_out0 && v$P$CD_10994_out0;
assign v$G5_4781_out0 = v$G$AB_9556_out0 && v$P$CD_10998_out0;
assign v$G5_4800_out0 = v$G$AB_9575_out0 && v$P$CD_11017_out0;
assign v$G5_4808_out0 = v$G$AB_9583_out0 && v$P$CD_11025_out0;
assign v$G5_4810_out0 = v$G$AB_9585_out0 && v$P$CD_11027_out0;
assign v$G5_4900_out0 = v$G$AB_9675_out0 && v$P$CD_11117_out0;
assign v$G5_4904_out0 = v$G$AB_9679_out0 && v$P$CD_11121_out0;
assign v$G5_4923_out0 = v$G$AB_9698_out0 && v$P$CD_11140_out0;
assign v$G5_4931_out0 = v$G$AB_9706_out0 && v$P$CD_11148_out0;
assign v$G5_4933_out0 = v$G$AB_9708_out0 && v$P$CD_11150_out0;
assign v$P22_4946_out0 = v$P_14493_out0;
assign v$P22_4949_out0 = v$P_14565_out0;
assign v$G1_5270_out0 = v$G_10512_out0;
assign v$G1_5273_out0 = v$G_10584_out0;
assign v$G1_5848_out0 = v$P$AB_2249_out0 && v$P$CD_10991_out0;
assign v$G1_5857_out0 = v$P$AB_2258_out0 && v$P$CD_11000_out0;
assign v$G1_5858_out0 = v$P$AB_2259_out0 && v$P$CD_11001_out0;
assign v$G1_5869_out0 = v$P$AB_2270_out0 && v$P$CD_11012_out0;
assign v$G1_5871_out0 = v$P$AB_2272_out0 && v$P$CD_11014_out0;
assign v$G1_5878_out0 = v$P$AB_2279_out0 && v$P$CD_11021_out0;
assign v$G1_5879_out0 = v$P$AB_2280_out0 && v$P$CD_11022_out0;
assign v$G1_5971_out0 = v$P$AB_2372_out0 && v$P$CD_11114_out0;
assign v$G1_5980_out0 = v$P$AB_2381_out0 && v$P$CD_11123_out0;
assign v$G1_5981_out0 = v$P$AB_2382_out0 && v$P$CD_11124_out0;
assign v$G1_5992_out0 = v$P$AB_2393_out0 && v$P$CD_11135_out0;
assign v$G1_5994_out0 = v$P$AB_2395_out0 && v$P$CD_11137_out0;
assign v$G1_6001_out0 = v$P$AB_2402_out0 && v$P$CD_11144_out0;
assign v$G1_6002_out0 = v$P$AB_2403_out0 && v$P$CD_11145_out0;
assign v$G4_6020_out0 = v$G_10520_out0;
assign v$G4_6023_out0 = v$G_10592_out0;
assign v$P23_6627_out0 = v$P_14488_out0;
assign v$P23_6630_out0 = v$P_14560_out0;
assign v$P16_7244_out0 = v$P_14500_out0;
assign v$P16_7247_out0 = v$P_14572_out0;
assign v$G20_8534_out0 = v$G_10525_out0;
assign v$G20_8537_out0 = v$G_10597_out0;
assign v$G$AB_9509_out0 = v$G0_16549_out0;
assign v$G$AB_9512_out0 = v$G18_13509_out0;
assign v$G$AB_9513_out0 = v$G21_14627_out0;
assign v$G$AB_9525_out0 = v$G12_7328_out0;
assign v$G$AB_9527_out0 = v$G15_11542_out0;
assign v$G$AB_9530_out0 = v$G6_16971_out0;
assign v$G$AB_9536_out0 = v$G3_11603_out0;
assign v$G$AB_9541_out0 = v$G9_9256_out0;
assign v$G$AB_9632_out0 = v$G0_16552_out0;
assign v$G$AB_9635_out0 = v$G18_13512_out0;
assign v$G$AB_9636_out0 = v$G21_14630_out0;
assign v$G$AB_9648_out0 = v$G12_7331_out0;
assign v$G$AB_9650_out0 = v$G15_11545_out0;
assign v$G$AB_9653_out0 = v$G6_16974_out0;
assign v$G$AB_9659_out0 = v$G3_11606_out0;
assign v$G$AB_9664_out0 = v$G9_9259_out0;
assign v$G17_9715_out0 = v$G_10516_out0;
assign v$G17_9718_out0 = v$G_10588_out0;
assign v$P11_9993_out0 = v$P_14498_out0;
assign v$P11_9996_out0 = v$P_14570_out0;
assign v$_10819_out0 = { v$_14023_out0,v$_19276_out0 };
assign v$_10822_out0 = { v$_14026_out0,v$_19279_out0 };
assign v$P$CD_10957_out0 = v$P6_8419_out0;
assign v$P$CD_10958_out0 = v$P3_15922_out0;
assign v$P$CD_10959_out0 = v$P12_244_out0;
assign v$P$CD_10960_out0 = v$P9_19054_out0;
assign v$P$CD_10963_out0 = v$P18_12291_out0;
assign v$P$CD_10974_out0 = v$P15_7184_out0;
assign v$P$CD_10975_out0 = v$P21_4982_out0;
assign v$P$CD_11080_out0 = v$P6_8422_out0;
assign v$P$CD_11081_out0 = v$P3_15925_out0;
assign v$P$CD_11082_out0 = v$P12_247_out0;
assign v$P$CD_11083_out0 = v$P9_19057_out0;
assign v$P$CD_11086_out0 = v$P18_12294_out0;
assign v$P$CD_11097_out0 = v$P15_7187_out0;
assign v$P$CD_11098_out0 = v$P21_4985_out0;
assign v$P20_11153_out0 = v$P_14496_out0;
assign v$P20_11156_out0 = v$P_14568_out0;
assign v$G5_11171_out0 = v$G_10528_out0;
assign v$G5_11174_out0 = v$G_10600_out0;
assign v$G11_11576_out0 = v$G_10527_out0;
assign v$G11_11579_out0 = v$G_10599_out0;
assign v$P17_12329_out0 = v$P_14487_out0;
assign v$P17_12332_out0 = v$P_14559_out0;
assign v$P7_12339_out0 = v$P_14482_out0;
assign v$P7_12342_out0 = v$P_14554_out0;
assign v$G22_13105_out0 = v$G_10522_out0;
assign v$G22_13108_out0 = v$G_10594_out0;
assign v$P4_14215_out0 = v$P_14491_out0;
assign v$P4_14218_out0 = v$P_14563_out0;
assign v$G23_14921_out0 = v$G_10517_out0;
assign v$G23_14924_out0 = v$G_10589_out0;
assign v$GATE2_16356_out0 = v$CIN_16718_out0 && v$P0_5024_out0;
assign v$GATE2_16359_out0 = v$CIN_16721_out0 && v$P0_5027_out0;
assign v$G2_16569_out0 = v$G_10526_out0;
assign v$G2_16572_out0 = v$G_10598_out0;
assign v$P19_16933_out0 = v$P_14492_out0;
assign v$P19_16936_out0 = v$P_14564_out0;
assign v$G16_17072_out0 = v$G_10529_out0;
assign v$G16_17075_out0 = v$G_10601_out0;
assign v$G14_18594_out0 = v$G_10513_out0;
assign v$G14_18597_out0 = v$G_10585_out0;
assign v$GATE1_721_out0 = v$GATE2_16356_out0 || v$G0_16549_out0;
assign v$GATE1_724_out0 = v$GATE2_16359_out0 || v$G0_16552_out0;
assign v$P$AD_835_out0 = v$G1_5848_out0;
assign v$P$AD_844_out0 = v$G1_5857_out0;
assign v$P$AD_845_out0 = v$G1_5858_out0;
assign v$P$AD_856_out0 = v$G1_5869_out0;
assign v$P$AD_858_out0 = v$G1_5871_out0;
assign v$P$AD_865_out0 = v$G1_5878_out0;
assign v$P$AD_866_out0 = v$G1_5879_out0;
assign v$P$AD_958_out0 = v$G1_5971_out0;
assign v$P$AD_967_out0 = v$G1_5980_out0;
assign v$P$AD_968_out0 = v$G1_5981_out0;
assign v$P$AD_979_out0 = v$G1_5992_out0;
assign v$P$AD_981_out0 = v$G1_5994_out0;
assign v$P$AD_988_out0 = v$G1_6001_out0;
assign v$P$AD_989_out0 = v$G1_6002_out0;
assign v$G$CD_1059_out0 = v$G14_18594_out0;
assign v$G$CD_1060_out0 = v$G8_2771_out0;
assign v$G$CD_1062_out0 = v$G1_5270_out0;
assign v$G$CD_1065_out0 = v$G19_2045_out0;
assign v$G$CD_1066_out0 = v$G22_13105_out0;
assign v$G$CD_1073_out0 = v$G23_14921_out0;
assign v$G$CD_1075_out0 = v$G2_16569_out0;
assign v$G$CD_1076_out0 = v$G5_11171_out0;
assign v$G$CD_1078_out0 = v$G13_3053_out0;
assign v$G$CD_1079_out0 = v$G17_9715_out0;
assign v$G$CD_1080_out0 = v$G16_17072_out0;
assign v$G$CD_1083_out0 = v$G7_1850_out0;
assign v$G$CD_1089_out0 = v$G4_6020_out0;
assign v$G$CD_1093_out0 = v$G20_8534_out0;
assign v$G$CD_1094_out0 = v$G10_1994_out0;
assign v$G$CD_1098_out0 = v$G11_11576_out0;
assign v$G$CD_1182_out0 = v$G14_18597_out0;
assign v$G$CD_1183_out0 = v$G8_2774_out0;
assign v$G$CD_1185_out0 = v$G1_5273_out0;
assign v$G$CD_1188_out0 = v$G19_2048_out0;
assign v$G$CD_1189_out0 = v$G22_13108_out0;
assign v$G$CD_1196_out0 = v$G23_14924_out0;
assign v$G$CD_1198_out0 = v$G2_16572_out0;
assign v$G$CD_1199_out0 = v$G5_11174_out0;
assign v$G$CD_1201_out0 = v$G13_3056_out0;
assign v$G$CD_1202_out0 = v$G17_9718_out0;
assign v$G$CD_1203_out0 = v$G16_17075_out0;
assign v$G$CD_1206_out0 = v$G7_1853_out0;
assign v$G$CD_1212_out0 = v$G4_6023_out0;
assign v$G$CD_1216_out0 = v$G20_8537_out0;
assign v$G$CD_1217_out0 = v$G10_1997_out0;
assign v$G$CD_1221_out0 = v$G11_11579_out0;
assign v$COUTD_7012_out0 = v$G6_534_out0;
assign v$COUTD_7017_out0 = v$G6_539_out0;
assign v$COUTD_7023_out0 = v$G6_545_out0;
assign v$COUTD_7026_out0 = v$G6_548_out0;
assign v$COUTD_7031_out0 = v$G6_553_out0;
assign v$COUTD_7044_out0 = v$G6_566_out0;
assign v$COUTD_7135_out0 = v$G6_657_out0;
assign v$COUTD_7140_out0 = v$G6_662_out0;
assign v$COUTD_7146_out0 = v$G6_668_out0;
assign v$COUTD_7149_out0 = v$G6_671_out0;
assign v$COUTD_7154_out0 = v$G6_676_out0;
assign v$COUTD_7167_out0 = v$G6_689_out0;
assign v$P$CD_10948_out0 = v$P14_3370_out0;
assign v$P$CD_10949_out0 = v$P8_1862_out0;
assign v$P$CD_10951_out0 = v$P1_3169_out0;
assign v$P$CD_10954_out0 = v$P19_16933_out0;
assign v$P$CD_10955_out0 = v$P22_4946_out0;
assign v$P$CD_10962_out0 = v$P23_6627_out0;
assign v$P$CD_10964_out0 = v$P2_2425_out0;
assign v$P$CD_10965_out0 = v$P5_229_out0;
assign v$P$CD_10967_out0 = v$P13_3246_out0;
assign v$P$CD_10968_out0 = v$P17_12329_out0;
assign v$P$CD_10969_out0 = v$P16_7244_out0;
assign v$P$CD_10972_out0 = v$P7_12339_out0;
assign v$P$CD_10978_out0 = v$P4_14215_out0;
assign v$P$CD_10982_out0 = v$P20_11153_out0;
assign v$P$CD_10983_out0 = v$P10_361_out0;
assign v$P$CD_10987_out0 = v$P11_9993_out0;
assign v$P$CD_11071_out0 = v$P14_3373_out0;
assign v$P$CD_11072_out0 = v$P8_1865_out0;
assign v$P$CD_11074_out0 = v$P1_3172_out0;
assign v$P$CD_11077_out0 = v$P19_16936_out0;
assign v$P$CD_11078_out0 = v$P22_4949_out0;
assign v$P$CD_11085_out0 = v$P23_6630_out0;
assign v$P$CD_11087_out0 = v$P2_2428_out0;
assign v$P$CD_11088_out0 = v$P5_232_out0;
assign v$P$CD_11090_out0 = v$P13_3249_out0;
assign v$P$CD_11091_out0 = v$P17_12332_out0;
assign v$P$CD_11092_out0 = v$P16_7247_out0;
assign v$P$CD_11095_out0 = v$P7_12342_out0;
assign v$P$CD_11101_out0 = v$P4_14218_out0;
assign v$P$CD_11105_out0 = v$P20_11156_out0;
assign v$P$CD_11106_out0 = v$P10_364_out0;
assign v$P$CD_11110_out0 = v$P11_9996_out0;
assign v$G4_11698_out0 = v$G5_4777_out0 || v$G$CD_1105_out0;
assign v$G4_11702_out0 = v$G5_4781_out0 || v$G$CD_1109_out0;
assign v$G4_11721_out0 = v$G5_4800_out0 || v$G$CD_1128_out0;
assign v$G4_11729_out0 = v$G5_4808_out0 || v$G$CD_1136_out0;
assign v$G4_11731_out0 = v$G5_4810_out0 || v$G$CD_1138_out0;
assign v$G4_11821_out0 = v$G5_4900_out0 || v$G$CD_1228_out0;
assign v$G4_11825_out0 = v$G5_4904_out0 || v$G$CD_1232_out0;
assign v$G4_11844_out0 = v$G5_4923_out0 || v$G$CD_1251_out0;
assign v$G4_11852_out0 = v$G5_4931_out0 || v$G$CD_1259_out0;
assign v$G4_11854_out0 = v$G5_4933_out0 || v$G$CD_1261_out0;
assign v$G8_11970_out0 = v$CINA_8815_out0 && v$P$AB_2209_out0;
assign v$G8_11973_out0 = v$CINA_8818_out0 && v$P$AB_2212_out0;
assign v$G8_11974_out0 = v$CINA_8819_out0 && v$P$AB_2213_out0;
assign v$G8_11986_out0 = v$CINA_8831_out0 && v$P$AB_2225_out0;
assign v$G8_11988_out0 = v$CINA_8833_out0 && v$P$AB_2227_out0;
assign v$G8_11991_out0 = v$CINA_8836_out0 && v$P$AB_2230_out0;
assign v$G8_11997_out0 = v$CINA_8842_out0 && v$P$AB_2236_out0;
assign v$G8_12002_out0 = v$CINA_8847_out0 && v$P$AB_2241_out0;
assign v$G8_12093_out0 = v$CINA_8938_out0 && v$P$AB_2332_out0;
assign v$G8_12096_out0 = v$CINA_8941_out0 && v$P$AB_2335_out0;
assign v$G8_12097_out0 = v$CINA_8942_out0 && v$P$AB_2336_out0;
assign v$G8_12109_out0 = v$CINA_8954_out0 && v$P$AB_2348_out0;
assign v$G8_12111_out0 = v$CINA_8956_out0 && v$P$AB_2350_out0;
assign v$G8_12114_out0 = v$CINA_8959_out0 && v$P$AB_2353_out0;
assign v$G8_12120_out0 = v$CINA_8965_out0 && v$P$AB_2359_out0;
assign v$G8_12125_out0 = v$CINA_8970_out0 && v$P$AB_2364_out0;
assign v$C4_1415_out0 = v$COUTD_7017_out0;
assign v$C4_1418_out0 = v$COUTD_7140_out0;
assign v$P$AB_2262_out0 = v$P$AD_835_out0;
assign v$P$AB_2269_out0 = v$P$AD_835_out0;
assign v$P$AB_2273_out0 = v$P$AD_856_out0;
assign v$P$AB_2276_out0 = v$P$AD_856_out0;
assign v$P$AB_2284_out0 = v$P$AD_835_out0;
assign v$P$AB_2385_out0 = v$P$AD_958_out0;
assign v$P$AB_2392_out0 = v$P$AD_958_out0;
assign v$P$AB_2396_out0 = v$P$AD_979_out0;
assign v$P$AB_2399_out0 = v$P$AD_979_out0;
assign v$P$AB_2407_out0 = v$P$AD_958_out0;
assign v$END27_2416_out0 = v$P$AD_865_out0;
assign v$END27_2419_out0 = v$P$AD_988_out0;
assign v$END21_4506_out0 = v$P$AD_845_out0;
assign v$END21_4509_out0 = v$P$AD_968_out0;
assign v$G5_4734_out0 = v$G$AB_9509_out0 && v$P$CD_10951_out0;
assign v$G5_4737_out0 = v$G$AB_9512_out0 && v$P$CD_10954_out0;
assign v$G5_4738_out0 = v$G$AB_9513_out0 && v$P$CD_10955_out0;
assign v$G5_4750_out0 = v$G$AB_9525_out0 && v$P$CD_10967_out0;
assign v$G5_4752_out0 = v$G$AB_9527_out0 && v$P$CD_10969_out0;
assign v$G5_4755_out0 = v$G$AB_9530_out0 && v$P$CD_10972_out0;
assign v$G5_4761_out0 = v$G$AB_9536_out0 && v$P$CD_10978_out0;
assign v$G5_4766_out0 = v$G$AB_9541_out0 && v$P$CD_10983_out0;
assign v$G5_4857_out0 = v$G$AB_9632_out0 && v$P$CD_11074_out0;
assign v$G5_4860_out0 = v$G$AB_9635_out0 && v$P$CD_11077_out0;
assign v$G5_4861_out0 = v$G$AB_9636_out0 && v$P$CD_11078_out0;
assign v$G5_4873_out0 = v$G$AB_9648_out0 && v$P$CD_11090_out0;
assign v$G5_4875_out0 = v$G$AB_9650_out0 && v$P$CD_11092_out0;
assign v$G5_4878_out0 = v$G$AB_9653_out0 && v$P$CD_11095_out0;
assign v$G5_4884_out0 = v$G$AB_9659_out0 && v$P$CD_11101_out0;
assign v$G5_4889_out0 = v$G$AB_9664_out0 && v$P$CD_11106_out0;
assign v$G1_5808_out0 = v$P$AB_2209_out0 && v$P$CD_10951_out0;
assign v$G1_5811_out0 = v$P$AB_2212_out0 && v$P$CD_10954_out0;
assign v$G1_5812_out0 = v$P$AB_2213_out0 && v$P$CD_10955_out0;
assign v$G1_5824_out0 = v$P$AB_2225_out0 && v$P$CD_10967_out0;
assign v$G1_5826_out0 = v$P$AB_2227_out0 && v$P$CD_10969_out0;
assign v$G1_5829_out0 = v$P$AB_2230_out0 && v$P$CD_10972_out0;
assign v$G1_5835_out0 = v$P$AB_2236_out0 && v$P$CD_10978_out0;
assign v$G1_5840_out0 = v$P$AB_2241_out0 && v$P$CD_10983_out0;
assign v$G1_5931_out0 = v$P$AB_2332_out0 && v$P$CD_11074_out0;
assign v$G1_5934_out0 = v$P$AB_2335_out0 && v$P$CD_11077_out0;
assign v$G1_5935_out0 = v$P$AB_2336_out0 && v$P$CD_11078_out0;
assign v$G1_5947_out0 = v$P$AB_2348_out0 && v$P$CD_11090_out0;
assign v$G1_5949_out0 = v$P$AB_2350_out0 && v$P$CD_11092_out0;
assign v$G1_5952_out0 = v$P$AB_2353_out0 && v$P$CD_11095_out0;
assign v$G1_5958_out0 = v$P$AB_2359_out0 && v$P$CD_11101_out0;
assign v$G1_5963_out0 = v$P$AB_2364_out0 && v$P$CD_11106_out0;
assign v$END40_6064_out0 = v$COUTD_7031_out0;
assign v$END40_6067_out0 = v$COUTD_7154_out0;
assign v$END29_6163_out0 = v$P$AD_856_out0;
assign v$END29_6166_out0 = v$P$AD_979_out0;
assign v$CINA_8858_out0 = v$COUTD_7044_out0;
assign v$CINA_8862_out0 = v$COUTD_7044_out0;
assign v$CINA_8881_out0 = v$COUTD_7044_out0;
assign v$CINA_8889_out0 = v$COUTD_7031_out0;
assign v$CINA_8891_out0 = v$COUTD_7044_out0;
assign v$CINA_8981_out0 = v$COUTD_7167_out0;
assign v$CINA_8985_out0 = v$COUTD_7167_out0;
assign v$CINA_9004_out0 = v$COUTD_7167_out0;
assign v$CINA_9012_out0 = v$COUTD_7154_out0;
assign v$CINA_9014_out0 = v$COUTD_7167_out0;
assign v$END4_9739_out0 = v$COUTD_7012_out0;
assign v$END4_9742_out0 = v$COUTD_7135_out0;
assign v$G7_10062_out0 = v$G8_11970_out0 && v$P$CD_10951_out0;
assign v$G7_10065_out0 = v$G8_11973_out0 && v$P$CD_10954_out0;
assign v$G7_10066_out0 = v$G8_11974_out0 && v$P$CD_10955_out0;
assign v$G7_10078_out0 = v$G8_11986_out0 && v$P$CD_10967_out0;
assign v$G7_10080_out0 = v$G8_11988_out0 && v$P$CD_10969_out0;
assign v$G7_10083_out0 = v$G8_11991_out0 && v$P$CD_10972_out0;
assign v$G7_10089_out0 = v$G8_11997_out0 && v$P$CD_10978_out0;
assign v$G7_10094_out0 = v$G8_12002_out0 && v$P$CD_10983_out0;
assign v$G7_10185_out0 = v$G8_12093_out0 && v$P$CD_11074_out0;
assign v$G7_10188_out0 = v$G8_12096_out0 && v$P$CD_11077_out0;
assign v$G7_10189_out0 = v$G8_12097_out0 && v$P$CD_11078_out0;
assign v$G7_10201_out0 = v$G8_12109_out0 && v$P$CD_11090_out0;
assign v$G7_10203_out0 = v$G8_12111_out0 && v$P$CD_11092_out0;
assign v$G7_10206_out0 = v$G8_12114_out0 && v$P$CD_11095_out0;
assign v$G7_10212_out0 = v$G8_12120_out0 && v$P$CD_11101_out0;
assign v$G7_10217_out0 = v$G8_12125_out0 && v$P$CD_11106_out0;
assign v$C0_11189_out0 = v$GATE1_721_out0;
assign v$C0_11192_out0 = v$GATE1_724_out0;
assign v$END52_12551_out0 = v$P$AD_858_out0;
assign v$END52_12554_out0 = v$P$AD_981_out0;
assign v$END60_15743_out0 = v$COUTD_7026_out0;
assign v$END60_15746_out0 = v$COUTD_7149_out0;
assign v$C3_16325_out0 = v$COUTD_7023_out0;
assign v$C3_16328_out0 = v$COUTD_7146_out0;
assign v$C5_16521_out0 = v$COUTD_7044_out0;
assign v$C5_16524_out0 = v$COUTD_7167_out0;
assign v$END23_17338_out0 = v$P$AD_866_out0;
assign v$END23_17341_out0 = v$P$AD_989_out0;
assign v$END25_17668_out0 = v$P$AD_844_out0;
assign v$END25_17671_out0 = v$P$AD_967_out0;
assign v$G$AD_17772_out0 = v$G4_11698_out0;
assign v$G$AD_17776_out0 = v$G4_11702_out0;
assign v$G$AD_17795_out0 = v$G4_11721_out0;
assign v$G$AD_17803_out0 = v$G4_11729_out0;
assign v$G$AD_17805_out0 = v$G4_11731_out0;
assign v$G$AD_17895_out0 = v$G4_11821_out0;
assign v$G$AD_17899_out0 = v$G4_11825_out0;
assign v$G$AD_17918_out0 = v$G4_11844_out0;
assign v$G$AD_17926_out0 = v$G4_11852_out0;
assign v$G$AD_17928_out0 = v$G4_11854_out0;
assign v$END16_224_out0 = v$G$AD_17805_out0;
assign v$END16_227_out0 = v$G$AD_17928_out0;
assign v$END14_286_out0 = v$G$AD_17776_out0;
assign v$END14_289_out0 = v$G$AD_17899_out0;
assign v$P$AD_795_out0 = v$G1_5808_out0;
assign v$P$AD_798_out0 = v$G1_5811_out0;
assign v$P$AD_799_out0 = v$G1_5812_out0;
assign v$P$AD_811_out0 = v$G1_5824_out0;
assign v$P$AD_813_out0 = v$G1_5826_out0;
assign v$P$AD_816_out0 = v$G1_5829_out0;
assign v$P$AD_822_out0 = v$G1_5835_out0;
assign v$P$AD_827_out0 = v$G1_5840_out0;
assign v$P$AD_918_out0 = v$G1_5931_out0;
assign v$P$AD_921_out0 = v$G1_5934_out0;
assign v$P$AD_922_out0 = v$G1_5935_out0;
assign v$P$AD_934_out0 = v$G1_5947_out0;
assign v$P$AD_936_out0 = v$G1_5949_out0;
assign v$P$AD_939_out0 = v$G1_5952_out0;
assign v$P$AD_945_out0 = v$G1_5958_out0;
assign v$P$AD_950_out0 = v$G1_5963_out0;
assign v$G$CD_1125_out0 = v$G$AD_17803_out0;
assign v$G$CD_1248_out0 = v$G$AD_17926_out0;
assign {v$A2A_1789_out1,v$A2A_1789_out0 } = v$A1_1870_out0 + v$B1_8427_out0 + v$C0_11189_out0;
assign {v$A2A_1792_out1,v$A2A_1792_out0 } = v$A1_1873_out0 + v$B1_8430_out0 + v$C0_11192_out0;
assign {v$A7A_1817_out1,v$A7A_1817_out0 } = v$A5_6903_out0 + v$B5_18980_out0 + v$C4_1415_out0;
assign {v$A7A_1820_out1,v$A7A_1820_out0 } = v$A5_6906_out0 + v$B5_18983_out0 + v$C4_1418_out0;
assign v$C4_2040_out0 = v$C4_1415_out0;
assign v$C4_2043_out0 = v$C4_1418_out0;
assign {v$A6A_3336_out1,v$A6A_3336_out0 } = v$A6_322_out0 + v$B6_13885_out0 + v$C5_16521_out0;
assign {v$A6A_3339_out1,v$A6A_3339_out0 } = v$A6_325_out0 + v$B6_13888_out0 + v$C5_16524_out0;
assign v$G1_5861_out0 = v$P$AB_2262_out0 && v$P$CD_11004_out0;
assign v$G1_5868_out0 = v$P$AB_2269_out0 && v$P$CD_11011_out0;
assign v$G1_5872_out0 = v$P$AB_2273_out0 && v$P$CD_11015_out0;
assign v$G1_5875_out0 = v$P$AB_2276_out0 && v$P$CD_11018_out0;
assign v$G1_5883_out0 = v$P$AB_2284_out0 && v$P$CD_11026_out0;
assign v$G1_5984_out0 = v$P$AB_2385_out0 && v$P$CD_11127_out0;
assign v$G1_5991_out0 = v$P$AB_2392_out0 && v$P$CD_11134_out0;
assign v$G1_5995_out0 = v$P$AB_2396_out0 && v$P$CD_11138_out0;
assign v$G1_5998_out0 = v$P$AB_2399_out0 && v$P$CD_11141_out0;
assign v$G1_6006_out0 = v$P$AB_2407_out0 && v$P$CD_11149_out0;
assign v$G$AB_9549_out0 = v$G$AD_17795_out0;
assign v$G$AB_9558_out0 = v$G$AD_17795_out0;
assign v$G$AB_9559_out0 = v$G$AD_17772_out0;
assign v$G$AB_9570_out0 = v$G$AD_17795_out0;
assign v$G$AB_9572_out0 = v$G$AD_17795_out0;
assign v$G$AB_9579_out0 = v$G$AD_17795_out0;
assign v$G$AB_9580_out0 = v$G$AD_17772_out0;
assign v$G$AB_9672_out0 = v$G$AD_17918_out0;
assign v$G$AB_9681_out0 = v$G$AD_17918_out0;
assign v$G$AB_9682_out0 = v$G$AD_17895_out0;
assign v$G$AB_9693_out0 = v$G$AD_17918_out0;
assign v$G$AB_9695_out0 = v$G$AD_17918_out0;
assign v$G$AB_9702_out0 = v$G$AD_17918_out0;
assign v$G$AB_9703_out0 = v$G$AD_17895_out0;
assign v$C0_9746_out0 = v$C0_11189_out0;
assign v$C0_9749_out0 = v$C0_11192_out0;
assign v$G4_11655_out0 = v$G5_4734_out0 || v$G$CD_1062_out0;
assign v$G4_11658_out0 = v$G5_4737_out0 || v$G$CD_1065_out0;
assign v$G4_11659_out0 = v$G5_4738_out0 || v$G$CD_1066_out0;
assign v$G4_11671_out0 = v$G5_4750_out0 || v$G$CD_1078_out0;
assign v$G4_11673_out0 = v$G5_4752_out0 || v$G$CD_1080_out0;
assign v$G4_11676_out0 = v$G5_4755_out0 || v$G$CD_1083_out0;
assign v$G4_11682_out0 = v$G5_4761_out0 || v$G$CD_1089_out0;
assign v$G4_11687_out0 = v$G5_4766_out0 || v$G$CD_1094_out0;
assign v$G4_11778_out0 = v$G5_4857_out0 || v$G$CD_1185_out0;
assign v$G4_11781_out0 = v$G5_4860_out0 || v$G$CD_1188_out0;
assign v$G4_11782_out0 = v$G5_4861_out0 || v$G$CD_1189_out0;
assign v$G4_11794_out0 = v$G5_4873_out0 || v$G$CD_1201_out0;
assign v$G4_11796_out0 = v$G5_4875_out0 || v$G$CD_1203_out0;
assign v$G4_11799_out0 = v$G5_4878_out0 || v$G$CD_1206_out0;
assign v$G4_11805_out0 = v$G5_4884_out0 || v$G$CD_1212_out0;
assign v$G4_11810_out0 = v$G5_4889_out0 || v$G$CD_1217_out0;
assign v$G8_12013_out0 = v$CINA_8858_out0 && v$P$AB_2252_out0;
assign v$G8_12017_out0 = v$CINA_8862_out0 && v$P$AB_2256_out0;
assign v$G8_12036_out0 = v$CINA_8881_out0 && v$P$AB_2275_out0;
assign v$G8_12044_out0 = v$CINA_8889_out0 && v$P$AB_2283_out0;
assign v$G8_12046_out0 = v$CINA_8891_out0 && v$P$AB_2285_out0;
assign v$G8_12136_out0 = v$CINA_8981_out0 && v$P$AB_2375_out0;
assign v$G8_12140_out0 = v$CINA_8985_out0 && v$P$AB_2379_out0;
assign v$G8_12159_out0 = v$CINA_9004_out0 && v$P$AB_2398_out0;
assign v$G8_12167_out0 = v$CINA_9012_out0 && v$P$AB_2406_out0;
assign v$G8_12169_out0 = v$CINA_9014_out0 && v$P$AB_2408_out0;
assign v$C5_12255_out0 = v$C5_16521_out0;
assign v$C5_12258_out0 = v$C5_16524_out0;
assign v$END18_12521_out0 = v$G$AD_17772_out0;
assign v$END18_12524_out0 = v$G$AD_17895_out0;
assign v$C3_16422_out0 = v$C3_16325_out0;
assign v$C3_16425_out0 = v$C3_16328_out0;
assign {v$A5A_16711_out1,v$A5A_16711_out0 } = v$A4_18140_out0 + v$B4_15268_out0 + v$C3_16325_out0;
assign {v$A5A_16714_out1,v$A5A_16714_out0 } = v$A4_18143_out0 + v$B4_15271_out0 + v$C3_16328_out0;
assign v$_84_out0 = { v$A5A_16711_out0,v$A7A_1817_out0 };
assign v$_87_out0 = { v$A5A_16714_out0,v$A7A_1820_out0 };
assign v$G6_497_out0 = v$G4_11655_out0 || v$G7_10062_out0;
assign v$G6_500_out0 = v$G4_11658_out0 || v$G7_10065_out0;
assign v$G6_501_out0 = v$G4_11659_out0 || v$G7_10066_out0;
assign v$G6_513_out0 = v$G4_11671_out0 || v$G7_10078_out0;
assign v$G6_515_out0 = v$G4_11673_out0 || v$G7_10080_out0;
assign v$G6_518_out0 = v$G4_11676_out0 || v$G7_10083_out0;
assign v$G6_524_out0 = v$G4_11682_out0 || v$G7_10089_out0;
assign v$G6_529_out0 = v$G4_11687_out0 || v$G7_10094_out0;
assign v$G6_620_out0 = v$G4_11778_out0 || v$G7_10185_out0;
assign v$G6_623_out0 = v$G4_11781_out0 || v$G7_10188_out0;
assign v$G6_624_out0 = v$G4_11782_out0 || v$G7_10189_out0;
assign v$G6_636_out0 = v$G4_11794_out0 || v$G7_10201_out0;
assign v$G6_638_out0 = v$G4_11796_out0 || v$G7_10203_out0;
assign v$G6_641_out0 = v$G4_11799_out0 || v$G7_10206_out0;
assign v$G6_647_out0 = v$G4_11805_out0 || v$G7_10212_out0;
assign v$G6_652_out0 = v$G4_11810_out0 || v$G7_10217_out0;
assign v$P$AD_848_out0 = v$G1_5861_out0;
assign v$P$AD_855_out0 = v$G1_5868_out0;
assign v$P$AD_859_out0 = v$G1_5872_out0;
assign v$P$AD_862_out0 = v$G1_5875_out0;
assign v$P$AD_870_out0 = v$G1_5883_out0;
assign v$P$AD_971_out0 = v$G1_5984_out0;
assign v$P$AD_978_out0 = v$G1_5991_out0;
assign v$P$AD_982_out0 = v$G1_5995_out0;
assign v$P$AD_985_out0 = v$G1_5998_out0;
assign v$P$AD_993_out0 = v$G1_6006_out0;
assign v$END1_1698_out0 = v$A2A_1789_out1;
assign v$END1_1701_out0 = v$A2A_1792_out1;
assign v$P$AB_2206_out0 = v$P$AD_811_out0;
assign v$P$AB_2207_out0 = v$P$AD_816_out0;
assign v$P$AB_2220_out0 = v$P$AD_799_out0;
assign v$P$AB_2222_out0 = v$P$AD_795_out0;
assign v$P$AB_2223_out0 = v$P$AD_822_out0;
assign v$P$AB_2226_out0 = v$P$AD_813_out0;
assign v$P$AB_2240_out0 = v$P$AD_798_out0;
assign v$P$AB_2245_out0 = v$P$AD_827_out0;
assign v$P$AB_2329_out0 = v$P$AD_934_out0;
assign v$P$AB_2330_out0 = v$P$AD_939_out0;
assign v$P$AB_2343_out0 = v$P$AD_922_out0;
assign v$P$AB_2345_out0 = v$P$AD_918_out0;
assign v$P$AB_2346_out0 = v$P$AD_945_out0;
assign v$P$AB_2349_out0 = v$P$AD_936_out0;
assign v$P$AB_2363_out0 = v$P$AD_921_out0;
assign v$P$AB_2368_out0 = v$P$AD_950_out0;
assign v$_2648_out0 = { v$C4_2040_out0,v$C5_12255_out0 };
assign v$_2651_out0 = { v$C4_2043_out0,v$C5_12258_out0 };
assign v$END5_4303_out0 = v$A7A_1817_out1;
assign v$END5_4306_out0 = v$A7A_1820_out1;
assign v$G5_4774_out0 = v$G$AB_9549_out0 && v$P$CD_10991_out0;
assign v$G5_4783_out0 = v$G$AB_9558_out0 && v$P$CD_11000_out0;
assign v$G5_4784_out0 = v$G$AB_9559_out0 && v$P$CD_11001_out0;
assign v$G5_4795_out0 = v$G$AB_9570_out0 && v$P$CD_11012_out0;
assign v$G5_4797_out0 = v$G$AB_9572_out0 && v$P$CD_11014_out0;
assign v$G5_4804_out0 = v$G$AB_9579_out0 && v$P$CD_11021_out0;
assign v$G5_4805_out0 = v$G$AB_9580_out0 && v$P$CD_11022_out0;
assign v$G5_4897_out0 = v$G$AB_9672_out0 && v$P$CD_11114_out0;
assign v$G5_4906_out0 = v$G$AB_9681_out0 && v$P$CD_11123_out0;
assign v$G5_4907_out0 = v$G$AB_9682_out0 && v$P$CD_11124_out0;
assign v$G5_4918_out0 = v$G$AB_9693_out0 && v$P$CD_11135_out0;
assign v$G5_4920_out0 = v$G$AB_9695_out0 && v$P$CD_11137_out0;
assign v$G5_4927_out0 = v$G$AB_9702_out0 && v$P$CD_11144_out0;
assign v$G5_4928_out0 = v$G$AB_9703_out0 && v$P$CD_11145_out0;
assign v$END4_5465_out0 = v$A5A_16711_out1;
assign v$END4_5468_out0 = v$A5A_16714_out1;
assign v$G7_10105_out0 = v$G8_12013_out0 && v$P$CD_10994_out0;
assign v$G7_10109_out0 = v$G8_12017_out0 && v$P$CD_10998_out0;
assign v$G7_10128_out0 = v$G8_12036_out0 && v$P$CD_11017_out0;
assign v$G7_10136_out0 = v$G8_12044_out0 && v$P$CD_11025_out0;
assign v$G7_10138_out0 = v$G8_12046_out0 && v$P$CD_11027_out0;
assign v$G7_10228_out0 = v$G8_12136_out0 && v$P$CD_11117_out0;
assign v$G7_10232_out0 = v$G8_12140_out0 && v$P$CD_11121_out0;
assign v$G7_10251_out0 = v$G8_12159_out0 && v$P$CD_11140_out0;
assign v$G7_10259_out0 = v$G8_12167_out0 && v$P$CD_11148_out0;
assign v$G7_10261_out0 = v$G8_12169_out0 && v$P$CD_11150_out0;
assign v$P$CD_10952_out0 = v$P$AD_822_out0;
assign v$P$CD_10956_out0 = v$P$AD_799_out0;
assign v$P$CD_10977_out0 = v$P$AD_813_out0;
assign v$P$CD_10980_out0 = v$P$AD_811_out0;
assign v$P$CD_10981_out0 = v$P$AD_827_out0;
assign v$P$CD_10985_out0 = v$P$AD_798_out0;
assign v$P$CD_10986_out0 = v$P$AD_816_out0;
assign v$P$CD_11075_out0 = v$P$AD_945_out0;
assign v$P$CD_11079_out0 = v$P$AD_922_out0;
assign v$P$CD_11100_out0 = v$P$AD_936_out0;
assign v$P$CD_11103_out0 = v$P$AD_934_out0;
assign v$P$CD_11104_out0 = v$P$AD_950_out0;
assign v$P$CD_11108_out0 = v$P$AD_921_out0;
assign v$P$CD_11109_out0 = v$P$AD_939_out0;
assign v$_14022_out0 = { v$A1A_12225_out0,v$A2A_1789_out0 };
assign v$_14025_out0 = { v$A1A_12228_out0,v$A2A_1792_out0 };
assign v$_15616_out0 = { v$C2_18779_out0,v$C3_16422_out0 };
assign v$_15619_out0 = { v$C2_18782_out0,v$C3_16425_out0 };
assign v$END6_15833_out0 = v$A6A_3336_out1;
assign v$END6_15836_out0 = v$A6A_3339_out1;
assign v$G$AD_17729_out0 = v$G4_11655_out0;
assign v$G$AD_17732_out0 = v$G4_11658_out0;
assign v$G$AD_17733_out0 = v$G4_11659_out0;
assign v$G$AD_17745_out0 = v$G4_11671_out0;
assign v$G$AD_17747_out0 = v$G4_11673_out0;
assign v$G$AD_17750_out0 = v$G4_11676_out0;
assign v$G$AD_17756_out0 = v$G4_11682_out0;
assign v$G$AD_17761_out0 = v$G4_11687_out0;
assign v$G$AD_17852_out0 = v$G4_11778_out0;
assign v$G$AD_17855_out0 = v$G4_11781_out0;
assign v$G$AD_17856_out0 = v$G4_11782_out0;
assign v$G$AD_17868_out0 = v$G4_11794_out0;
assign v$G$AD_17870_out0 = v$G4_11796_out0;
assign v$G$AD_17873_out0 = v$G4_11799_out0;
assign v$G$AD_17879_out0 = v$G4_11805_out0;
assign v$G$AD_17884_out0 = v$G4_11810_out0;
assign v$END33_275_out0 = v$P$AD_862_out0;
assign v$END33_278_out0 = v$P$AD_985_out0;
assign v$G6_540_out0 = v$G4_11698_out0 || v$G7_10105_out0;
assign v$G6_544_out0 = v$G4_11702_out0 || v$G7_10109_out0;
assign v$G6_563_out0 = v$G4_11721_out0 || v$G7_10128_out0;
assign v$G6_571_out0 = v$G4_11729_out0 || v$G7_10136_out0;
assign v$G6_573_out0 = v$G4_11731_out0 || v$G7_10138_out0;
assign v$G6_663_out0 = v$G4_11821_out0 || v$G7_10228_out0;
assign v$G6_667_out0 = v$G4_11825_out0 || v$G7_10232_out0;
assign v$G6_686_out0 = v$G4_11844_out0 || v$G7_10251_out0;
assign v$G6_694_out0 = v$G4_11852_out0 || v$G7_10259_out0;
assign v$G6_696_out0 = v$G4_11854_out0 || v$G7_10261_out0;
assign v$G$CD_1063_out0 = v$G$AD_17756_out0;
assign v$G$CD_1067_out0 = v$G$AD_17733_out0;
assign v$G$CD_1088_out0 = v$G$AD_17747_out0;
assign v$G$CD_1091_out0 = v$G$AD_17745_out0;
assign v$G$CD_1092_out0 = v$G$AD_17761_out0;
assign v$G$CD_1096_out0 = v$G$AD_17732_out0;
assign v$G$CD_1097_out0 = v$G$AD_17750_out0;
assign v$G$CD_1186_out0 = v$G$AD_17879_out0;
assign v$G$CD_1190_out0 = v$G$AD_17856_out0;
assign v$G$CD_1211_out0 = v$G$AD_17870_out0;
assign v$G$CD_1214_out0 = v$G$AD_17868_out0;
assign v$G$CD_1215_out0 = v$G$AD_17884_out0;
assign v$G$CD_1219_out0 = v$G$AD_17855_out0;
assign v$G$CD_1220_out0 = v$G$AD_17873_out0;
assign v$P$AB_2255_out0 = v$P$AD_855_out0;
assign v$P$AB_2274_out0 = v$P$AD_855_out0;
assign v$P$AB_2378_out0 = v$P$AD_978_out0;
assign v$P$AB_2397_out0 = v$P$AD_978_out0;
assign v$END47_2878_out0 = v$P$AD_855_out0;
assign v$END47_2881_out0 = v$P$AD_978_out0;
assign v$G1_5805_out0 = v$P$AB_2206_out0 && v$P$CD_10948_out0;
assign v$G1_5806_out0 = v$P$AB_2207_out0 && v$P$CD_10949_out0;
assign v$G1_5819_out0 = v$P$AB_2220_out0 && v$P$CD_10962_out0;
assign v$G1_5821_out0 = v$P$AB_2222_out0 && v$P$CD_10964_out0;
assign v$G1_5822_out0 = v$P$AB_2223_out0 && v$P$CD_10965_out0;
assign v$G1_5825_out0 = v$P$AB_2226_out0 && v$P$CD_10968_out0;
assign v$G1_5839_out0 = v$P$AB_2240_out0 && v$P$CD_10982_out0;
assign v$G1_5844_out0 = v$P$AB_2245_out0 && v$P$CD_10987_out0;
assign v$G1_5928_out0 = v$P$AB_2329_out0 && v$P$CD_11071_out0;
assign v$G1_5929_out0 = v$P$AB_2330_out0 && v$P$CD_11072_out0;
assign v$G1_5942_out0 = v$P$AB_2343_out0 && v$P$CD_11085_out0;
assign v$G1_5944_out0 = v$P$AB_2345_out0 && v$P$CD_11087_out0;
assign v$G1_5945_out0 = v$P$AB_2346_out0 && v$P$CD_11088_out0;
assign v$G1_5948_out0 = v$P$AB_2349_out0 && v$P$CD_11091_out0;
assign v$G1_5962_out0 = v$P$AB_2363_out0 && v$P$CD_11105_out0;
assign v$G1_5967_out0 = v$P$AB_2368_out0 && v$P$CD_11110_out0;
assign v$COUTD_6975_out0 = v$G6_497_out0;
assign v$COUTD_6978_out0 = v$G6_500_out0;
assign v$COUTD_6979_out0 = v$G6_501_out0;
assign v$COUTD_6991_out0 = v$G6_513_out0;
assign v$COUTD_6993_out0 = v$G6_515_out0;
assign v$COUTD_6996_out0 = v$G6_518_out0;
assign v$COUTD_7002_out0 = v$G6_524_out0;
assign v$COUTD_7007_out0 = v$G6_529_out0;
assign v$COUTD_7098_out0 = v$G6_620_out0;
assign v$COUTD_7101_out0 = v$G6_623_out0;
assign v$COUTD_7102_out0 = v$G6_624_out0;
assign v$COUTD_7114_out0 = v$G6_636_out0;
assign v$COUTD_7116_out0 = v$G6_638_out0;
assign v$COUTD_7119_out0 = v$G6_641_out0;
assign v$COUTD_7125_out0 = v$G6_647_out0;
assign v$COUTD_7130_out0 = v$G6_652_out0;
assign v$_7570_out0 = { v$_9237_out0,v$_15616_out0 };
assign v$_7573_out0 = { v$_9240_out0,v$_15619_out0 };
assign v$G$AB_9506_out0 = v$G$AD_17745_out0;
assign v$G$AB_9507_out0 = v$G$AD_17750_out0;
assign v$G$AB_9520_out0 = v$G$AD_17733_out0;
assign v$G$AB_9522_out0 = v$G$AD_17729_out0;
assign v$G$AB_9523_out0 = v$G$AD_17756_out0;
assign v$G$AB_9526_out0 = v$G$AD_17747_out0;
assign v$G$AB_9540_out0 = v$G$AD_17732_out0;
assign v$G$AB_9545_out0 = v$G$AD_17761_out0;
assign v$G$AB_9629_out0 = v$G$AD_17868_out0;
assign v$G$AB_9630_out0 = v$G$AD_17873_out0;
assign v$G$AB_9643_out0 = v$G$AD_17856_out0;
assign v$G$AB_9645_out0 = v$G$AD_17852_out0;
assign v$G$AB_9646_out0 = v$G$AD_17879_out0;
assign v$G$AB_9649_out0 = v$G$AD_17870_out0;
assign v$G$AB_9663_out0 = v$G$AD_17855_out0;
assign v$G$AB_9668_out0 = v$G$AD_17884_out0;
assign v$G4_11695_out0 = v$G5_4774_out0 || v$G$CD_1102_out0;
assign v$G4_11704_out0 = v$G5_4783_out0 || v$G$CD_1111_out0;
assign v$G4_11705_out0 = v$G5_4784_out0 || v$G$CD_1112_out0;
assign v$G4_11716_out0 = v$G5_4795_out0 || v$G$CD_1123_out0;
assign v$G4_11718_out0 = v$G5_4797_out0 || v$G$CD_1125_out0;
assign v$G4_11725_out0 = v$G5_4804_out0 || v$G$CD_1132_out0;
assign v$G4_11726_out0 = v$G5_4805_out0 || v$G$CD_1133_out0;
assign v$G4_11818_out0 = v$G5_4897_out0 || v$G$CD_1225_out0;
assign v$G4_11827_out0 = v$G5_4906_out0 || v$G$CD_1234_out0;
assign v$G4_11828_out0 = v$G5_4907_out0 || v$G$CD_1235_out0;
assign v$G4_11839_out0 = v$G5_4918_out0 || v$G$CD_1246_out0;
assign v$G4_11841_out0 = v$G5_4920_out0 || v$G$CD_1248_out0;
assign v$G4_11848_out0 = v$G5_4927_out0 || v$G$CD_1255_out0;
assign v$G4_11849_out0 = v$G5_4928_out0 || v$G$CD_1256_out0;
assign v$END44_16260_out0 = v$P$AD_870_out0;
assign v$END44_16263_out0 = v$P$AD_993_out0;
assign v$END42_18918_out0 = v$P$AD_848_out0;
assign v$END42_18921_out0 = v$P$AD_971_out0;
assign v$END31_19133_out0 = v$P$AD_859_out0;
assign v$END31_19136_out0 = v$P$AD_982_out0;
assign v$P$AD_792_out0 = v$G1_5805_out0;
assign v$P$AD_793_out0 = v$G1_5806_out0;
assign v$P$AD_806_out0 = v$G1_5819_out0;
assign v$P$AD_808_out0 = v$G1_5821_out0;
assign v$P$AD_809_out0 = v$G1_5822_out0;
assign v$P$AD_812_out0 = v$G1_5825_out0;
assign v$P$AD_826_out0 = v$G1_5839_out0;
assign v$P$AD_831_out0 = v$G1_5844_out0;
assign v$P$AD_915_out0 = v$G1_5928_out0;
assign v$P$AD_916_out0 = v$G1_5929_out0;
assign v$P$AD_929_out0 = v$G1_5942_out0;
assign v$P$AD_931_out0 = v$G1_5944_out0;
assign v$P$AD_932_out0 = v$G1_5945_out0;
assign v$P$AD_935_out0 = v$G1_5948_out0;
assign v$P$AD_949_out0 = v$G1_5962_out0;
assign v$P$AD_954_out0 = v$G1_5967_out0;
assign v$G5_4731_out0 = v$G$AB_9506_out0 && v$P$CD_10948_out0;
assign v$G5_4732_out0 = v$G$AB_9507_out0 && v$P$CD_10949_out0;
assign v$G5_4745_out0 = v$G$AB_9520_out0 && v$P$CD_10962_out0;
assign v$G5_4747_out0 = v$G$AB_9522_out0 && v$P$CD_10964_out0;
assign v$G5_4748_out0 = v$G$AB_9523_out0 && v$P$CD_10965_out0;
assign v$G5_4751_out0 = v$G$AB_9526_out0 && v$P$CD_10968_out0;
assign v$G5_4765_out0 = v$G$AB_9540_out0 && v$P$CD_10982_out0;
assign v$G5_4770_out0 = v$G$AB_9545_out0 && v$P$CD_10987_out0;
assign v$G5_4854_out0 = v$G$AB_9629_out0 && v$P$CD_11071_out0;
assign v$G5_4855_out0 = v$G$AB_9630_out0 && v$P$CD_11072_out0;
assign v$G5_4868_out0 = v$G$AB_9643_out0 && v$P$CD_11085_out0;
assign v$G5_4870_out0 = v$G$AB_9645_out0 && v$P$CD_11087_out0;
assign v$G5_4871_out0 = v$G$AB_9646_out0 && v$P$CD_11088_out0;
assign v$G5_4874_out0 = v$G$AB_9649_out0 && v$P$CD_11091_out0;
assign v$G5_4888_out0 = v$G$AB_9663_out0 && v$P$CD_11105_out0;
assign v$G5_4893_out0 = v$G$AB_9668_out0 && v$P$CD_11110_out0;
assign v$G1_5854_out0 = v$P$AB_2255_out0 && v$P$CD_10997_out0;
assign v$G1_5873_out0 = v$P$AB_2274_out0 && v$P$CD_11016_out0;
assign v$G1_5977_out0 = v$P$AB_2378_out0 && v$P$CD_11120_out0;
assign v$G1_5996_out0 = v$P$AB_2397_out0 && v$P$CD_11139_out0;
assign v$COUTD_7018_out0 = v$G6_540_out0;
assign v$COUTD_7022_out0 = v$G6_544_out0;
assign v$COUTD_7041_out0 = v$G6_563_out0;
assign v$COUTD_7049_out0 = v$G6_571_out0;
assign v$COUTD_7051_out0 = v$G6_573_out0;
assign v$COUTD_7141_out0 = v$G6_663_out0;
assign v$COUTD_7145_out0 = v$G6_667_out0;
assign v$COUTD_7164_out0 = v$G6_686_out0;
assign v$COUTD_7172_out0 = v$G6_694_out0;
assign v$COUTD_7174_out0 = v$G6_696_out0;
assign v$CINA_8812_out0 = v$COUTD_6991_out0;
assign v$CINA_8813_out0 = v$COUTD_6996_out0;
assign v$CINA_8826_out0 = v$COUTD_6979_out0;
assign v$CINA_8828_out0 = v$COUTD_6975_out0;
assign v$CINA_8829_out0 = v$COUTD_7002_out0;
assign v$CINA_8832_out0 = v$COUTD_6993_out0;
assign v$CINA_8846_out0 = v$COUTD_6978_out0;
assign v$CINA_8851_out0 = v$COUTD_7007_out0;
assign v$CINA_8935_out0 = v$COUTD_7114_out0;
assign v$CINA_8936_out0 = v$COUTD_7119_out0;
assign v$CINA_8949_out0 = v$COUTD_7102_out0;
assign v$CINA_8951_out0 = v$COUTD_7098_out0;
assign v$CINA_8952_out0 = v$COUTD_7125_out0;
assign v$CINA_8955_out0 = v$COUTD_7116_out0;
assign v$CINA_8969_out0 = v$COUTD_7101_out0;
assign v$CINA_8974_out0 = v$COUTD_7130_out0;
assign v$C1_17402_out0 = v$COUTD_6975_out0;
assign v$C1_17405_out0 = v$COUTD_7098_out0;
assign v$G$AD_17769_out0 = v$G4_11695_out0;
assign v$G$AD_17778_out0 = v$G4_11704_out0;
assign v$G$AD_17779_out0 = v$G4_11705_out0;
assign v$G$AD_17790_out0 = v$G4_11716_out0;
assign v$G$AD_17792_out0 = v$G4_11718_out0;
assign v$G$AD_17799_out0 = v$G4_11725_out0;
assign v$G$AD_17800_out0 = v$G4_11726_out0;
assign v$G$AD_17892_out0 = v$G4_11818_out0;
assign v$G$AD_17901_out0 = v$G4_11827_out0;
assign v$G$AD_17902_out0 = v$G4_11828_out0;
assign v$G$AD_17913_out0 = v$G4_11839_out0;
assign v$G$AD_17915_out0 = v$G4_11841_out0;
assign v$G$AD_17922_out0 = v$G4_11848_out0;
assign v$G$AD_17923_out0 = v$G4_11849_out0;
assign v$END53_332_out0 = v$G$AD_17792_out0;
assign v$END53_335_out0 = v$G$AD_17915_out0;
assign v$P$AD_841_out0 = v$G1_5854_out0;
assign v$P$AD_860_out0 = v$G1_5873_out0;
assign v$P$AD_964_out0 = v$G1_5977_out0;
assign v$P$AD_983_out0 = v$G1_5996_out0;
assign v$P$AB_2205_out0 = v$P$AD_793_out0;
assign v$P$AB_2210_out0 = v$P$AD_808_out0;
assign v$P$AB_2216_out0 = v$P$AD_808_out0;
assign v$P$AB_2219_out0 = v$P$AD_826_out0;
assign v$P$AB_2224_out0 = v$P$AD_792_out0;
assign v$P$AB_2237_out0 = v$P$AD_808_out0;
assign v$P$AB_2328_out0 = v$P$AD_916_out0;
assign v$P$AB_2333_out0 = v$P$AD_931_out0;
assign v$P$AB_2339_out0 = v$P$AD_931_out0;
assign v$P$AB_2342_out0 = v$P$AD_949_out0;
assign v$P$AB_2347_out0 = v$P$AD_915_out0;
assign v$P$AB_2360_out0 = v$P$AD_931_out0;
assign v$END26_6680_out0 = v$G$AD_17799_out0;
assign v$END26_6683_out0 = v$G$AD_17922_out0;
assign v$C8_7750_out0 = v$COUTD_7018_out0;
assign v$C8_7753_out0 = v$COUTD_7141_out0;
assign v$CINA_8855_out0 = v$COUTD_7041_out0;
assign v$CINA_8864_out0 = v$COUTD_7041_out0;
assign v$CINA_8865_out0 = v$COUTD_7018_out0;
assign v$CINA_8876_out0 = v$COUTD_7041_out0;
assign v$CINA_8878_out0 = v$COUTD_7041_out0;
assign v$CINA_8885_out0 = v$COUTD_7041_out0;
assign v$CINA_8886_out0 = v$COUTD_7018_out0;
assign v$CINA_8978_out0 = v$COUTD_7164_out0;
assign v$CINA_8987_out0 = v$COUTD_7164_out0;
assign v$CINA_8988_out0 = v$COUTD_7141_out0;
assign v$CINA_8999_out0 = v$COUTD_7164_out0;
assign v$CINA_9001_out0 = v$COUTD_7164_out0;
assign v$CINA_9008_out0 = v$COUTD_7164_out0;
assign v$CINA_9009_out0 = v$COUTD_7141_out0;
assign v$G$AB_9562_out0 = v$G$AD_17769_out0;
assign v$G$AB_9569_out0 = v$G$AD_17769_out0;
assign v$G$AB_9573_out0 = v$G$AD_17790_out0;
assign v$G$AB_9576_out0 = v$G$AD_17790_out0;
assign v$G$AB_9584_out0 = v$G$AD_17769_out0;
assign v$G$AB_9685_out0 = v$G$AD_17892_out0;
assign v$G$AB_9692_out0 = v$G$AD_17892_out0;
assign v$G$AB_9696_out0 = v$G$AD_17913_out0;
assign v$G$AB_9699_out0 = v$G$AD_17913_out0;
assign v$G$AB_9707_out0 = v$G$AD_17892_out0;
assign v$C6_9968_out0 = v$COUTD_7022_out0;
assign v$C6_9971_out0 = v$COUTD_7145_out0;
assign v$P$CD_10947_out0 = v$P$AD_831_out0;
assign v$P$CD_10953_out0 = v$P$AD_793_out0;
assign v$P$CD_10961_out0 = v$P$AD_806_out0;
assign v$P$CD_10966_out0 = v$P$AD_812_out0;
assign v$P$CD_10970_out0 = v$P$AD_826_out0;
assign v$P$CD_10971_out0 = v$P$AD_792_out0;
assign v$P$CD_10979_out0 = v$P$AD_809_out0;
assign v$P$CD_11070_out0 = v$P$AD_954_out0;
assign v$P$CD_11076_out0 = v$P$AD_916_out0;
assign v$P$CD_11084_out0 = v$P$AD_929_out0;
assign v$P$CD_11089_out0 = v$P$AD_935_out0;
assign v$P$CD_11093_out0 = v$P$AD_949_out0;
assign v$P$CD_11094_out0 = v$P$AD_915_out0;
assign v$P$CD_11102_out0 = v$P$AD_932_out0;
assign v$C7_11477_out0 = v$COUTD_7051_out0;
assign v$C7_11480_out0 = v$COUTD_7174_out0;
assign v$G4_11652_out0 = v$G5_4731_out0 || v$G$CD_1059_out0;
assign v$G4_11653_out0 = v$G5_4732_out0 || v$G$CD_1060_out0;
assign v$G4_11666_out0 = v$G5_4745_out0 || v$G$CD_1073_out0;
assign v$G4_11668_out0 = v$G5_4747_out0 || v$G$CD_1075_out0;
assign v$G4_11669_out0 = v$G5_4748_out0 || v$G$CD_1076_out0;
assign v$G4_11672_out0 = v$G5_4751_out0 || v$G$CD_1079_out0;
assign v$G4_11686_out0 = v$G5_4765_out0 || v$G$CD_1093_out0;
assign v$G4_11691_out0 = v$G5_4770_out0 || v$G$CD_1098_out0;
assign v$G4_11775_out0 = v$G5_4854_out0 || v$G$CD_1182_out0;
assign v$G4_11776_out0 = v$G5_4855_out0 || v$G$CD_1183_out0;
assign v$G4_11789_out0 = v$G5_4868_out0 || v$G$CD_1196_out0;
assign v$G4_11791_out0 = v$G5_4870_out0 || v$G$CD_1198_out0;
assign v$G4_11792_out0 = v$G5_4871_out0 || v$G$CD_1199_out0;
assign v$G4_11795_out0 = v$G5_4874_out0 || v$G$CD_1202_out0;
assign v$G4_11809_out0 = v$G5_4888_out0 || v$G$CD_1216_out0;
assign v$G4_11814_out0 = v$G5_4893_out0 || v$G$CD_1221_out0;
assign v$G8_11967_out0 = v$CINA_8812_out0 && v$P$AB_2206_out0;
assign v$G8_11968_out0 = v$CINA_8813_out0 && v$P$AB_2207_out0;
assign v$G8_11981_out0 = v$CINA_8826_out0 && v$P$AB_2220_out0;
assign v$G8_11983_out0 = v$CINA_8828_out0 && v$P$AB_2222_out0;
assign v$G8_11984_out0 = v$CINA_8829_out0 && v$P$AB_2223_out0;
assign v$G8_11987_out0 = v$CINA_8832_out0 && v$P$AB_2226_out0;
assign v$G8_12001_out0 = v$CINA_8846_out0 && v$P$AB_2240_out0;
assign v$G8_12006_out0 = v$CINA_8851_out0 && v$P$AB_2245_out0;
assign v$G8_12090_out0 = v$CINA_8935_out0 && v$P$AB_2329_out0;
assign v$G8_12091_out0 = v$CINA_8936_out0 && v$P$AB_2330_out0;
assign v$G8_12104_out0 = v$CINA_8949_out0 && v$P$AB_2343_out0;
assign v$G8_12106_out0 = v$CINA_8951_out0 && v$P$AB_2345_out0;
assign v$G8_12107_out0 = v$CINA_8952_out0 && v$P$AB_2346_out0;
assign v$G8_12110_out0 = v$CINA_8955_out0 && v$P$AB_2349_out0;
assign v$G8_12124_out0 = v$CINA_8969_out0 && v$P$AB_2363_out0;
assign v$G8_12129_out0 = v$CINA_8974_out0 && v$P$AB_2368_out0;
assign v$C1_12422_out0 = v$C1_17402_out0;
assign v$C1_12425_out0 = v$C1_17405_out0;
assign {v$A3A_12526_out1,v$A3A_12526_out0 } = v$A2_18869_out0 + v$B2_3327_out0 + v$C1_17402_out0;
assign {v$A3A_12529_out1,v$A3A_12529_out0 } = v$A2_18872_out0 + v$B2_3330_out0 + v$C1_17405_out0;
assign v$END20_13849_out0 = v$G$AD_17779_out0;
assign v$END20_13852_out0 = v$G$AD_17902_out0;
assign v$END28_14250_out0 = v$G$AD_17790_out0;
assign v$END28_14253_out0 = v$G$AD_17913_out0;
assign v$C11_15406_out0 = v$COUTD_7041_out0;
assign v$C11_15409_out0 = v$COUTD_7164_out0;
assign v$END22_16075_out0 = v$G$AD_17800_out0;
assign v$END22_16078_out0 = v$G$AD_17923_out0;
assign v$END24_17024_out0 = v$G$AD_17778_out0;
assign v$END24_17027_out0 = v$G$AD_17901_out0;
assign v$END61_18572_out0 = v$COUTD_7049_out0;
assign v$END61_18575_out0 = v$COUTD_7172_out0;
assign {v$A8A_1661_out1,v$A8A_1661_out0 } = v$A7_15893_out0 + v$B7_17636_out0 + v$C6_9968_out0;
assign {v$A8A_1664_out1,v$A8A_1664_out0 } = v$A7_15896_out0 + v$B7_17639_out0 + v$C6_9971_out0;
assign {v$A17A_2684_out1,v$A17A_2684_out0 } = v$A12_3357_out0 + v$B12_2116_out0 + v$C11_15406_out0;
assign {v$A17A_2687_out1,v$A17A_2687_out0 } = v$A12_3360_out0 + v$B12_2119_out0 + v$C11_15409_out0;
assign v$G5_4787_out0 = v$G$AB_9562_out0 && v$P$CD_11004_out0;
assign v$G5_4794_out0 = v$G$AB_9569_out0 && v$P$CD_11011_out0;
assign v$G5_4798_out0 = v$G$AB_9573_out0 && v$P$CD_11015_out0;
assign v$G5_4801_out0 = v$G$AB_9576_out0 && v$P$CD_11018_out0;
assign v$G5_4809_out0 = v$G$AB_9584_out0 && v$P$CD_11026_out0;
assign v$G5_4910_out0 = v$G$AB_9685_out0 && v$P$CD_11127_out0;
assign v$G5_4917_out0 = v$G$AB_9692_out0 && v$P$CD_11134_out0;
assign v$G5_4921_out0 = v$G$AB_9696_out0 && v$P$CD_11138_out0;
assign v$G5_4924_out0 = v$G$AB_9699_out0 && v$P$CD_11141_out0;
assign v$G5_4932_out0 = v$G$AB_9707_out0 && v$P$CD_11149_out0;
assign v$END2_5450_out0 = v$A3A_12526_out1;
assign v$END2_5453_out0 = v$A3A_12529_out1;
assign v$G1_5804_out0 = v$P$AB_2205_out0 && v$P$CD_10947_out0;
assign v$G1_5809_out0 = v$P$AB_2210_out0 && v$P$CD_10952_out0;
assign v$G1_5815_out0 = v$P$AB_2216_out0 && v$P$CD_10958_out0;
assign v$G1_5818_out0 = v$P$AB_2219_out0 && v$P$CD_10961_out0;
assign v$G1_5823_out0 = v$P$AB_2224_out0 && v$P$CD_10966_out0;
assign v$G1_5836_out0 = v$P$AB_2237_out0 && v$P$CD_10979_out0;
assign v$G1_5927_out0 = v$P$AB_2328_out0 && v$P$CD_11070_out0;
assign v$G1_5932_out0 = v$P$AB_2333_out0 && v$P$CD_11075_out0;
assign v$G1_5938_out0 = v$P$AB_2339_out0 && v$P$CD_11081_out0;
assign v$G1_5941_out0 = v$P$AB_2342_out0 && v$P$CD_11084_out0;
assign v$G1_5946_out0 = v$P$AB_2347_out0 && v$P$CD_11089_out0;
assign v$G1_5959_out0 = v$P$AB_2360_out0 && v$P$CD_11102_out0;
assign v$C6_7343_out0 = v$C6_9968_out0;
assign v$C6_7346_out0 = v$C6_9971_out0;
assign v$_9236_out0 = { v$C0_9746_out0,v$C1_12422_out0 };
assign v$_9239_out0 = { v$C0_9749_out0,v$C1_12425_out0 };
assign v$C11_9889_out0 = v$C11_15406_out0;
assign v$C11_9892_out0 = v$C11_15409_out0;
assign v$G7_10059_out0 = v$G8_11967_out0 && v$P$CD_10948_out0;
assign v$G7_10060_out0 = v$G8_11968_out0 && v$P$CD_10949_out0;
assign v$G7_10073_out0 = v$G8_11981_out0 && v$P$CD_10962_out0;
assign v$G7_10075_out0 = v$G8_11983_out0 && v$P$CD_10964_out0;
assign v$G7_10076_out0 = v$G8_11984_out0 && v$P$CD_10965_out0;
assign v$G7_10079_out0 = v$G8_11987_out0 && v$P$CD_10968_out0;
assign v$G7_10093_out0 = v$G8_12001_out0 && v$P$CD_10982_out0;
assign v$G7_10098_out0 = v$G8_12006_out0 && v$P$CD_10987_out0;
assign v$G7_10182_out0 = v$G8_12090_out0 && v$P$CD_11071_out0;
assign v$G7_10183_out0 = v$G8_12091_out0 && v$P$CD_11072_out0;
assign v$G7_10196_out0 = v$G8_12104_out0 && v$P$CD_11085_out0;
assign v$G7_10198_out0 = v$G8_12106_out0 && v$P$CD_11087_out0;
assign v$G7_10199_out0 = v$G8_12107_out0 && v$P$CD_11088_out0;
assign v$G7_10202_out0 = v$G8_12110_out0 && v$P$CD_11091_out0;
assign v$G7_10216_out0 = v$G8_12124_out0 && v$P$CD_11105_out0;
assign v$G7_10221_out0 = v$G8_12129_out0 && v$P$CD_11110_out0;
assign {v$A9A_10864_out1,v$A9A_10864_out0 } = v$A8_18699_out0 + v$B8_13717_out0 + v$C7_11477_out0;
assign {v$A9A_10867_out1,v$A9A_10867_out0 } = v$A8_18702_out0 + v$B8_13720_out0 + v$C7_11480_out0;
assign v$G8_12010_out0 = v$CINA_8855_out0 && v$P$AB_2249_out0;
assign v$G8_12019_out0 = v$CINA_8864_out0 && v$P$AB_2258_out0;
assign v$G8_12020_out0 = v$CINA_8865_out0 && v$P$AB_2259_out0;
assign v$G8_12031_out0 = v$CINA_8876_out0 && v$P$AB_2270_out0;
assign v$G8_12033_out0 = v$CINA_8878_out0 && v$P$AB_2272_out0;
assign v$G8_12040_out0 = v$CINA_8885_out0 && v$P$AB_2279_out0;
assign v$G8_12041_out0 = v$CINA_8886_out0 && v$P$AB_2280_out0;
assign v$G8_12133_out0 = v$CINA_8978_out0 && v$P$AB_2372_out0;
assign v$G8_12142_out0 = v$CINA_8987_out0 && v$P$AB_2381_out0;
assign v$G8_12143_out0 = v$CINA_8988_out0 && v$P$AB_2382_out0;
assign v$G8_12154_out0 = v$CINA_8999_out0 && v$P$AB_2393_out0;
assign v$G8_12156_out0 = v$CINA_9001_out0 && v$P$AB_2395_out0;
assign v$G8_12163_out0 = v$CINA_9008_out0 && v$P$AB_2402_out0;
assign v$G8_12164_out0 = v$CINA_9009_out0 && v$P$AB_2403_out0;
assign v$END51_12244_out0 = v$P$AD_841_out0;
assign v$END51_12247_out0 = v$P$AD_964_out0;
assign {v$A10A_16614_out1,v$A10A_16614_out0 } = v$A9_3645_out0 + v$B9_4222_out0 + v$C8_7750_out0;
assign {v$A10A_16617_out1,v$A10A_16617_out0 } = v$A9_3648_out0 + v$B9_4225_out0 + v$C8_7753_out0;
assign v$C7_17053_out0 = v$C7_11477_out0;
assign v$C7_17056_out0 = v$C7_11480_out0;
assign v$G$AD_17726_out0 = v$G4_11652_out0;
assign v$G$AD_17727_out0 = v$G4_11653_out0;
assign v$G$AD_17740_out0 = v$G4_11666_out0;
assign v$G$AD_17742_out0 = v$G4_11668_out0;
assign v$G$AD_17743_out0 = v$G4_11669_out0;
assign v$G$AD_17746_out0 = v$G4_11672_out0;
assign v$G$AD_17760_out0 = v$G4_11686_out0;
assign v$G$AD_17765_out0 = v$G4_11691_out0;
assign v$G$AD_17849_out0 = v$G4_11775_out0;
assign v$G$AD_17850_out0 = v$G4_11776_out0;
assign v$G$AD_17863_out0 = v$G4_11789_out0;
assign v$G$AD_17865_out0 = v$G4_11791_out0;
assign v$G$AD_17866_out0 = v$G4_11792_out0;
assign v$G$AD_17869_out0 = v$G4_11795_out0;
assign v$G$AD_17883_out0 = v$G4_11809_out0;
assign v$G$AD_17888_out0 = v$G4_11814_out0;
assign v$END49_19061_out0 = v$P$AD_860_out0;
assign v$END49_19064_out0 = v$P$AD_983_out0;
assign v$C8_19109_out0 = v$C8_7750_out0;
assign v$C8_19112_out0 = v$C8_7753_out0;
assign v$G6_494_out0 = v$G4_11652_out0 || v$G7_10059_out0;
assign v$G6_495_out0 = v$G4_11653_out0 || v$G7_10060_out0;
assign v$G6_508_out0 = v$G4_11666_out0 || v$G7_10073_out0;
assign v$G6_510_out0 = v$G4_11668_out0 || v$G7_10075_out0;
assign v$G6_511_out0 = v$G4_11669_out0 || v$G7_10076_out0;
assign v$G6_514_out0 = v$G4_11672_out0 || v$G7_10079_out0;
assign v$G6_528_out0 = v$G4_11686_out0 || v$G7_10093_out0;
assign v$G6_533_out0 = v$G4_11691_out0 || v$G7_10098_out0;
assign v$G6_617_out0 = v$G4_11775_out0 || v$G7_10182_out0;
assign v$G6_618_out0 = v$G4_11776_out0 || v$G7_10183_out0;
assign v$G6_631_out0 = v$G4_11789_out0 || v$G7_10196_out0;
assign v$G6_633_out0 = v$G4_11791_out0 || v$G7_10198_out0;
assign v$G6_634_out0 = v$G4_11792_out0 || v$G7_10199_out0;
assign v$G6_637_out0 = v$G4_11795_out0 || v$G7_10202_out0;
assign v$G6_651_out0 = v$G4_11809_out0 || v$G7_10216_out0;
assign v$G6_656_out0 = v$G4_11814_out0 || v$G7_10221_out0;
assign v$P$AD_791_out0 = v$G1_5804_out0;
assign v$P$AD_796_out0 = v$G1_5809_out0;
assign v$P$AD_802_out0 = v$G1_5815_out0;
assign v$P$AD_805_out0 = v$G1_5818_out0;
assign v$P$AD_810_out0 = v$G1_5823_out0;
assign v$P$AD_823_out0 = v$G1_5836_out0;
assign v$P$AD_914_out0 = v$G1_5927_out0;
assign v$P$AD_919_out0 = v$G1_5932_out0;
assign v$P$AD_925_out0 = v$G1_5938_out0;
assign v$P$AD_928_out0 = v$G1_5941_out0;
assign v$P$AD_933_out0 = v$G1_5946_out0;
assign v$P$AD_946_out0 = v$G1_5959_out0;
assign v$G$CD_1058_out0 = v$G$AD_17765_out0;
assign v$G$CD_1064_out0 = v$G$AD_17727_out0;
assign v$G$CD_1072_out0 = v$G$AD_17740_out0;
assign v$G$CD_1077_out0 = v$G$AD_17746_out0;
assign v$G$CD_1081_out0 = v$G$AD_17760_out0;
assign v$G$CD_1082_out0 = v$G$AD_17726_out0;
assign v$G$CD_1090_out0 = v$G$AD_17743_out0;
assign v$G$CD_1181_out0 = v$G$AD_17888_out0;
assign v$G$CD_1187_out0 = v$G$AD_17850_out0;
assign v$G$CD_1195_out0 = v$G$AD_17863_out0;
assign v$G$CD_1200_out0 = v$G$AD_17869_out0;
assign v$G$CD_1204_out0 = v$G$AD_17883_out0;
assign v$G$CD_1205_out0 = v$G$AD_17849_out0;
assign v$G$CD_1213_out0 = v$G$AD_17866_out0;
assign v$END7_3584_out0 = v$A8A_1661_out1;
assign v$END7_3587_out0 = v$A8A_1664_out1;
assign v$_3828_out0 = { v$A6A_3336_out0,v$A8A_1661_out0 };
assign v$_3831_out0 = { v$A6A_3339_out0,v$A8A_1664_out0 };
assign v$END8_4072_out0 = v$A9A_10864_out1;
assign v$END8_4075_out0 = v$A9A_10867_out1;
assign v$END9_4394_out0 = v$A10A_16614_out1;
assign v$END9_4397_out0 = v$A10A_16617_out1;
assign v$G$AB_9505_out0 = v$G$AD_17727_out0;
assign v$G$AB_9510_out0 = v$G$AD_17742_out0;
assign v$G$AB_9516_out0 = v$G$AD_17742_out0;
assign v$G$AB_9519_out0 = v$G$AD_17760_out0;
assign v$G$AB_9524_out0 = v$G$AD_17726_out0;
assign v$G$AB_9537_out0 = v$G$AD_17742_out0;
assign v$G$AB_9628_out0 = v$G$AD_17850_out0;
assign v$G$AB_9633_out0 = v$G$AD_17865_out0;
assign v$G$AB_9639_out0 = v$G$AD_17865_out0;
assign v$G$AB_9642_out0 = v$G$AD_17883_out0;
assign v$G$AB_9647_out0 = v$G$AD_17849_out0;
assign v$G$AB_9660_out0 = v$G$AD_17865_out0;
assign v$ENDw_9932_out0 = v$A17A_2684_out1;
assign v$ENDw_9935_out0 = v$A17A_2687_out1;
assign v$G7_10102_out0 = v$G8_12010_out0 && v$P$CD_10991_out0;
assign v$G7_10111_out0 = v$G8_12019_out0 && v$P$CD_11000_out0;
assign v$G7_10112_out0 = v$G8_12020_out0 && v$P$CD_11001_out0;
assign v$G7_10123_out0 = v$G8_12031_out0 && v$P$CD_11012_out0;
assign v$G7_10125_out0 = v$G8_12033_out0 && v$P$CD_11014_out0;
assign v$G7_10132_out0 = v$G8_12040_out0 && v$P$CD_11021_out0;
assign v$G7_10133_out0 = v$G8_12041_out0 && v$P$CD_11022_out0;
assign v$G7_10225_out0 = v$G8_12133_out0 && v$P$CD_11114_out0;
assign v$G7_10234_out0 = v$G8_12142_out0 && v$P$CD_11123_out0;
assign v$G7_10235_out0 = v$G8_12143_out0 && v$P$CD_11124_out0;
assign v$G7_10246_out0 = v$G8_12154_out0 && v$P$CD_11135_out0;
assign v$G7_10248_out0 = v$G8_12156_out0 && v$P$CD_11137_out0;
assign v$G7_10255_out0 = v$G8_12163_out0 && v$P$CD_11144_out0;
assign v$G7_10256_out0 = v$G8_12164_out0 && v$P$CD_11145_out0;
assign v$G4_11708_out0 = v$G5_4787_out0 || v$G$CD_1115_out0;
assign v$G4_11715_out0 = v$G5_4794_out0 || v$G$CD_1122_out0;
assign v$G4_11719_out0 = v$G5_4798_out0 || v$G$CD_1126_out0;
assign v$G4_11722_out0 = v$G5_4801_out0 || v$G$CD_1129_out0;
assign v$G4_11730_out0 = v$G5_4809_out0 || v$G$CD_1137_out0;
assign v$G4_11831_out0 = v$G5_4910_out0 || v$G$CD_1238_out0;
assign v$G4_11838_out0 = v$G5_4917_out0 || v$G$CD_1245_out0;
assign v$G4_11842_out0 = v$G5_4921_out0 || v$G$CD_1249_out0;
assign v$G4_11845_out0 = v$G5_4924_out0 || v$G$CD_1252_out0;
assign v$G4_11853_out0 = v$G5_4932_out0 || v$G$CD_1260_out0;
assign v$_15632_out0 = { v$A9A_10864_out0,v$A10A_16614_out0 };
assign v$_15635_out0 = { v$A9A_10867_out0,v$A10A_16617_out0 };
assign v$_16926_out0 = { v$C6_7343_out0,v$C7_17053_out0 };
assign v$_16929_out0 = { v$C6_7346_out0,v$C7_17056_out0 };
assign v$G6_537_out0 = v$G4_11695_out0 || v$G7_10102_out0;
assign v$G6_546_out0 = v$G4_11704_out0 || v$G7_10111_out0;
assign v$G6_547_out0 = v$G4_11705_out0 || v$G7_10112_out0;
assign v$G6_558_out0 = v$G4_11716_out0 || v$G7_10123_out0;
assign v$G6_560_out0 = v$G4_11718_out0 || v$G7_10125_out0;
assign v$G6_567_out0 = v$G4_11725_out0 || v$G7_10132_out0;
assign v$G6_568_out0 = v$G4_11726_out0 || v$G7_10133_out0;
assign v$G6_660_out0 = v$G4_11818_out0 || v$G7_10225_out0;
assign v$G6_669_out0 = v$G4_11827_out0 || v$G7_10234_out0;
assign v$G6_670_out0 = v$G4_11828_out0 || v$G7_10235_out0;
assign v$G6_681_out0 = v$G4_11839_out0 || v$G7_10246_out0;
assign v$G6_683_out0 = v$G4_11841_out0 || v$G7_10248_out0;
assign v$G6_690_out0 = v$G4_11848_out0 || v$G7_10255_out0;
assign v$G6_691_out0 = v$G4_11849_out0 || v$G7_10256_out0;
assign v$P$AB_2211_out0 = v$P$AD_823_out0;
assign v$P$AB_2215_out0 = v$P$AD_823_out0;
assign v$P$AB_2234_out0 = v$P$AD_823_out0;
assign v$P$AB_2242_out0 = v$P$AD_810_out0;
assign v$P$AB_2244_out0 = v$P$AD_823_out0;
assign v$P$AB_2334_out0 = v$P$AD_946_out0;
assign v$P$AB_2338_out0 = v$P$AD_946_out0;
assign v$P$AB_2357_out0 = v$P$AD_946_out0;
assign v$P$AB_2365_out0 = v$P$AD_933_out0;
assign v$P$AB_2367_out0 = v$P$AD_946_out0;
assign v$G5_4730_out0 = v$G$AB_9505_out0 && v$P$CD_10947_out0;
assign v$G5_4735_out0 = v$G$AB_9510_out0 && v$P$CD_10952_out0;
assign v$G5_4741_out0 = v$G$AB_9516_out0 && v$P$CD_10958_out0;
assign v$G5_4744_out0 = v$G$AB_9519_out0 && v$P$CD_10961_out0;
assign v$G5_4749_out0 = v$G$AB_9524_out0 && v$P$CD_10966_out0;
assign v$G5_4762_out0 = v$G$AB_9537_out0 && v$P$CD_10979_out0;
assign v$G5_4853_out0 = v$G$AB_9628_out0 && v$P$CD_11070_out0;
assign v$G5_4858_out0 = v$G$AB_9633_out0 && v$P$CD_11075_out0;
assign v$G5_4864_out0 = v$G$AB_9639_out0 && v$P$CD_11081_out0;
assign v$G5_4867_out0 = v$G$AB_9642_out0 && v$P$CD_11084_out0;
assign v$G5_4872_out0 = v$G$AB_9647_out0 && v$P$CD_11089_out0;
assign v$G5_4885_out0 = v$G$AB_9660_out0 && v$P$CD_11102_out0;
assign v$COUTD_6972_out0 = v$G6_494_out0;
assign v$COUTD_6973_out0 = v$G6_495_out0;
assign v$COUTD_6986_out0 = v$G6_508_out0;
assign v$COUTD_6988_out0 = v$G6_510_out0;
assign v$COUTD_6989_out0 = v$G6_511_out0;
assign v$COUTD_6992_out0 = v$G6_514_out0;
assign v$COUTD_7006_out0 = v$G6_528_out0;
assign v$COUTD_7011_out0 = v$G6_533_out0;
assign v$COUTD_7095_out0 = v$G6_617_out0;
assign v$COUTD_7096_out0 = v$G6_618_out0;
assign v$COUTD_7109_out0 = v$G6_631_out0;
assign v$COUTD_7111_out0 = v$G6_633_out0;
assign v$COUTD_7112_out0 = v$G6_634_out0;
assign v$COUTD_7115_out0 = v$G6_637_out0;
assign v$COUTD_7129_out0 = v$G6_651_out0;
assign v$COUTD_7134_out0 = v$G6_656_out0;
assign v$_7721_out0 = { v$_2648_out0,v$_16926_out0 };
assign v$_7724_out0 = { v$_2651_out0,v$_16929_out0 };
assign v$P$CD_10950_out0 = v$P$AD_810_out0;
assign v$P$CD_10976_out0 = v$P$AD_791_out0;
assign v$P$CD_10984_out0 = v$P$AD_805_out0;
assign v$P$CD_11073_out0 = v$P$AD_933_out0;
assign v$P$CD_11099_out0 = v$P$AD_914_out0;
assign v$P$CD_11107_out0 = v$P$AD_928_out0;
assign v$END11_12656_out0 = v$P$AD_802_out0;
assign v$END11_12659_out0 = v$P$AD_925_out0;
assign v$G$AD_17782_out0 = v$G4_11708_out0;
assign v$G$AD_17789_out0 = v$G4_11715_out0;
assign v$G$AD_17793_out0 = v$G4_11719_out0;
assign v$G$AD_17796_out0 = v$G4_11722_out0;
assign v$G$AD_17804_out0 = v$G4_11730_out0;
assign v$G$AD_17905_out0 = v$G4_11831_out0;
assign v$G$AD_17912_out0 = v$G4_11838_out0;
assign v$G$AD_17916_out0 = v$G4_11842_out0;
assign v$G$AD_17919_out0 = v$G4_11845_out0;
assign v$G$AD_17927_out0 = v$G4_11853_out0;
assign v$_18581_out0 = { v$_84_out0,v$_3828_out0 };
assign v$_18584_out0 = { v$_87_out0,v$_3831_out0 };
assign v$END13_18674_out0 = v$P$AD_796_out0;
assign v$END13_18677_out0 = v$P$AD_919_out0;
assign v$END1_1451_out0 = v$COUTD_7011_out0;
assign v$END1_1454_out0 = v$COUTD_7134_out0;
assign v$END32_2666_out0 = v$G$AD_17796_out0;
assign v$END32_2669_out0 = v$G$AD_17919_out0;
assign v$C2_2885_out0 = v$COUTD_6988_out0;
assign v$C2_2888_out0 = v$COUTD_7111_out0;
assign v$END_3542_out0 = v$COUTD_6989_out0;
assign v$END_3545_out0 = v$COUTD_7112_out0;
assign v$END3_3656_out0 = v$COUTD_6986_out0;
assign v$END3_3659_out0 = v$COUTD_7109_out0;
assign v$G1_5810_out0 = v$P$AB_2211_out0 && v$P$CD_10953_out0;
assign v$G1_5814_out0 = v$P$AB_2215_out0 && v$P$CD_10957_out0;
assign v$G1_5833_out0 = v$P$AB_2234_out0 && v$P$CD_10976_out0;
assign v$G1_5841_out0 = v$P$AB_2242_out0 && v$P$CD_10984_out0;
assign v$G1_5843_out0 = v$P$AB_2244_out0 && v$P$CD_10986_out0;
assign v$G1_5933_out0 = v$P$AB_2334_out0 && v$P$CD_11076_out0;
assign v$G1_5937_out0 = v$P$AB_2338_out0 && v$P$CD_11080_out0;
assign v$G1_5956_out0 = v$P$AB_2357_out0 && v$P$CD_11099_out0;
assign v$G1_5964_out0 = v$P$AB_2365_out0 && v$P$CD_11107_out0;
assign v$G1_5966_out0 = v$P$AB_2367_out0 && v$P$CD_11109_out0;
assign v$COUTD_7015_out0 = v$G6_537_out0;
assign v$COUTD_7024_out0 = v$G6_546_out0;
assign v$COUTD_7025_out0 = v$G6_547_out0;
assign v$COUTD_7036_out0 = v$G6_558_out0;
assign v$COUTD_7038_out0 = v$G6_560_out0;
assign v$COUTD_7045_out0 = v$G6_567_out0;
assign v$COUTD_7046_out0 = v$G6_568_out0;
assign v$COUTD_7138_out0 = v$G6_660_out0;
assign v$COUTD_7147_out0 = v$G6_669_out0;
assign v$COUTD_7148_out0 = v$G6_670_out0;
assign v$COUTD_7159_out0 = v$G6_681_out0;
assign v$COUTD_7161_out0 = v$G6_683_out0;
assign v$COUTD_7168_out0 = v$G6_690_out0;
assign v$COUTD_7169_out0 = v$G6_691_out0;
assign v$END2_8069_out0 = v$COUTD_6992_out0;
assign v$END2_8072_out0 = v$COUTD_7115_out0;
assign v$_8114_out0 = { v$_7570_out0,v$_7721_out0 };
assign v$_8117_out0 = { v$_7573_out0,v$_7724_out0 };
assign v$CINA_8811_out0 = v$COUTD_6973_out0;
assign v$CINA_8816_out0 = v$COUTD_6988_out0;
assign v$CINA_8822_out0 = v$COUTD_6988_out0;
assign v$CINA_8825_out0 = v$COUTD_7006_out0;
assign v$CINA_8830_out0 = v$COUTD_6972_out0;
assign v$CINA_8843_out0 = v$COUTD_6988_out0;
assign v$CINA_8934_out0 = v$COUTD_7096_out0;
assign v$CINA_8939_out0 = v$COUTD_7111_out0;
assign v$CINA_8945_out0 = v$COUTD_7111_out0;
assign v$CINA_8948_out0 = v$COUTD_7129_out0;
assign v$CINA_8953_out0 = v$COUTD_7095_out0;
assign v$CINA_8966_out0 = v$COUTD_7111_out0;
assign v$END45_9384_out0 = v$COUTD_7006_out0;
assign v$END45_9387_out0 = v$COUTD_7129_out0;
assign v$G$AB_9555_out0 = v$G$AD_17789_out0;
assign v$G$AB_9574_out0 = v$G$AD_17789_out0;
assign v$G$AB_9678_out0 = v$G$AD_17912_out0;
assign v$G$AB_9697_out0 = v$G$AD_17912_out0;
assign v$G4_11651_out0 = v$G5_4730_out0 || v$G$CD_1058_out0;
assign v$G4_11656_out0 = v$G5_4735_out0 || v$G$CD_1063_out0;
assign v$G4_11662_out0 = v$G5_4741_out0 || v$G$CD_1069_out0;
assign v$G4_11665_out0 = v$G5_4744_out0 || v$G$CD_1072_out0;
assign v$G4_11670_out0 = v$G5_4749_out0 || v$G$CD_1077_out0;
assign v$G4_11683_out0 = v$G5_4762_out0 || v$G$CD_1090_out0;
assign v$G4_11774_out0 = v$G5_4853_out0 || v$G$CD_1181_out0;
assign v$G4_11779_out0 = v$G5_4858_out0 || v$G$CD_1186_out0;
assign v$G4_11785_out0 = v$G5_4864_out0 || v$G$CD_1192_out0;
assign v$G4_11788_out0 = v$G5_4867_out0 || v$G$CD_1195_out0;
assign v$G4_11793_out0 = v$G5_4872_out0 || v$G$CD_1200_out0;
assign v$G4_11806_out0 = v$G5_4885_out0 || v$G$CD_1213_out0;
assign v$END43_13773_out0 = v$G$AD_17804_out0;
assign v$END43_13776_out0 = v$G$AD_17927_out0;
assign v$END46_15665_out0 = v$G$AD_17789_out0;
assign v$END46_15668_out0 = v$G$AD_17912_out0;
assign v$END30_16311_out0 = v$G$AD_17793_out0;
assign v$END30_16314_out0 = v$G$AD_17916_out0;
assign v$END41_17288_out0 = v$G$AD_17782_out0;
assign v$END41_17291_out0 = v$G$AD_17905_out0;
assign v$_18360_out0 = { v$_10819_out0,v$_18581_out0 };
assign v$_18363_out0 = { v$_10822_out0,v$_18584_out0 };
assign v$C14_292_out0 = v$COUTD_7036_out0;
assign v$C14_295_out0 = v$COUTD_7159_out0;
assign v$P$AD_797_out0 = v$G1_5810_out0;
assign v$P$AD_801_out0 = v$G1_5814_out0;
assign v$P$AD_820_out0 = v$G1_5833_out0;
assign v$P$AD_828_out0 = v$G1_5841_out0;
assign v$P$AD_830_out0 = v$G1_5843_out0;
assign v$P$AD_920_out0 = v$G1_5933_out0;
assign v$P$AD_924_out0 = v$G1_5937_out0;
assign v$P$AD_943_out0 = v$G1_5956_out0;
assign v$P$AD_951_out0 = v$G1_5964_out0;
assign v$P$AD_953_out0 = v$G1_5966_out0;
assign v$C17_2718_out0 = v$COUTD_7015_out0;
assign v$C17_2721_out0 = v$COUTD_7138_out0;
assign v$G5_4780_out0 = v$G$AB_9555_out0 && v$P$CD_10997_out0;
assign v$G5_4799_out0 = v$G$AB_9574_out0 && v$P$CD_11016_out0;
assign v$G5_4903_out0 = v$G$AB_9678_out0 && v$P$CD_11120_out0;
assign v$G5_4922_out0 = v$G$AB_9697_out0 && v$P$CD_11139_out0;
assign v$C23_5058_out0 = v$COUTD_7038_out0;
assign v$C23_5061_out0 = v$COUTD_7161_out0;
assign v$C9_6218_out0 = v$COUTD_7025_out0;
assign v$C9_6221_out0 = v$COUTD_7148_out0;
assign v$CINA_8868_out0 = v$COUTD_7015_out0;
assign v$CINA_8875_out0 = v$COUTD_7015_out0;
assign v$CINA_8879_out0 = v$COUTD_7036_out0;
assign v$CINA_8882_out0 = v$COUTD_7036_out0;
assign v$CINA_8890_out0 = v$COUTD_7015_out0;
assign v$CINA_8991_out0 = v$COUTD_7138_out0;
assign v$CINA_8998_out0 = v$COUTD_7138_out0;
assign v$CINA_9002_out0 = v$COUTD_7159_out0;
assign v$CINA_9005_out0 = v$COUTD_7159_out0;
assign v$CINA_9013_out0 = v$COUTD_7138_out0;
assign v$G8_11966_out0 = v$CINA_8811_out0 && v$P$AB_2205_out0;
assign v$G8_11971_out0 = v$CINA_8816_out0 && v$P$AB_2210_out0;
assign v$G8_11977_out0 = v$CINA_8822_out0 && v$P$AB_2216_out0;
assign v$G8_11980_out0 = v$CINA_8825_out0 && v$P$AB_2219_out0;
assign v$G8_11985_out0 = v$CINA_8830_out0 && v$P$AB_2224_out0;
assign v$G8_11998_out0 = v$CINA_8843_out0 && v$P$AB_2237_out0;
assign v$G8_12089_out0 = v$CINA_8934_out0 && v$P$AB_2328_out0;
assign v$G8_12094_out0 = v$CINA_8939_out0 && v$P$AB_2333_out0;
assign v$G8_12100_out0 = v$CINA_8945_out0 && v$P$AB_2339_out0;
assign v$G8_12103_out0 = v$CINA_8948_out0 && v$P$AB_2342_out0;
assign v$G8_12108_out0 = v$CINA_8953_out0 && v$P$AB_2347_out0;
assign v$G8_12121_out0 = v$CINA_8966_out0 && v$P$AB_2360_out0;
assign v$C13_12348_out0 = v$COUTD_7045_out0;
assign v$C13_12351_out0 = v$COUTD_7168_out0;
assign v$C10_13303_out0 = v$COUTD_7046_out0;
assign v$C10_13306_out0 = v$COUTD_7169_out0;
assign {v$A4A_13732_out1,v$A4A_13732_out0 } = v$A3_15210_out0 + v$B3_9846_out0 + v$C2_2885_out0;
assign {v$A4A_13735_out1,v$A4A_13735_out0 } = v$A3_15213_out0 + v$B3_9849_out0 + v$C2_2888_out0;
assign v$C12_14096_out0 = v$COUTD_7024_out0;
assign v$C12_14099_out0 = v$COUTD_7147_out0;
assign v$G$AD_17725_out0 = v$G4_11651_out0;
assign v$G$AD_17730_out0 = v$G4_11656_out0;
assign v$G$AD_17736_out0 = v$G4_11662_out0;
assign v$G$AD_17739_out0 = v$G4_11665_out0;
assign v$G$AD_17744_out0 = v$G4_11670_out0;
assign v$G$AD_17757_out0 = v$G4_11683_out0;
assign v$G$AD_17848_out0 = v$G4_11774_out0;
assign v$G$AD_17853_out0 = v$G4_11779_out0;
assign v$G$AD_17859_out0 = v$G4_11785_out0;
assign v$G$AD_17862_out0 = v$G4_11788_out0;
assign v$G$AD_17867_out0 = v$G4_11793_out0;
assign v$G$AD_17880_out0 = v$G4_11806_out0;
assign v$C2_18778_out0 = v$C2_2885_out0;
assign v$C2_18781_out0 = v$C2_2888_out0;
assign v$C14_342_out0 = v$C14_292_out0;
assign v$C14_345_out0 = v$C14_295_out0;
assign v$G$CD_1061_out0 = v$G$AD_17744_out0;
assign v$G$CD_1087_out0 = v$G$AD_17725_out0;
assign v$G$CD_1095_out0 = v$G$AD_17739_out0;
assign v$G$CD_1184_out0 = v$G$AD_17867_out0;
assign v$G$CD_1210_out0 = v$G$AD_17848_out0;
assign v$G$CD_1218_out0 = v$G$AD_17862_out0;
assign v$END10_1296_out0 = v$G$AD_17736_out0;
assign v$END10_1299_out0 = v$G$AD_17859_out0;
assign v$C10_2105_out0 = v$C10_13303_out0;
assign v$C10_2108_out0 = v$C10_13306_out0;
assign v$P$AB_2208_out0 = v$P$AD_820_out0;
assign v$P$AB_2217_out0 = v$P$AD_820_out0;
assign v$P$AB_2218_out0 = v$P$AD_797_out0;
assign v$P$AB_2229_out0 = v$P$AD_820_out0;
assign v$P$AB_2231_out0 = v$P$AD_820_out0;
assign v$P$AB_2238_out0 = v$P$AD_820_out0;
assign v$P$AB_2239_out0 = v$P$AD_797_out0;
assign v$P$AB_2331_out0 = v$P$AD_943_out0;
assign v$P$AB_2340_out0 = v$P$AD_943_out0;
assign v$P$AB_2341_out0 = v$P$AD_920_out0;
assign v$P$AB_2352_out0 = v$P$AD_943_out0;
assign v$P$AB_2354_out0 = v$P$AD_943_out0;
assign v$P$AB_2361_out0 = v$P$AD_943_out0;
assign v$P$AB_2362_out0 = v$P$AD_920_out0;
assign {v$A12A_4615_out1,v$A12A_4615_out0 } = v$A11_10388_out0 + v$B11_9445_out0 + v$C10_13303_out0;
assign {v$A12A_4618_out1,v$A12A_4618_out0 } = v$A11_10391_out0 + v$B11_9448_out0 + v$C10_13306_out0;
assign v$C17_6344_out0 = v$C17_2718_out0;
assign v$C17_6347_out0 = v$C17_2721_out0;
assign {v$A13_7556_out1,v$A13_7556_out0 } = v$A15_17959_out0 + v$B15_10448_out0 + v$C14_292_out0;
assign {v$A13_7559_out1,v$A13_7559_out0 } = v$A15_17962_out0 + v$B15_10451_out0 + v$C14_295_out0;
assign v$END15_7697_out0 = v$P$AD_801_out0;
assign v$END15_7700_out0 = v$P$AD_924_out0;
assign v$END17_7966_out0 = v$P$AD_830_out0;
assign v$END17_7969_out0 = v$P$AD_953_out0;
assign v$END3_8258_out0 = v$A4A_13732_out1;
assign v$END3_8261_out0 = v$A4A_13735_out1;
assign v$G$AB_9511_out0 = v$G$AD_17757_out0;
assign v$G$AB_9515_out0 = v$G$AD_17757_out0;
assign v$G$AB_9534_out0 = v$G$AD_17757_out0;
assign v$G$AB_9542_out0 = v$G$AD_17744_out0;
assign v$G$AB_9544_out0 = v$G$AD_17757_out0;
assign v$G$AB_9634_out0 = v$G$AD_17880_out0;
assign v$G$AB_9638_out0 = v$G$AD_17880_out0;
assign v$G$AB_9657_out0 = v$G$AD_17880_out0;
assign v$G$AB_9665_out0 = v$G$AD_17867_out0;
assign v$G$AB_9667_out0 = v$G$AD_17880_out0;
assign v$C12_9769_out0 = v$C12_14096_out0;
assign v$C12_9772_out0 = v$C12_14099_out0;
assign v$G7_10058_out0 = v$G8_11966_out0 && v$P$CD_10947_out0;
assign v$G7_10063_out0 = v$G8_11971_out0 && v$P$CD_10952_out0;
assign v$G7_10069_out0 = v$G8_11977_out0 && v$P$CD_10958_out0;
assign v$G7_10072_out0 = v$G8_11980_out0 && v$P$CD_10961_out0;
assign v$G7_10077_out0 = v$G8_11985_out0 && v$P$CD_10966_out0;
assign v$G7_10090_out0 = v$G8_11998_out0 && v$P$CD_10979_out0;
assign v$G7_10181_out0 = v$G8_12089_out0 && v$P$CD_11070_out0;
assign v$G7_10186_out0 = v$G8_12094_out0 && v$P$CD_11075_out0;
assign v$G7_10192_out0 = v$G8_12100_out0 && v$P$CD_11081_out0;
assign v$G7_10195_out0 = v$G8_12103_out0 && v$P$CD_11084_out0;
assign v$G7_10200_out0 = v$G8_12108_out0 && v$P$CD_11089_out0;
assign v$G7_10213_out0 = v$G8_12121_out0 && v$P$CD_11102_out0;
assign {v$A18_10460_out1,v$A18_10460_out0 } = v$A13_14447_out0 + v$B13_9024_out0 + v$C12_14096_out0;
assign {v$A18_10463_out1,v$A18_10463_out0 } = v$A13_14450_out0 + v$B13_9027_out0 + v$C12_14099_out0;
assign v$P$CD_10973_out0 = v$P$AD_828_out0;
assign v$P$CD_11096_out0 = v$P$AD_951_out0;
assign v$END12_11275_out0 = v$G$AD_17730_out0;
assign v$END12_11278_out0 = v$G$AD_17853_out0;
assign v$G4_11701_out0 = v$G5_4780_out0 || v$G$CD_1108_out0;
assign v$G4_11720_out0 = v$G5_4799_out0 || v$G$CD_1127_out0;
assign v$G4_11824_out0 = v$G5_4903_out0 || v$G$CD_1231_out0;
assign v$G4_11843_out0 = v$G5_4922_out0 || v$G$CD_1250_out0;
assign v$G8_12023_out0 = v$CINA_8868_out0 && v$P$AB_2262_out0;
assign v$G8_12030_out0 = v$CINA_8875_out0 && v$P$AB_2269_out0;
assign v$G8_12034_out0 = v$CINA_8879_out0 && v$P$AB_2273_out0;
assign v$G8_12037_out0 = v$CINA_8882_out0 && v$P$AB_2276_out0;
assign v$G8_12045_out0 = v$CINA_8890_out0 && v$P$AB_2284_out0;
assign v$G8_12146_out0 = v$CINA_8991_out0 && v$P$AB_2385_out0;
assign v$G8_12153_out0 = v$CINA_8998_out0 && v$P$AB_2392_out0;
assign v$G8_12157_out0 = v$CINA_9002_out0 && v$P$AB_2396_out0;
assign v$G8_12160_out0 = v$CINA_9005_out0 && v$P$AB_2399_out0;
assign v$G8_12168_out0 = v$CINA_9013_out0 && v$P$AB_2407_out0;
assign v$END19_12219_out0 = v$P$AD_797_out0;
assign v$END19_12222_out0 = v$P$AD_920_out0;
assign v$C9_12718_out0 = v$C9_6218_out0;
assign v$C9_12721_out0 = v$C9_6221_out0;
assign {v$A15_13799_out1,v$A15_13799_out0 } = v$A18_18302_out0 + v$B18_11370_out0 + v$C17_2718_out0;
assign {v$A15_13802_out1,v$A15_13802_out0 } = v$A18_18305_out0 + v$B18_11373_out0 + v$C17_2721_out0;
assign {v$A16A_15160_out1,v$A16A_15160_out0 } = v$A10_1705_out0 + v$B10_10299_out0 + v$C9_6218_out0;
assign {v$A16A_15163_out1,v$A16A_15163_out0 } = v$A10_1708_out0 + v$B10_10302_out0 + v$C9_6221_out0;
assign v$C23_16760_out0 = v$C23_5058_out0;
assign v$C23_16763_out0 = v$C23_5061_out0;
assign {v$A20_16994_out1,v$A20_16994_out0 } = v$A14_740_out0 + v$B14_4160_out0 + v$C13_12348_out0;
assign {v$A20_16997_out1,v$A20_16997_out0 } = v$A14_743_out0 + v$B14_4163_out0 + v$C13_12351_out0;
assign v$C13_19199_out0 = v$C13_12348_out0;
assign v$C13_19202_out0 = v$C13_12351_out0;
assign v$_19275_out0 = { v$A3A_12526_out0,v$A4A_13732_out0 };
assign v$_19278_out0 = { v$A3A_12529_out0,v$A4A_13735_out0 };
assign v$G6_493_out0 = v$G4_11651_out0 || v$G7_10058_out0;
assign v$G6_498_out0 = v$G4_11656_out0 || v$G7_10063_out0;
assign v$G6_504_out0 = v$G4_11662_out0 || v$G7_10069_out0;
assign v$G6_507_out0 = v$G4_11665_out0 || v$G7_10072_out0;
assign v$G6_512_out0 = v$G4_11670_out0 || v$G7_10077_out0;
assign v$G6_525_out0 = v$G4_11683_out0 || v$G7_10090_out0;
assign v$G6_616_out0 = v$G4_11774_out0 || v$G7_10181_out0;
assign v$G6_621_out0 = v$G4_11779_out0 || v$G7_10186_out0;
assign v$G6_627_out0 = v$G4_11785_out0 || v$G7_10192_out0;
assign v$G6_630_out0 = v$G4_11788_out0 || v$G7_10195_out0;
assign v$G6_635_out0 = v$G4_11793_out0 || v$G7_10200_out0;
assign v$G6_648_out0 = v$G4_11806_out0 || v$G7_10213_out0;
assign v$ENDq_1611_out0 = v$A12A_4615_out1;
assign v$ENDq_1614_out0 = v$A12A_4618_out1;
assign v$G5_4736_out0 = v$G$AB_9511_out0 && v$P$CD_10953_out0;
assign v$G5_4740_out0 = v$G$AB_9515_out0 && v$P$CD_10957_out0;
assign v$G5_4759_out0 = v$G$AB_9534_out0 && v$P$CD_10976_out0;
assign v$G5_4767_out0 = v$G$AB_9542_out0 && v$P$CD_10984_out0;
assign v$G5_4769_out0 = v$G$AB_9544_out0 && v$P$CD_10986_out0;
assign v$G5_4859_out0 = v$G$AB_9634_out0 && v$P$CD_11076_out0;
assign v$G5_4863_out0 = v$G$AB_9638_out0 && v$P$CD_11080_out0;
assign v$G5_4882_out0 = v$G$AB_9657_out0 && v$P$CD_11099_out0;
assign v$G5_4890_out0 = v$G$AB_9665_out0 && v$P$CD_11107_out0;
assign v$G5_4892_out0 = v$G$AB_9667_out0 && v$P$CD_11109_out0;
assign v$G1_5807_out0 = v$P$AB_2208_out0 && v$P$CD_10950_out0;
assign v$G1_5816_out0 = v$P$AB_2217_out0 && v$P$CD_10959_out0;
assign v$G1_5817_out0 = v$P$AB_2218_out0 && v$P$CD_10960_out0;
assign v$G1_5828_out0 = v$P$AB_2229_out0 && v$P$CD_10971_out0;
assign v$G1_5830_out0 = v$P$AB_2231_out0 && v$P$CD_10973_out0;
assign v$G1_5837_out0 = v$P$AB_2238_out0 && v$P$CD_10980_out0;
assign v$G1_5838_out0 = v$P$AB_2239_out0 && v$P$CD_10981_out0;
assign v$G1_5930_out0 = v$P$AB_2331_out0 && v$P$CD_11073_out0;
assign v$G1_5939_out0 = v$P$AB_2340_out0 && v$P$CD_11082_out0;
assign v$G1_5940_out0 = v$P$AB_2341_out0 && v$P$CD_11083_out0;
assign v$G1_5951_out0 = v$P$AB_2352_out0 && v$P$CD_11094_out0;
assign v$G1_5953_out0 = v$P$AB_2354_out0 && v$P$CD_11096_out0;
assign v$G1_5960_out0 = v$P$AB_2361_out0 && v$P$CD_11103_out0;
assign v$G1_5961_out0 = v$P$AB_2362_out0 && v$P$CD_11104_out0;
assign v$_6175_out0 = { v$A17A_2684_out0,v$A18_10460_out0 };
assign v$_6178_out0 = { v$A17A_2687_out0,v$A18_10463_out0 };
assign v$CARRY_6584_out0 = v$C23_16760_out0;
assign v$CARRY_6587_out0 = v$C23_16763_out0;
assign v$ENDr_7844_out0 = v$A20_16994_out1;
assign v$ENDr_7847_out0 = v$A20_16997_out1;
assign v$_7876_out0 = { v$C8_19109_out0,v$C9_12718_out0 };
assign v$_7879_out0 = { v$C8_19112_out0,v$C9_12721_out0 };
assign v$ENDi_9032_out0 = v$A15_13799_out1;
assign v$ENDi_9035_out0 = v$A15_13802_out1;
assign v$END0_9723_out0 = v$A16A_15160_out1;
assign v$END0_9726_out0 = v$A16A_15163_out1;
assign v$G7_10115_out0 = v$G8_12023_out0 && v$P$CD_11004_out0;
assign v$G7_10122_out0 = v$G8_12030_out0 && v$P$CD_11011_out0;
assign v$G7_10126_out0 = v$G8_12034_out0 && v$P$CD_11015_out0;
assign v$G7_10129_out0 = v$G8_12037_out0 && v$P$CD_11018_out0;
assign v$G7_10137_out0 = v$G8_12045_out0 && v$P$CD_11026_out0;
assign v$G7_10238_out0 = v$G8_12146_out0 && v$P$CD_11127_out0;
assign v$G7_10245_out0 = v$G8_12153_out0 && v$P$CD_11134_out0;
assign v$G7_10249_out0 = v$G8_12157_out0 && v$P$CD_11138_out0;
assign v$G7_10252_out0 = v$G8_12160_out0 && v$P$CD_11141_out0;
assign v$G7_10260_out0 = v$G8_12168_out0 && v$P$CD_11149_out0;
assign v$_10691_out0 = { v$C12_9769_out0,v$C13_19199_out0 };
assign v$_10694_out0 = { v$C12_9772_out0,v$C13_19202_out0 };
assign v$ENDt_10713_out0 = v$A13_7556_out1;
assign v$ENDt_10716_out0 = v$A13_7559_out1;
assign v$_10818_out0 = { v$_14022_out0,v$_19275_out0 };
assign v$_10821_out0 = { v$_14025_out0,v$_19278_out0 };
assign v$_11465_out0 = { v$A16A_15160_out0,v$A12A_4615_out0 };
assign v$_11468_out0 = { v$A16A_15163_out0,v$A12A_4618_out0 };
assign v$_15448_out0 = { v$C10_2105_out0,v$C11_9889_out0 };
assign v$_15451_out0 = { v$C10_2108_out0,v$C11_9892_out0 };
assign v$G$AD_17775_out0 = v$G4_11701_out0;
assign v$G$AD_17794_out0 = v$G4_11720_out0;
assign v$G$AD_17898_out0 = v$G4_11824_out0;
assign v$G$AD_17917_out0 = v$G4_11843_out0;
assign v$_18100_out0 = { v$A20_16994_out0,v$A13_7556_out0 };
assign v$_18103_out0 = { v$A20_16997_out0,v$A13_7559_out0 };
assign v$ENDe_18506_out0 = v$A18_10460_out1;
assign v$ENDe_18509_out0 = v$A18_10463_out1;
assign v$G6_550_out0 = v$G4_11708_out0 || v$G7_10115_out0;
assign v$G6_557_out0 = v$G4_11715_out0 || v$G7_10122_out0;
assign v$G6_561_out0 = v$G4_11719_out0 || v$G7_10126_out0;
assign v$G6_564_out0 = v$G4_11722_out0 || v$G7_10129_out0;
assign v$G6_572_out0 = v$G4_11730_out0 || v$G7_10137_out0;
assign v$G6_673_out0 = v$G4_11831_out0 || v$G7_10238_out0;
assign v$G6_680_out0 = v$G4_11838_out0 || v$G7_10245_out0;
assign v$G6_684_out0 = v$G4_11842_out0 || v$G7_10249_out0;
assign v$G6_687_out0 = v$G4_11845_out0 || v$G7_10252_out0;
assign v$G6_695_out0 = v$G4_11853_out0 || v$G7_10260_out0;
assign v$P$AD_794_out0 = v$G1_5807_out0;
assign v$P$AD_803_out0 = v$G1_5816_out0;
assign v$P$AD_804_out0 = v$G1_5817_out0;
assign v$P$AD_815_out0 = v$G1_5828_out0;
assign v$P$AD_817_out0 = v$G1_5830_out0;
assign v$P$AD_824_out0 = v$G1_5837_out0;
assign v$P$AD_825_out0 = v$G1_5838_out0;
assign v$P$AD_917_out0 = v$G1_5930_out0;
assign v$P$AD_926_out0 = v$G1_5939_out0;
assign v$P$AD_927_out0 = v$G1_5940_out0;
assign v$P$AD_938_out0 = v$G1_5951_out0;
assign v$P$AD_940_out0 = v$G1_5953_out0;
assign v$P$AD_947_out0 = v$G1_5960_out0;
assign v$P$AD_948_out0 = v$G1_5961_out0;
assign v$_1715_out0 = { v$_15632_out0,v$_11465_out0 };
assign v$_1718_out0 = { v$_15635_out0,v$_11468_out0 };
assign v$COUTD_6971_out0 = v$G6_493_out0;
assign v$COUTD_6976_out0 = v$G6_498_out0;
assign v$COUTD_6982_out0 = v$G6_504_out0;
assign v$COUTD_6985_out0 = v$G6_507_out0;
assign v$COUTD_6990_out0 = v$G6_512_out0;
assign v$COUTD_7003_out0 = v$G6_525_out0;
assign v$COUTD_7094_out0 = v$G6_616_out0;
assign v$COUTD_7099_out0 = v$G6_621_out0;
assign v$COUTD_7105_out0 = v$G6_627_out0;
assign v$COUTD_7108_out0 = v$G6_630_out0;
assign v$COUTD_7113_out0 = v$G6_635_out0;
assign v$COUTD_7126_out0 = v$G6_648_out0;
assign v$END50_7731_out0 = v$G$AD_17775_out0;
assign v$END50_7734_out0 = v$G$AD_17898_out0;
assign v$END48_10829_out0 = v$G$AD_17794_out0;
assign v$END48_10832_out0 = v$G$AD_17917_out0;
assign v$G4_11657_out0 = v$G5_4736_out0 || v$G$CD_1064_out0;
assign v$G4_11661_out0 = v$G5_4740_out0 || v$G$CD_1068_out0;
assign v$G4_11680_out0 = v$G5_4759_out0 || v$G$CD_1087_out0;
assign v$G4_11688_out0 = v$G5_4767_out0 || v$G$CD_1095_out0;
assign v$G4_11690_out0 = v$G5_4769_out0 || v$G$CD_1097_out0;
assign v$G4_11780_out0 = v$G5_4859_out0 || v$G$CD_1187_out0;
assign v$G4_11784_out0 = v$G5_4863_out0 || v$G$CD_1191_out0;
assign v$G4_11803_out0 = v$G5_4882_out0 || v$G$CD_1210_out0;
assign v$G4_11811_out0 = v$G5_4890_out0 || v$G$CD_1218_out0;
assign v$G4_11813_out0 = v$G5_4892_out0 || v$G$CD_1220_out0;
assign v$_14898_out0 = { v$_6175_out0,v$_18100_out0 };
assign v$_14901_out0 = { v$_6178_out0,v$_18103_out0 };
assign v$_18909_out0 = { v$_7876_out0,v$_15448_out0 };
assign v$_18912_out0 = { v$_7879_out0,v$_15451_out0 };
assign v$_1321_out0 = { v$_1715_out0,v$_14898_out0 };
assign v$_1324_out0 = { v$_1718_out0,v$_14901_out0 };
assign v$C4_1414_out0 = v$COUTD_6976_out0;
assign v$C4_1417_out0 = v$COUTD_7099_out0;
assign v$P$AB_2221_out0 = v$P$AD_794_out0;
assign v$P$AB_2228_out0 = v$P$AD_794_out0;
assign v$P$AB_2232_out0 = v$P$AD_815_out0;
assign v$P$AB_2235_out0 = v$P$AD_815_out0;
assign v$P$AB_2243_out0 = v$P$AD_794_out0;
assign v$P$AB_2344_out0 = v$P$AD_917_out0;
assign v$P$AB_2351_out0 = v$P$AD_917_out0;
assign v$P$AB_2355_out0 = v$P$AD_938_out0;
assign v$P$AB_2358_out0 = v$P$AD_938_out0;
assign v$P$AB_2366_out0 = v$P$AD_917_out0;
assign v$END27_2415_out0 = v$P$AD_824_out0;
assign v$END27_2418_out0 = v$P$AD_947_out0;
assign v$END21_4505_out0 = v$P$AD_804_out0;
assign v$END21_4508_out0 = v$P$AD_927_out0;
assign v$END40_6063_out0 = v$COUTD_6990_out0;
assign v$END40_6066_out0 = v$COUTD_7113_out0;
assign v$END29_6162_out0 = v$P$AD_815_out0;
assign v$END29_6165_out0 = v$P$AD_938_out0;
assign v$COUTD_7028_out0 = v$G6_550_out0;
assign v$COUTD_7035_out0 = v$G6_557_out0;
assign v$COUTD_7039_out0 = v$G6_561_out0;
assign v$COUTD_7042_out0 = v$G6_564_out0;
assign v$COUTD_7050_out0 = v$G6_572_out0;
assign v$COUTD_7151_out0 = v$G6_673_out0;
assign v$COUTD_7158_out0 = v$G6_680_out0;
assign v$COUTD_7162_out0 = v$G6_684_out0;
assign v$COUTD_7165_out0 = v$G6_687_out0;
assign v$COUTD_7173_out0 = v$G6_695_out0;
assign v$CINA_8817_out0 = v$COUTD_7003_out0;
assign v$CINA_8821_out0 = v$COUTD_7003_out0;
assign v$CINA_8840_out0 = v$COUTD_7003_out0;
assign v$CINA_8848_out0 = v$COUTD_6990_out0;
assign v$CINA_8850_out0 = v$COUTD_7003_out0;
assign v$CINA_8940_out0 = v$COUTD_7126_out0;
assign v$CINA_8944_out0 = v$COUTD_7126_out0;
assign v$CINA_8963_out0 = v$COUTD_7126_out0;
assign v$CINA_8971_out0 = v$COUTD_7113_out0;
assign v$CINA_8973_out0 = v$COUTD_7126_out0;
assign v$END4_9738_out0 = v$COUTD_6971_out0;
assign v$END4_9741_out0 = v$COUTD_7094_out0;
assign v$END52_12550_out0 = v$P$AD_817_out0;
assign v$END52_12553_out0 = v$P$AD_940_out0;
assign v$END60_15742_out0 = v$COUTD_6985_out0;
assign v$END60_15745_out0 = v$COUTD_7108_out0;
assign v$C3_16324_out0 = v$COUTD_6982_out0;
assign v$C3_16327_out0 = v$COUTD_7105_out0;
assign v$C5_16520_out0 = v$COUTD_7003_out0;
assign v$C5_16523_out0 = v$COUTD_7126_out0;
assign v$END23_17337_out0 = v$P$AD_825_out0;
assign v$END23_17340_out0 = v$P$AD_948_out0;
assign v$END25_17667_out0 = v$P$AD_803_out0;
assign v$END25_17670_out0 = v$P$AD_926_out0;
assign v$G$AD_17731_out0 = v$G4_11657_out0;
assign v$G$AD_17735_out0 = v$G4_11661_out0;
assign v$G$AD_17754_out0 = v$G4_11680_out0;
assign v$G$AD_17762_out0 = v$G4_11688_out0;
assign v$G$AD_17764_out0 = v$G4_11690_out0;
assign v$G$AD_17854_out0 = v$G4_11780_out0;
assign v$G$AD_17858_out0 = v$G4_11784_out0;
assign v$G$AD_17877_out0 = v$G4_11803_out0;
assign v$G$AD_17885_out0 = v$G4_11811_out0;
assign v$G$AD_17887_out0 = v$G4_11813_out0;
assign v$END16_223_out0 = v$G$AD_17764_out0;
assign v$END16_226_out0 = v$G$AD_17887_out0;
assign v$END14_285_out0 = v$G$AD_17735_out0;
assign v$END14_288_out0 = v$G$AD_17858_out0;
assign v$G$CD_1084_out0 = v$G$AD_17762_out0;
assign v$G$CD_1207_out0 = v$G$AD_17885_out0;
assign v$C16_1425_out0 = v$COUTD_7042_out0;
assign v$C16_1428_out0 = v$COUTD_7165_out0;
assign {v$A7A_1816_out1,v$A7A_1816_out0 } = v$A5_6902_out0 + v$B5_18979_out0 + v$C4_1414_out0;
assign {v$A7A_1819_out1,v$A7A_1819_out0 } = v$A5_6905_out0 + v$B5_18982_out0 + v$C4_1417_out0;
assign v$C4_2039_out0 = v$C4_1414_out0;
assign v$C4_2042_out0 = v$C4_1417_out0;
assign {v$A6A_3335_out1,v$A6A_3335_out0 } = v$A6_321_out0 + v$B6_13884_out0 + v$C5_16520_out0;
assign {v$A6A_3338_out1,v$A6A_3338_out0 } = v$A6_324_out0 + v$B6_13887_out0 + v$C5_16523_out0;
assign v$G1_5820_out0 = v$P$AB_2221_out0 && v$P$CD_10963_out0;
assign v$G1_5827_out0 = v$P$AB_2228_out0 && v$P$CD_10970_out0;
assign v$G1_5831_out0 = v$P$AB_2232_out0 && v$P$CD_10974_out0;
assign v$G1_5834_out0 = v$P$AB_2235_out0 && v$P$CD_10977_out0;
assign v$G1_5842_out0 = v$P$AB_2243_out0 && v$P$CD_10985_out0;
assign v$G1_5943_out0 = v$P$AB_2344_out0 && v$P$CD_11086_out0;
assign v$G1_5950_out0 = v$P$AB_2351_out0 && v$P$CD_11093_out0;
assign v$G1_5954_out0 = v$P$AB_2355_out0 && v$P$CD_11097_out0;
assign v$G1_5957_out0 = v$P$AB_2358_out0 && v$P$CD_11100_out0;
assign v$G1_5965_out0 = v$P$AB_2366_out0 && v$P$CD_11108_out0;
assign v$C15_8449_out0 = v$COUTD_7039_out0;
assign v$C15_8452_out0 = v$COUTD_7162_out0;
assign v$C19_8469_out0 = v$COUTD_7050_out0;
assign v$C19_8472_out0 = v$COUTD_7173_out0;
assign v$CINA_8861_out0 = v$COUTD_7035_out0;
assign v$CINA_8880_out0 = v$COUTD_7035_out0;
assign v$CINA_8984_out0 = v$COUTD_7158_out0;
assign v$CINA_9003_out0 = v$COUTD_7158_out0;
assign v$G$AB_9508_out0 = v$G$AD_17754_out0;
assign v$G$AB_9517_out0 = v$G$AD_17754_out0;
assign v$G$AB_9518_out0 = v$G$AD_17731_out0;
assign v$G$AB_9529_out0 = v$G$AD_17754_out0;
assign v$G$AB_9531_out0 = v$G$AD_17754_out0;
assign v$G$AB_9538_out0 = v$G$AD_17754_out0;
assign v$G$AB_9539_out0 = v$G$AD_17731_out0;
assign v$G$AB_9631_out0 = v$G$AD_17877_out0;
assign v$G$AB_9640_out0 = v$G$AD_17877_out0;
assign v$G$AB_9641_out0 = v$G$AD_17854_out0;
assign v$G$AB_9652_out0 = v$G$AD_17877_out0;
assign v$G$AB_9654_out0 = v$G$AD_17877_out0;
assign v$G$AB_9661_out0 = v$G$AD_17877_out0;
assign v$G$AB_9662_out0 = v$G$AD_17854_out0;
assign v$G8_11972_out0 = v$CINA_8817_out0 && v$P$AB_2211_out0;
assign v$G8_11976_out0 = v$CINA_8821_out0 && v$P$AB_2215_out0;
assign v$G8_11995_out0 = v$CINA_8840_out0 && v$P$AB_2234_out0;
assign v$G8_12003_out0 = v$CINA_8848_out0 && v$P$AB_2242_out0;
assign v$G8_12005_out0 = v$CINA_8850_out0 && v$P$AB_2244_out0;
assign v$G8_12095_out0 = v$CINA_8940_out0 && v$P$AB_2334_out0;
assign v$G8_12099_out0 = v$CINA_8944_out0 && v$P$AB_2338_out0;
assign v$G8_12118_out0 = v$CINA_8963_out0 && v$P$AB_2357_out0;
assign v$G8_12126_out0 = v$CINA_8971_out0 && v$P$AB_2365_out0;
assign v$G8_12128_out0 = v$CINA_8973_out0 && v$P$AB_2367_out0;
assign v$C5_12254_out0 = v$C5_16520_out0;
assign v$C5_12257_out0 = v$C5_16523_out0;
assign v$END18_12520_out0 = v$G$AD_17731_out0;
assign v$END18_12523_out0 = v$G$AD_17854_out0;
assign v$C20_16081_out0 = v$COUTD_7035_out0;
assign v$C20_16084_out0 = v$COUTD_7158_out0;
assign v$C3_16421_out0 = v$C3_16324_out0;
assign v$C3_16424_out0 = v$C3_16327_out0;
assign {v$A5A_16710_out1,v$A5A_16710_out0 } = v$A4_18139_out0 + v$B4_15267_out0 + v$C3_16324_out0;
assign {v$A5A_16713_out1,v$A5A_16713_out0 } = v$A4_18142_out0 + v$B4_15270_out0 + v$C3_16327_out0;
assign v$C18_16904_out0 = v$COUTD_7028_out0;
assign v$C18_16907_out0 = v$COUTD_7151_out0;
assign v$_18836_out0 = { v$_18360_out0,v$_1321_out0 };
assign v$_18839_out0 = { v$_18363_out0,v$_1324_out0 };
assign v$_83_out0 = { v$A5A_16710_out0,v$A7A_1816_out0 };
assign v$_86_out0 = { v$A5A_16713_out0,v$A7A_1819_out0 };
assign v$P$AD_807_out0 = v$G1_5820_out0;
assign v$P$AD_814_out0 = v$G1_5827_out0;
assign v$P$AD_818_out0 = v$G1_5831_out0;
assign v$P$AD_821_out0 = v$G1_5834_out0;
assign v$P$AD_829_out0 = v$G1_5842_out0;
assign v$P$AD_930_out0 = v$G1_5943_out0;
assign v$P$AD_937_out0 = v$G1_5950_out0;
assign v$P$AD_941_out0 = v$G1_5954_out0;
assign v$P$AD_944_out0 = v$G1_5957_out0;
assign v$P$AD_952_out0 = v$G1_5965_out0;
assign v$_2647_out0 = { v$C4_2039_out0,v$C5_12254_out0 };
assign v$_2650_out0 = { v$C4_2042_out0,v$C5_12257_out0 };
assign v$END5_4302_out0 = v$A7A_1816_out1;
assign v$END5_4305_out0 = v$A7A_1819_out1;
assign v$G5_4733_out0 = v$G$AB_9508_out0 && v$P$CD_10950_out0;
assign v$G5_4742_out0 = v$G$AB_9517_out0 && v$P$CD_10959_out0;
assign v$G5_4743_out0 = v$G$AB_9518_out0 && v$P$CD_10960_out0;
assign v$G5_4754_out0 = v$G$AB_9529_out0 && v$P$CD_10971_out0;
assign v$G5_4756_out0 = v$G$AB_9531_out0 && v$P$CD_10973_out0;
assign v$G5_4763_out0 = v$G$AB_9538_out0 && v$P$CD_10980_out0;
assign v$G5_4764_out0 = v$G$AB_9539_out0 && v$P$CD_10981_out0;
assign v$G5_4856_out0 = v$G$AB_9631_out0 && v$P$CD_11073_out0;
assign v$G5_4865_out0 = v$G$AB_9640_out0 && v$P$CD_11082_out0;
assign v$G5_4866_out0 = v$G$AB_9641_out0 && v$P$CD_11083_out0;
assign v$G5_4877_out0 = v$G$AB_9652_out0 && v$P$CD_11094_out0;
assign v$G5_4879_out0 = v$G$AB_9654_out0 && v$P$CD_11096_out0;
assign v$G5_4886_out0 = v$G$AB_9661_out0 && v$P$CD_11103_out0;
assign v$G5_4887_out0 = v$G$AB_9662_out0 && v$P$CD_11104_out0;
assign v$END4_5464_out0 = v$A5A_16710_out1;
assign v$END4_5467_out0 = v$A5A_16713_out1;
assign v$G7_10064_out0 = v$G8_11972_out0 && v$P$CD_10953_out0;
assign v$G7_10068_out0 = v$G8_11976_out0 && v$P$CD_10957_out0;
assign v$G7_10087_out0 = v$G8_11995_out0 && v$P$CD_10976_out0;
assign v$G7_10095_out0 = v$G8_12003_out0 && v$P$CD_10984_out0;
assign v$G7_10097_out0 = v$G8_12005_out0 && v$P$CD_10986_out0;
assign v$G7_10187_out0 = v$G8_12095_out0 && v$P$CD_11076_out0;
assign v$G7_10191_out0 = v$G8_12099_out0 && v$P$CD_11080_out0;
assign v$G7_10210_out0 = v$G8_12118_out0 && v$P$CD_11099_out0;
assign v$G7_10218_out0 = v$G8_12126_out0 && v$P$CD_11107_out0;
assign v$G7_10220_out0 = v$G8_12128_out0 && v$P$CD_11109_out0;
assign v$G8_12016_out0 = v$CINA_8861_out0 && v$P$AB_2255_out0;
assign v$G8_12035_out0 = v$CINA_8880_out0 && v$P$AB_2274_out0;
assign v$G8_12139_out0 = v$CINA_8984_out0 && v$P$AB_2378_out0;
assign v$G8_12158_out0 = v$CINA_9003_out0 && v$P$AB_2397_out0;
assign v$C15_13709_out0 = v$C15_8449_out0;
assign v$C15_13712_out0 = v$C15_8452_out0;
assign v$C19_14423_out0 = v$C19_8469_out0;
assign v$C19_14426_out0 = v$C19_8472_out0;
assign v$C20_15594_out0 = v$C20_16081_out0;
assign v$C20_15597_out0 = v$C20_16084_out0;
assign v$_15615_out0 = { v$C2_18778_out0,v$C3_16421_out0 };
assign v$_15618_out0 = { v$C2_18781_out0,v$C3_16424_out0 };
assign v$C16_15770_out0 = v$C16_1425_out0;
assign v$C16_15773_out0 = v$C16_1428_out0;
assign v$END6_15832_out0 = v$A6A_3335_out1;
assign v$END6_15835_out0 = v$A6A_3338_out1;
assign {v$A14_15943_out1,v$A14_15943_out0 } = v$A16_14193_out0 + v$B16_17036_out0 + v$C15_8449_out0;
assign {v$A14_15946_out1,v$A14_15946_out0 } = v$A16_14196_out0 + v$B16_17039_out0 + v$C15_8452_out0;
assign {v$A19_16513_out1,v$A19_16513_out0 } = v$A19_1365_out0 + v$B19_17412_out0 + v$C18_16904_out0;
assign {v$A19_16516_out1,v$A19_16516_out0 } = v$A19_1368_out0 + v$B19_17415_out0 + v$C18_16907_out0;
assign {v$A24_17571_out1,v$A24_17571_out0 } = v$A21_2794_out0 + v$B21_18691_out0 + v$C20_16081_out0;
assign {v$A24_17574_out1,v$A24_17574_out0 } = v$A21_2797_out0 + v$B21_18694_out0 + v$C20_16084_out0;
assign {v$A22_18129_out1,v$A22_18129_out0 } = v$A20_4605_out0 + v$B20_4114_out0 + v$C19_8469_out0;
assign {v$A22_18132_out1,v$A22_18132_out0 } = v$A20_4608_out0 + v$B20_4117_out0 + v$C19_8472_out0;
assign {v$A11_18486_out1,v$A11_18486_out0 } = v$A17_17344_out0 + v$B17_16127_out0 + v$C16_1425_out0;
assign {v$A11_18489_out1,v$A11_18489_out0 } = v$A17_17347_out0 + v$B17_16130_out0 + v$C16_1428_out0;
assign v$C18_18611_out0 = v$C18_16904_out0;
assign v$C18_18614_out0 = v$C18_16907_out0;
assign v$END33_274_out0 = v$P$AD_821_out0;
assign v$END33_277_out0 = v$P$AD_944_out0;
assign v$G6_499_out0 = v$G4_11657_out0 || v$G7_10064_out0;
assign v$G6_503_out0 = v$G4_11661_out0 || v$G7_10068_out0;
assign v$G6_522_out0 = v$G4_11680_out0 || v$G7_10087_out0;
assign v$G6_530_out0 = v$G4_11688_out0 || v$G7_10095_out0;
assign v$G6_532_out0 = v$G4_11690_out0 || v$G7_10097_out0;
assign v$G6_622_out0 = v$G4_11780_out0 || v$G7_10187_out0;
assign v$G6_626_out0 = v$G4_11784_out0 || v$G7_10191_out0;
assign v$G6_645_out0 = v$G4_11803_out0 || v$G7_10210_out0;
assign v$G6_653_out0 = v$G4_11811_out0 || v$G7_10218_out0;
assign v$G6_655_out0 = v$G4_11813_out0 || v$G7_10220_out0;
assign v$_1349_out0 = { v$A15_13799_out0,v$A19_16513_out0 };
assign v$_1352_out0 = { v$A15_13802_out0,v$A19_16516_out0 };
assign v$_1956_out0 = { v$A22_18129_out0,v$A24_17571_out0 };
assign v$_1959_out0 = { v$A22_18132_out0,v$A24_17574_out0 };
assign v$P$AB_2214_out0 = v$P$AD_814_out0;
assign v$P$AB_2233_out0 = v$P$AD_814_out0;
assign v$P$AB_2337_out0 = v$P$AD_937_out0;
assign v$P$AB_2356_out0 = v$P$AD_937_out0;
assign v$END47_2877_out0 = v$P$AD_814_out0;
assign v$END47_2880_out0 = v$P$AD_937_out0;
assign v$_3066_out0 = { v$C14_342_out0,v$C15_13709_out0 };
assign v$_3069_out0 = { v$C14_345_out0,v$C15_13712_out0 };
assign v$ENDp_3411_out0 = v$A22_18129_out1;
assign v$ENDp_3414_out0 = v$A22_18132_out1;
assign v$ENDy_4273_out0 = v$A14_15943_out1;
assign v$ENDy_4276_out0 = v$A14_15946_out1;
assign v$ENDu_7315_out0 = v$A11_18486_out1;
assign v$ENDu_7318_out0 = v$A11_18489_out1;
assign v$_7569_out0 = { v$_9236_out0,v$_15615_out0 };
assign v$_7572_out0 = { v$_9239_out0,v$_15618_out0 };
assign v$_8195_out0 = { v$C16_15770_out0,v$C17_6344_out0 };
assign v$_8198_out0 = { v$C16_15773_out0,v$C17_6347_out0 };
assign v$_8643_out0 = { v$C18_18611_out0,v$C19_14423_out0 };
assign v$_8646_out0 = { v$C18_18614_out0,v$C19_14426_out0 };
assign v$G7_10108_out0 = v$G8_12016_out0 && v$P$CD_10997_out0;
assign v$G7_10127_out0 = v$G8_12035_out0 && v$P$CD_11016_out0;
assign v$G7_10231_out0 = v$G8_12139_out0 && v$P$CD_11120_out0;
assign v$G7_10250_out0 = v$G8_12158_out0 && v$P$CD_11139_out0;
assign v$G4_11654_out0 = v$G5_4733_out0 || v$G$CD_1061_out0;
assign v$G4_11663_out0 = v$G5_4742_out0 || v$G$CD_1070_out0;
assign v$G4_11664_out0 = v$G5_4743_out0 || v$G$CD_1071_out0;
assign v$G4_11675_out0 = v$G5_4754_out0 || v$G$CD_1082_out0;
assign v$G4_11677_out0 = v$G5_4756_out0 || v$G$CD_1084_out0;
assign v$G4_11684_out0 = v$G5_4763_out0 || v$G$CD_1091_out0;
assign v$G4_11685_out0 = v$G5_4764_out0 || v$G$CD_1092_out0;
assign v$G4_11777_out0 = v$G5_4856_out0 || v$G$CD_1184_out0;
assign v$G4_11786_out0 = v$G5_4865_out0 || v$G$CD_1193_out0;
assign v$G4_11787_out0 = v$G5_4866_out0 || v$G$CD_1194_out0;
assign v$G4_11798_out0 = v$G5_4877_out0 || v$G$CD_1205_out0;
assign v$G4_11800_out0 = v$G5_4879_out0 || v$G$CD_1207_out0;
assign v$G4_11807_out0 = v$G5_4886_out0 || v$G$CD_1214_out0;
assign v$G4_11808_out0 = v$G5_4887_out0 || v$G$CD_1215_out0;
assign v$_13879_out0 = { v$A14_15943_out0,v$A11_18486_out0 };
assign v$_13882_out0 = { v$A14_15946_out0,v$A11_18489_out0 };
assign v$END44_16259_out0 = v$P$AD_829_out0;
assign v$END44_16262_out0 = v$P$AD_952_out0;
assign v$ENDa_17185_out0 = v$A24_17571_out1;
assign v$ENDa_17188_out0 = v$A24_17574_out1;
assign v$END42_18917_out0 = v$P$AD_807_out0;
assign v$END42_18920_out0 = v$P$AD_930_out0;
assign v$END31_19132_out0 = v$P$AD_818_out0;
assign v$END31_19135_out0 = v$P$AD_941_out0;
assign v$ENDo_19306_out0 = v$A19_16513_out1;
assign v$ENDo_19309_out0 = v$A19_16516_out1;
assign v$G6_543_out0 = v$G4_11701_out0 || v$G7_10108_out0;
assign v$G6_562_out0 = v$G4_11720_out0 || v$G7_10127_out0;
assign v$G6_666_out0 = v$G4_11824_out0 || v$G7_10231_out0;
assign v$G6_685_out0 = v$G4_11843_out0 || v$G7_10250_out0;
assign v$_1397_out0 = { v$_10691_out0,v$_3066_out0 };
assign v$_1400_out0 = { v$_10694_out0,v$_3069_out0 };
assign v$G1_5813_out0 = v$P$AB_2214_out0 && v$P$CD_10956_out0;
assign v$G1_5832_out0 = v$P$AB_2233_out0 && v$P$CD_10975_out0;
assign v$G1_5936_out0 = v$P$AB_2337_out0 && v$P$CD_11079_out0;
assign v$G1_5955_out0 = v$P$AB_2356_out0 && v$P$CD_11098_out0;
assign v$COUTD_6977_out0 = v$G6_499_out0;
assign v$COUTD_6981_out0 = v$G6_503_out0;
assign v$COUTD_7000_out0 = v$G6_522_out0;
assign v$COUTD_7008_out0 = v$G6_530_out0;
assign v$COUTD_7010_out0 = v$G6_532_out0;
assign v$COUTD_7100_out0 = v$G6_622_out0;
assign v$COUTD_7104_out0 = v$G6_626_out0;
assign v$COUTD_7123_out0 = v$G6_645_out0;
assign v$COUTD_7131_out0 = v$G6_653_out0;
assign v$COUTD_7133_out0 = v$G6_655_out0;
assign v$_10813_out0 = { v$_8195_out0,v$_8643_out0 };
assign v$_10816_out0 = { v$_8198_out0,v$_8646_out0 };
assign v$_16868_out0 = { v$_13879_out0,v$_1349_out0 };
assign v$_16871_out0 = { v$_13882_out0,v$_1352_out0 };
assign v$G$AD_17728_out0 = v$G4_11654_out0;
assign v$G$AD_17737_out0 = v$G4_11663_out0;
assign v$G$AD_17738_out0 = v$G4_11664_out0;
assign v$G$AD_17749_out0 = v$G4_11675_out0;
assign v$G$AD_17751_out0 = v$G4_11677_out0;
assign v$G$AD_17758_out0 = v$G4_11684_out0;
assign v$G$AD_17759_out0 = v$G4_11685_out0;
assign v$G$AD_17851_out0 = v$G4_11777_out0;
assign v$G$AD_17860_out0 = v$G4_11786_out0;
assign v$G$AD_17861_out0 = v$G4_11787_out0;
assign v$G$AD_17872_out0 = v$G4_11798_out0;
assign v$G$AD_17874_out0 = v$G4_11800_out0;
assign v$G$AD_17881_out0 = v$G4_11807_out0;
assign v$G$AD_17882_out0 = v$G4_11808_out0;
assign v$END53_331_out0 = v$G$AD_17751_out0;
assign v$END53_334_out0 = v$G$AD_17874_out0;
assign v$P$AD_800_out0 = v$G1_5813_out0;
assign v$P$AD_819_out0 = v$G1_5832_out0;
assign v$P$AD_923_out0 = v$G1_5936_out0;
assign v$P$AD_942_out0 = v$G1_5955_out0;
assign v$END26_6679_out0 = v$G$AD_17758_out0;
assign v$END26_6682_out0 = v$G$AD_17881_out0;
assign v$COUTD_7021_out0 = v$G6_543_out0;
assign v$COUTD_7040_out0 = v$G6_562_out0;
assign v$COUTD_7144_out0 = v$G6_666_out0;
assign v$COUTD_7163_out0 = v$G6_685_out0;
assign v$C8_7749_out0 = v$COUTD_6977_out0;
assign v$C8_7752_out0 = v$COUTD_7100_out0;
assign v$CINA_8814_out0 = v$COUTD_7000_out0;
assign v$CINA_8823_out0 = v$COUTD_7000_out0;
assign v$CINA_8824_out0 = v$COUTD_6977_out0;
assign v$CINA_8835_out0 = v$COUTD_7000_out0;
assign v$CINA_8837_out0 = v$COUTD_7000_out0;
assign v$CINA_8844_out0 = v$COUTD_7000_out0;
assign v$CINA_8845_out0 = v$COUTD_6977_out0;
assign v$CINA_8937_out0 = v$COUTD_7123_out0;
assign v$CINA_8946_out0 = v$COUTD_7123_out0;
assign v$CINA_8947_out0 = v$COUTD_7100_out0;
assign v$CINA_8958_out0 = v$COUTD_7123_out0;
assign v$CINA_8960_out0 = v$COUTD_7123_out0;
assign v$CINA_8967_out0 = v$COUTD_7123_out0;
assign v$CINA_8968_out0 = v$COUTD_7100_out0;
assign v$G$AB_9521_out0 = v$G$AD_17728_out0;
assign v$G$AB_9528_out0 = v$G$AD_17728_out0;
assign v$G$AB_9532_out0 = v$G$AD_17749_out0;
assign v$G$AB_9535_out0 = v$G$AD_17749_out0;
assign v$G$AB_9543_out0 = v$G$AD_17728_out0;
assign v$G$AB_9644_out0 = v$G$AD_17851_out0;
assign v$G$AB_9651_out0 = v$G$AD_17851_out0;
assign v$G$AB_9655_out0 = v$G$AD_17872_out0;
assign v$G$AB_9658_out0 = v$G$AD_17872_out0;
assign v$G$AB_9666_out0 = v$G$AD_17851_out0;
assign v$C6_9967_out0 = v$COUTD_6981_out0;
assign v$C6_9970_out0 = v$COUTD_7104_out0;
assign v$C7_11476_out0 = v$COUTD_7010_out0;
assign v$C7_11479_out0 = v$COUTD_7133_out0;
assign v$END20_13848_out0 = v$G$AD_17738_out0;
assign v$END20_13851_out0 = v$G$AD_17861_out0;
assign v$END28_14249_out0 = v$G$AD_17749_out0;
assign v$END28_14252_out0 = v$G$AD_17872_out0;
assign v$C11_15405_out0 = v$COUTD_7000_out0;
assign v$C11_15408_out0 = v$COUTD_7123_out0;
assign v$END22_16074_out0 = v$G$AD_17759_out0;
assign v$END22_16077_out0 = v$G$AD_17882_out0;
assign v$END24_17023_out0 = v$G$AD_17737_out0;
assign v$END24_17026_out0 = v$G$AD_17860_out0;
assign v$_17997_out0 = { v$_18909_out0,v$_1397_out0 };
assign v$_18000_out0 = { v$_18912_out0,v$_1400_out0 };
assign v$END61_18571_out0 = v$COUTD_7008_out0;
assign v$END61_18574_out0 = v$COUTD_7131_out0;
assign {v$A8A_1660_out1,v$A8A_1660_out0 } = v$A7_15892_out0 + v$B7_17635_out0 + v$C6_9967_out0;
assign {v$A8A_1663_out1,v$A8A_1663_out0 } = v$A7_15895_out0 + v$B7_17638_out0 + v$C6_9970_out0;
assign {v$A17A_2683_out1,v$A17A_2683_out0 } = v$A12_3356_out0 + v$B12_2115_out0 + v$C11_15405_out0;
assign {v$A17A_2686_out1,v$A17A_2686_out0 } = v$A12_3359_out0 + v$B12_2118_out0 + v$C11_15408_out0;
assign v$G5_4746_out0 = v$G$AB_9521_out0 && v$P$CD_10963_out0;
assign v$G5_4753_out0 = v$G$AB_9528_out0 && v$P$CD_10970_out0;
assign v$G5_4757_out0 = v$G$AB_9532_out0 && v$P$CD_10974_out0;
assign v$G5_4760_out0 = v$G$AB_9535_out0 && v$P$CD_10977_out0;
assign v$G5_4768_out0 = v$G$AB_9543_out0 && v$P$CD_10985_out0;
assign v$G5_4869_out0 = v$G$AB_9644_out0 && v$P$CD_11086_out0;
assign v$G5_4876_out0 = v$G$AB_9651_out0 && v$P$CD_11093_out0;
assign v$G5_4880_out0 = v$G$AB_9655_out0 && v$P$CD_11097_out0;
assign v$G5_4883_out0 = v$G$AB_9658_out0 && v$P$CD_11100_out0;
assign v$G5_4891_out0 = v$G$AB_9666_out0 && v$P$CD_11108_out0;
assign v$_5084_out0 = { v$_8114_out0,v$_17997_out0 };
assign v$_5087_out0 = { v$_8117_out0,v$_18000_out0 };
assign v$C6_7342_out0 = v$C6_9967_out0;
assign v$C6_7345_out0 = v$C6_9970_out0;
assign v$C11_9888_out0 = v$C11_15405_out0;
assign v$C11_9891_out0 = v$C11_15408_out0;
assign {v$A9A_10863_out1,v$A9A_10863_out0 } = v$A8_18698_out0 + v$B8_13716_out0 + v$C7_11476_out0;
assign {v$A9A_10866_out1,v$A9A_10866_out0 } = v$A8_18701_out0 + v$B8_13719_out0 + v$C7_11479_out0;
assign v$C21_11260_out0 = v$COUTD_7040_out0;
assign v$C21_11263_out0 = v$COUTD_7163_out0;
assign v$C22_11490_out0 = v$COUTD_7021_out0;
assign v$C22_11493_out0 = v$COUTD_7144_out0;
assign v$G8_11969_out0 = v$CINA_8814_out0 && v$P$AB_2208_out0;
assign v$G8_11978_out0 = v$CINA_8823_out0 && v$P$AB_2217_out0;
assign v$G8_11979_out0 = v$CINA_8824_out0 && v$P$AB_2218_out0;
assign v$G8_11990_out0 = v$CINA_8835_out0 && v$P$AB_2229_out0;
assign v$G8_11992_out0 = v$CINA_8837_out0 && v$P$AB_2231_out0;
assign v$G8_11999_out0 = v$CINA_8844_out0 && v$P$AB_2238_out0;
assign v$G8_12000_out0 = v$CINA_8845_out0 && v$P$AB_2239_out0;
assign v$G8_12092_out0 = v$CINA_8937_out0 && v$P$AB_2331_out0;
assign v$G8_12101_out0 = v$CINA_8946_out0 && v$P$AB_2340_out0;
assign v$G8_12102_out0 = v$CINA_8947_out0 && v$P$AB_2341_out0;
assign v$G8_12113_out0 = v$CINA_8958_out0 && v$P$AB_2352_out0;
assign v$G8_12115_out0 = v$CINA_8960_out0 && v$P$AB_2354_out0;
assign v$G8_12122_out0 = v$CINA_8967_out0 && v$P$AB_2361_out0;
assign v$G8_12123_out0 = v$CINA_8968_out0 && v$P$AB_2362_out0;
assign v$END51_12243_out0 = v$P$AD_800_out0;
assign v$END51_12246_out0 = v$P$AD_923_out0;
assign {v$A10A_16613_out1,v$A10A_16613_out0 } = v$A9_3644_out0 + v$B9_4221_out0 + v$C8_7749_out0;
assign {v$A10A_16616_out1,v$A10A_16616_out0 } = v$A9_3647_out0 + v$B9_4224_out0 + v$C8_7752_out0;
assign v$C7_17052_out0 = v$C7_11476_out0;
assign v$C7_17055_out0 = v$C7_11479_out0;
assign v$END49_19060_out0 = v$P$AD_819_out0;
assign v$END49_19063_out0 = v$P$AD_942_out0;
assign v$C8_19108_out0 = v$C8_7749_out0;
assign v$C8_19111_out0 = v$C8_7752_out0;
assign v$END7_3583_out0 = v$A8A_1660_out1;
assign v$END7_3586_out0 = v$A8A_1663_out1;
assign v$_3827_out0 = { v$A6A_3335_out0,v$A8A_1660_out0 };
assign v$_3830_out0 = { v$A6A_3338_out0,v$A8A_1663_out0 };
assign v$END8_4071_out0 = v$A9A_10863_out1;
assign v$END8_4074_out0 = v$A9A_10866_out1;
assign v$END9_4393_out0 = v$A10A_16613_out1;
assign v$END9_4396_out0 = v$A10A_16616_out1;
assign v$C21_6610_out0 = v$C21_11260_out0;
assign v$C21_6613_out0 = v$C21_11263_out0;
assign v$C22_8716_out0 = v$C22_11490_out0;
assign v$C22_8719_out0 = v$C22_11493_out0;
assign {v$A23_9926_out1,v$A23_9926_out0 } = v$A23_5283_out0 + v$B23_1443_out0 + v$C22_11490_out0;
assign {v$A23_9929_out1,v$A23_9929_out0 } = v$A23_5286_out0 + v$B23_1446_out0 + v$C22_11493_out0;
assign v$ENDw_9931_out0 = v$A17A_2683_out1;
assign v$ENDw_9934_out0 = v$A17A_2686_out1;
assign v$G7_10061_out0 = v$G8_11969_out0 && v$P$CD_10950_out0;
assign v$G7_10070_out0 = v$G8_11978_out0 && v$P$CD_10959_out0;
assign v$G7_10071_out0 = v$G8_11979_out0 && v$P$CD_10960_out0;
assign v$G7_10082_out0 = v$G8_11990_out0 && v$P$CD_10971_out0;
assign v$G7_10084_out0 = v$G8_11992_out0 && v$P$CD_10973_out0;
assign v$G7_10091_out0 = v$G8_11999_out0 && v$P$CD_10980_out0;
assign v$G7_10092_out0 = v$G8_12000_out0 && v$P$CD_10981_out0;
assign v$G7_10184_out0 = v$G8_12092_out0 && v$P$CD_11073_out0;
assign v$G7_10193_out0 = v$G8_12101_out0 && v$P$CD_11082_out0;
assign v$G7_10194_out0 = v$G8_12102_out0 && v$P$CD_11083_out0;
assign v$G7_10205_out0 = v$G8_12113_out0 && v$P$CD_11094_out0;
assign v$G7_10207_out0 = v$G8_12115_out0 && v$P$CD_11096_out0;
assign v$G7_10214_out0 = v$G8_12122_out0 && v$P$CD_11103_out0;
assign v$G7_10215_out0 = v$G8_12123_out0 && v$P$CD_11104_out0;
assign v$G4_11667_out0 = v$G5_4746_out0 || v$G$CD_1074_out0;
assign v$G4_11674_out0 = v$G5_4753_out0 || v$G$CD_1081_out0;
assign v$G4_11678_out0 = v$G5_4757_out0 || v$G$CD_1085_out0;
assign v$G4_11681_out0 = v$G5_4760_out0 || v$G$CD_1088_out0;
assign v$G4_11689_out0 = v$G5_4768_out0 || v$G$CD_1096_out0;
assign v$G4_11790_out0 = v$G5_4869_out0 || v$G$CD_1197_out0;
assign v$G4_11797_out0 = v$G5_4876_out0 || v$G$CD_1204_out0;
assign v$G4_11801_out0 = v$G5_4880_out0 || v$G$CD_1208_out0;
assign v$G4_11804_out0 = v$G5_4883_out0 || v$G$CD_1211_out0;
assign v$G4_11812_out0 = v$G5_4891_out0 || v$G$CD_1219_out0;
assign v$_15631_out0 = { v$A9A_10863_out0,v$A10A_16613_out0 };
assign v$_15634_out0 = { v$A9A_10866_out0,v$A10A_16616_out0 };
assign v$_16925_out0 = { v$C6_7342_out0,v$C7_17052_out0 };
assign v$_16928_out0 = { v$C6_7345_out0,v$C7_17055_out0 };
assign {v$A21_19181_out1,v$A21_19181_out0 } = v$A22_4592_out0 + v$B22_11302_out0 + v$C21_11260_out0;
assign {v$A21_19184_out1,v$A21_19184_out0 } = v$A22_4595_out0 + v$B22_11305_out0 + v$C21_11263_out0;
assign v$G6_496_out0 = v$G4_11654_out0 || v$G7_10061_out0;
assign v$G6_505_out0 = v$G4_11663_out0 || v$G7_10070_out0;
assign v$G6_506_out0 = v$G4_11664_out0 || v$G7_10071_out0;
assign v$G6_517_out0 = v$G4_11675_out0 || v$G7_10082_out0;
assign v$G6_519_out0 = v$G4_11677_out0 || v$G7_10084_out0;
assign v$G6_526_out0 = v$G4_11684_out0 || v$G7_10091_out0;
assign v$G6_527_out0 = v$G4_11685_out0 || v$G7_10092_out0;
assign v$G6_619_out0 = v$G4_11777_out0 || v$G7_10184_out0;
assign v$G6_628_out0 = v$G4_11786_out0 || v$G7_10193_out0;
assign v$G6_629_out0 = v$G4_11787_out0 || v$G7_10194_out0;
assign v$G6_640_out0 = v$G4_11798_out0 || v$G7_10205_out0;
assign v$G6_642_out0 = v$G4_11800_out0 || v$G7_10207_out0;
assign v$G6_649_out0 = v$G4_11807_out0 || v$G7_10214_out0;
assign v$G6_650_out0 = v$G4_11808_out0 || v$G7_10215_out0;
assign v$_712_out0 = { v$C20_15594_out0,v$C21_6610_out0 };
assign v$_715_out0 = { v$C20_15597_out0,v$C21_6613_out0 };
assign v$_1735_out0 = { v$A21_19181_out0,v$A23_9926_out0 };
assign v$_1738_out0 = { v$A21_19184_out0,v$A23_9929_out0 };
assign v$ENDs_3437_out0 = v$A21_19181_out1;
assign v$ENDs_3440_out0 = v$A21_19184_out1;
assign v$_7720_out0 = { v$_2647_out0,v$_16925_out0 };
assign v$_7723_out0 = { v$_2650_out0,v$_16928_out0 };
assign v$ENDd_11332_out0 = v$A23_9926_out1;
assign v$ENDd_11335_out0 = v$A23_9929_out1;
assign v$_16305_out0 = { v$C22_8716_out0,v$C23_16760_out0 };
assign v$_16308_out0 = { v$C22_8719_out0,v$C23_16763_out0 };
assign v$G$AD_17741_out0 = v$G4_11667_out0;
assign v$G$AD_17748_out0 = v$G4_11674_out0;
assign v$G$AD_17752_out0 = v$G4_11678_out0;
assign v$G$AD_17755_out0 = v$G4_11681_out0;
assign v$G$AD_17763_out0 = v$G4_11689_out0;
assign v$G$AD_17864_out0 = v$G4_11790_out0;
assign v$G$AD_17871_out0 = v$G4_11797_out0;
assign v$G$AD_17875_out0 = v$G4_11801_out0;
assign v$G$AD_17878_out0 = v$G4_11804_out0;
assign v$G$AD_17886_out0 = v$G4_11812_out0;
assign v$_18580_out0 = { v$_83_out0,v$_3827_out0 };
assign v$_18583_out0 = { v$_86_out0,v$_3830_out0 };
assign v$END32_2665_out0 = v$G$AD_17755_out0;
assign v$END32_2668_out0 = v$G$AD_17878_out0;
assign v$COUTD_6974_out0 = v$G6_496_out0;
assign v$COUTD_6983_out0 = v$G6_505_out0;
assign v$COUTD_6984_out0 = v$G6_506_out0;
assign v$COUTD_6995_out0 = v$G6_517_out0;
assign v$COUTD_6997_out0 = v$G6_519_out0;
assign v$COUTD_7004_out0 = v$G6_526_out0;
assign v$COUTD_7005_out0 = v$G6_527_out0;
assign v$COUTD_7097_out0 = v$G6_619_out0;
assign v$COUTD_7106_out0 = v$G6_628_out0;
assign v$COUTD_7107_out0 = v$G6_629_out0;
assign v$COUTD_7118_out0 = v$G6_640_out0;
assign v$COUTD_7120_out0 = v$G6_642_out0;
assign v$COUTD_7127_out0 = v$G6_649_out0;
assign v$COUTD_7128_out0 = v$G6_650_out0;
assign v$_8113_out0 = { v$_7569_out0,v$_7720_out0 };
assign v$_8116_out0 = { v$_7572_out0,v$_7723_out0 };
assign v$G$AB_9514_out0 = v$G$AD_17748_out0;
assign v$G$AB_9533_out0 = v$G$AD_17748_out0;
assign v$G$AB_9637_out0 = v$G$AD_17871_out0;
assign v$G$AB_9656_out0 = v$G$AD_17871_out0;
assign v$_9867_out0 = { v$_1956_out0,v$_1735_out0 };
assign v$_9870_out0 = { v$_1959_out0,v$_1738_out0 };
assign v$END43_13772_out0 = v$G$AD_17763_out0;
assign v$END43_13775_out0 = v$G$AD_17886_out0;
assign v$_14316_out0 = { v$_712_out0,v$_16305_out0 };
assign v$_14319_out0 = { v$_715_out0,v$_16308_out0 };
assign v$END46_15664_out0 = v$G$AD_17748_out0;
assign v$END46_15667_out0 = v$G$AD_17871_out0;
assign v$END30_16310_out0 = v$G$AD_17752_out0;
assign v$END30_16313_out0 = v$G$AD_17875_out0;
assign v$END41_17287_out0 = v$G$AD_17741_out0;
assign v$END41_17290_out0 = v$G$AD_17864_out0;
assign v$_18359_out0 = { v$_10818_out0,v$_18580_out0 };
assign v$_18362_out0 = { v$_10821_out0,v$_18583_out0 };
assign v$C14_291_out0 = v$COUTD_6995_out0;
assign v$C14_294_out0 = v$COUTD_7118_out0;
assign v$C17_2717_out0 = v$COUTD_6974_out0;
assign v$C17_2720_out0 = v$COUTD_7097_out0;
assign v$_4250_out0 = { v$_10813_out0,v$_14316_out0 };
assign v$_4253_out0 = { v$_10816_out0,v$_14319_out0 };
assign v$G5_4739_out0 = v$G$AB_9514_out0 && v$P$CD_10956_out0;
assign v$G5_4758_out0 = v$G$AB_9533_out0 && v$P$CD_10975_out0;
assign v$G5_4862_out0 = v$G$AB_9637_out0 && v$P$CD_11079_out0;
assign v$G5_4881_out0 = v$G$AB_9656_out0 && v$P$CD_11098_out0;
assign v$C23_5057_out0 = v$COUTD_6997_out0;
assign v$C23_5060_out0 = v$COUTD_7120_out0;
assign v$C9_6217_out0 = v$COUTD_6984_out0;
assign v$C9_6220_out0 = v$COUTD_7107_out0;
assign v$_6895_out0 = { v$_16868_out0,v$_9867_out0 };
assign v$_6898_out0 = { v$_16871_out0,v$_9870_out0 };
assign v$CINA_8827_out0 = v$COUTD_6974_out0;
assign v$CINA_8834_out0 = v$COUTD_6974_out0;
assign v$CINA_8838_out0 = v$COUTD_6995_out0;
assign v$CINA_8841_out0 = v$COUTD_6995_out0;
assign v$CINA_8849_out0 = v$COUTD_6974_out0;
assign v$CINA_8950_out0 = v$COUTD_7097_out0;
assign v$CINA_8957_out0 = v$COUTD_7097_out0;
assign v$CINA_8961_out0 = v$COUTD_7118_out0;
assign v$CINA_8964_out0 = v$COUTD_7118_out0;
assign v$CINA_8972_out0 = v$COUTD_7097_out0;
assign v$C13_12347_out0 = v$COUTD_7004_out0;
assign v$C13_12350_out0 = v$COUTD_7127_out0;
assign v$C10_13302_out0 = v$COUTD_7005_out0;
assign v$C10_13305_out0 = v$COUTD_7128_out0;
assign v$C12_14095_out0 = v$COUTD_6983_out0;
assign v$C12_14098_out0 = v$COUTD_7106_out0;
assign v$C14_341_out0 = v$C14_291_out0;
assign v$C14_344_out0 = v$C14_294_out0;
assign v$C10_2104_out0 = v$C10_13302_out0;
assign v$C10_2107_out0 = v$C10_13305_out0;
assign v$_3941_out0 = { v$_5084_out0,v$_4250_out0 };
assign v$_3944_out0 = { v$_5087_out0,v$_4253_out0 };
assign {v$A12A_4614_out1,v$A12A_4614_out0 } = v$A11_10387_out0 + v$B11_9444_out0 + v$C10_13302_out0;
assign {v$A12A_4617_out1,v$A12A_4617_out0 } = v$A11_10390_out0 + v$B11_9447_out0 + v$C10_13305_out0;
assign v$C17_6343_out0 = v$C17_2717_out0;
assign v$C17_6346_out0 = v$C17_2720_out0;
assign {v$A13_7555_out1,v$A13_7555_out0 } = v$A15_17958_out0 + v$B15_10447_out0 + v$C14_291_out0;
assign {v$A13_7558_out1,v$A13_7558_out0 } = v$A15_17961_out0 + v$B15_10450_out0 + v$C14_294_out0;
assign v$C12_9768_out0 = v$C12_14095_out0;
assign v$C12_9771_out0 = v$C12_14098_out0;
assign v$_10329_out0 = { v$_18836_out0,v$_6895_out0 };
assign v$_10332_out0 = { v$_18839_out0,v$_6898_out0 };
assign {v$A18_10459_out1,v$A18_10459_out0 } = v$A13_14446_out0 + v$B13_9023_out0 + v$C12_14095_out0;
assign {v$A18_10462_out1,v$A18_10462_out0 } = v$A13_14449_out0 + v$B13_9026_out0 + v$C12_14098_out0;
assign v$G4_11660_out0 = v$G5_4739_out0 || v$G$CD_1067_out0;
assign v$G4_11679_out0 = v$G5_4758_out0 || v$G$CD_1086_out0;
assign v$G4_11783_out0 = v$G5_4862_out0 || v$G$CD_1190_out0;
assign v$G4_11802_out0 = v$G5_4881_out0 || v$G$CD_1209_out0;
assign v$G8_11982_out0 = v$CINA_8827_out0 && v$P$AB_2221_out0;
assign v$G8_11989_out0 = v$CINA_8834_out0 && v$P$AB_2228_out0;
assign v$G8_11993_out0 = v$CINA_8838_out0 && v$P$AB_2232_out0;
assign v$G8_11996_out0 = v$CINA_8841_out0 && v$P$AB_2235_out0;
assign v$G8_12004_out0 = v$CINA_8849_out0 && v$P$AB_2243_out0;
assign v$G8_12105_out0 = v$CINA_8950_out0 && v$P$AB_2344_out0;
assign v$G8_12112_out0 = v$CINA_8957_out0 && v$P$AB_2351_out0;
assign v$G8_12116_out0 = v$CINA_8961_out0 && v$P$AB_2355_out0;
assign v$G8_12119_out0 = v$CINA_8964_out0 && v$P$AB_2358_out0;
assign v$G8_12127_out0 = v$CINA_8972_out0 && v$P$AB_2366_out0;
assign v$C9_12717_out0 = v$C9_6217_out0;
assign v$C9_12720_out0 = v$C9_6220_out0;
assign {v$A15_13798_out1,v$A15_13798_out0 } = v$A18_18301_out0 + v$B18_11369_out0 + v$C17_2717_out0;
assign {v$A15_13801_out1,v$A15_13801_out0 } = v$A18_18304_out0 + v$B18_11372_out0 + v$C17_2720_out0;
assign {v$A16A_15159_out1,v$A16A_15159_out0 } = v$A10_1704_out0 + v$B10_10298_out0 + v$C9_6217_out0;
assign {v$A16A_15162_out1,v$A16A_15162_out0 } = v$A10_1707_out0 + v$B10_10301_out0 + v$C9_6220_out0;
assign v$C23_16759_out0 = v$C23_5057_out0;
assign v$C23_16762_out0 = v$C23_5060_out0;
assign {v$A20_16993_out1,v$A20_16993_out0 } = v$A14_739_out0 + v$B14_4159_out0 + v$C13_12347_out0;
assign {v$A20_16996_out1,v$A20_16996_out0 } = v$A14_742_out0 + v$B14_4162_out0 + v$C13_12350_out0;
assign v$C13_19198_out0 = v$C13_12347_out0;
assign v$C13_19201_out0 = v$C13_12350_out0;
assign v$ENDq_1610_out0 = v$A12A_4614_out1;
assign v$ENDq_1613_out0 = v$A12A_4617_out1;
assign v$_6174_out0 = { v$A17A_2683_out0,v$A18_10459_out0 };
assign v$_6177_out0 = { v$A17A_2686_out0,v$A18_10462_out0 };
assign v$CARRY_6583_out0 = v$C23_16759_out0;
assign v$CARRY_6586_out0 = v$C23_16762_out0;
assign v$ENDr_7843_out0 = v$A20_16993_out1;
assign v$ENDr_7846_out0 = v$A20_16996_out1;
assign v$_7875_out0 = { v$C8_19108_out0,v$C9_12717_out0 };
assign v$_7878_out0 = { v$C8_19111_out0,v$C9_12720_out0 };
assign v$ENDi_9031_out0 = v$A15_13798_out1;
assign v$ENDi_9034_out0 = v$A15_13801_out1;
assign v$END0_9722_out0 = v$A16A_15159_out1;
assign v$END0_9725_out0 = v$A16A_15162_out1;
assign v$SUM_9733_out0 = v$_10329_out0;
assign v$SUM_9736_out0 = v$_10332_out0;
assign v$G7_10074_out0 = v$G8_11982_out0 && v$P$CD_10963_out0;
assign v$G7_10081_out0 = v$G8_11989_out0 && v$P$CD_10970_out0;
assign v$G7_10085_out0 = v$G8_11993_out0 && v$P$CD_10974_out0;
assign v$G7_10088_out0 = v$G8_11996_out0 && v$P$CD_10977_out0;
assign v$G7_10096_out0 = v$G8_12004_out0 && v$P$CD_10985_out0;
assign v$G7_10197_out0 = v$G8_12105_out0 && v$P$CD_11086_out0;
assign v$G7_10204_out0 = v$G8_12112_out0 && v$P$CD_11093_out0;
assign v$G7_10208_out0 = v$G8_12116_out0 && v$P$CD_11097_out0;
assign v$G7_10211_out0 = v$G8_12119_out0 && v$P$CD_11100_out0;
assign v$G7_10219_out0 = v$G8_12127_out0 && v$P$CD_11108_out0;
assign v$_10690_out0 = { v$C12_9768_out0,v$C13_19198_out0 };
assign v$_10693_out0 = { v$C12_9771_out0,v$C13_19201_out0 };
assign v$ENDt_10712_out0 = v$A13_7555_out1;
assign v$ENDt_10715_out0 = v$A13_7558_out1;
assign v$_11464_out0 = { v$A16A_15159_out0,v$A12A_4614_out0 };
assign v$_11467_out0 = { v$A16A_15162_out0,v$A12A_4617_out0 };
assign v$SUM1_13399_out0 = v$_3941_out0;
assign v$SUM1_13402_out0 = v$_3944_out0;
assign v$_15447_out0 = { v$C10_2104_out0,v$C11_9888_out0 };
assign v$_15450_out0 = { v$C10_2107_out0,v$C11_9891_out0 };
assign v$G$AD_17734_out0 = v$G4_11660_out0;
assign v$G$AD_17753_out0 = v$G4_11679_out0;
assign v$G$AD_17857_out0 = v$G4_11783_out0;
assign v$G$AD_17876_out0 = v$G4_11802_out0;
assign v$_18099_out0 = { v$A20_16993_out0,v$A13_7555_out0 };
assign v$_18102_out0 = { v$A20_16996_out0,v$A13_7558_out0 };
assign v$ENDe_18505_out0 = v$A18_10459_out1;
assign v$ENDe_18508_out0 = v$A18_10462_out1;
assign v$G6_509_out0 = v$G4_11667_out0 || v$G7_10074_out0;
assign v$G6_516_out0 = v$G4_11674_out0 || v$G7_10081_out0;
assign v$G6_520_out0 = v$G4_11678_out0 || v$G7_10085_out0;
assign v$G6_523_out0 = v$G4_11681_out0 || v$G7_10088_out0;
assign v$G6_531_out0 = v$G4_11689_out0 || v$G7_10096_out0;
assign v$G6_632_out0 = v$G4_11790_out0 || v$G7_10197_out0;
assign v$G6_639_out0 = v$G4_11797_out0 || v$G7_10204_out0;
assign v$G6_643_out0 = v$G4_11801_out0 || v$G7_10208_out0;
assign v$G6_646_out0 = v$G4_11804_out0 || v$G7_10211_out0;
assign v$G6_654_out0 = v$G4_11812_out0 || v$G7_10219_out0;
assign v$_1714_out0 = { v$_15631_out0,v$_11464_out0 };
assign v$_1717_out0 = { v$_15634_out0,v$_11467_out0 };
assign v$END50_7730_out0 = v$G$AD_17734_out0;
assign v$END50_7733_out0 = v$G$AD_17857_out0;
assign v$SEL4_7880_out0 = v$SUM_9733_out0[23:1];
assign v$SEL4_7881_out0 = v$SUM_9736_out0[23:1];
assign v$END48_10828_out0 = v$G$AD_17753_out0;
assign v$END48_10831_out0 = v$G$AD_17876_out0;
assign v$IGNORE_13217_out0 = v$SUM1_13399_out0;
assign v$IGNORE_13218_out0 = v$SUM1_13402_out0;
assign v$_14897_out0 = { v$_6174_out0,v$_18099_out0 };
assign v$_14900_out0 = { v$_6177_out0,v$_18102_out0 };
assign v$OVERFLOW_15590_out0 = v$CARRY_6583_out0;
assign v$OVERFLOW_15591_out0 = v$CARRY_6586_out0;
assign v$_18908_out0 = { v$_7875_out0,v$_15447_out0 };
assign v$_18911_out0 = { v$_7878_out0,v$_15450_out0 };
assign v$OVERFLOW_445_out0 = v$OVERFLOW_15590_out0;
assign v$OVERFLOW_446_out0 = v$OVERFLOW_15591_out0;
assign v$_1320_out0 = { v$_1714_out0,v$_14897_out0 };
assign v$_1323_out0 = { v$_1717_out0,v$_14900_out0 };
assign v$COUTD_6987_out0 = v$G6_509_out0;
assign v$COUTD_6994_out0 = v$G6_516_out0;
assign v$COUTD_6998_out0 = v$G6_520_out0;
assign v$COUTD_7001_out0 = v$G6_523_out0;
assign v$COUTD_7009_out0 = v$G6_531_out0;
assign v$COUTD_7110_out0 = v$G6_632_out0;
assign v$COUTD_7117_out0 = v$G6_639_out0;
assign v$COUTD_7121_out0 = v$G6_643_out0;
assign v$COUTD_7124_out0 = v$G6_646_out0;
assign v$COUTD_7132_out0 = v$G6_654_out0;
assign v$_7693_out0 = { v$SEL4_7880_out0,v$CARRY_6584_out0 };
assign v$_7694_out0 = { v$SEL4_7881_out0,v$CARRY_6587_out0 };
assign v$C16_1424_out0 = v$COUTD_7001_out0;
assign v$C16_1427_out0 = v$COUTD_7124_out0;
assign v$FINAL$RESULT_2764_out0 = v$_7693_out0;
assign v$FINAL$RESULT_2765_out0 = v$_7694_out0;
assign v$OVERFLOW_3820_out0 = v$OVERFLOW_445_out0;
assign v$OVERFLOW_3821_out0 = v$OVERFLOW_446_out0;
assign v$C15_8448_out0 = v$COUTD_6998_out0;
assign v$C15_8451_out0 = v$COUTD_7121_out0;
assign v$C19_8468_out0 = v$COUTD_7009_out0;
assign v$C19_8471_out0 = v$COUTD_7132_out0;
assign v$CINA_8820_out0 = v$COUTD_6994_out0;
assign v$CINA_8839_out0 = v$COUTD_6994_out0;
assign v$CINA_8943_out0 = v$COUTD_7117_out0;
assign v$CINA_8962_out0 = v$COUTD_7117_out0;
assign v$C20_16080_out0 = v$COUTD_6994_out0;
assign v$C20_16083_out0 = v$COUTD_7117_out0;
assign v$C18_16903_out0 = v$COUTD_6987_out0;
assign v$C18_16906_out0 = v$COUTD_7110_out0;
assign v$_18835_out0 = { v$_18359_out0,v$_1320_out0 };
assign v$_18838_out0 = { v$_18362_out0,v$_1323_out0 };
assign v$MULTIPLIER$OUT_9712_out0 = v$FINAL$RESULT_2764_out0;
assign v$MULTIPLIER$OUT_9713_out0 = v$FINAL$RESULT_2765_out0;
assign v$G8_11975_out0 = v$CINA_8820_out0 && v$P$AB_2214_out0;
assign v$G8_11994_out0 = v$CINA_8839_out0 && v$P$AB_2233_out0;
assign v$G8_12098_out0 = v$CINA_8943_out0 && v$P$AB_2337_out0;
assign v$G8_12117_out0 = v$CINA_8962_out0 && v$P$AB_2356_out0;
assign v$C15_13708_out0 = v$C15_8448_out0;
assign v$C15_13711_out0 = v$C15_8451_out0;
assign v$C19_14422_out0 = v$C19_8468_out0;
assign v$C19_14425_out0 = v$C19_8471_out0;
assign v$C20_15593_out0 = v$C20_16080_out0;
assign v$C20_15596_out0 = v$C20_16083_out0;
assign v$C16_15769_out0 = v$C16_1424_out0;
assign v$C16_15772_out0 = v$C16_1427_out0;
assign {v$A14_15942_out1,v$A14_15942_out0 } = v$A16_14192_out0 + v$B16_17035_out0 + v$C15_8448_out0;
assign {v$A14_15945_out1,v$A14_15945_out0 } = v$A16_14195_out0 + v$B16_17038_out0 + v$C15_8451_out0;
assign {v$A19_16512_out1,v$A19_16512_out0 } = v$A19_1364_out0 + v$B19_17411_out0 + v$C18_16903_out0;
assign {v$A19_16515_out1,v$A19_16515_out0 } = v$A19_1367_out0 + v$B19_17414_out0 + v$C18_16906_out0;
assign {v$A24_17570_out1,v$A24_17570_out0 } = v$A21_2793_out0 + v$B21_18690_out0 + v$C20_16080_out0;
assign {v$A24_17573_out1,v$A24_17573_out0 } = v$A21_2796_out0 + v$B21_18693_out0 + v$C20_16083_out0;
assign {v$A22_18128_out1,v$A22_18128_out0 } = v$A20_4604_out0 + v$B20_4113_out0 + v$C19_8468_out0;
assign {v$A22_18131_out1,v$A22_18131_out0 } = v$A20_4607_out0 + v$B20_4116_out0 + v$C19_8471_out0;
assign {v$A11_18485_out1,v$A11_18485_out0 } = v$A17_17343_out0 + v$B17_16126_out0 + v$C16_1424_out0;
assign {v$A11_18488_out1,v$A11_18488_out0 } = v$A17_17346_out0 + v$B17_16129_out0 + v$C16_1427_out0;
assign v$C18_18610_out0 = v$C18_16903_out0;
assign v$C18_18613_out0 = v$C18_16906_out0;
assign v$OVERFLOW_19065_out0 = v$OVERFLOW_3820_out0;
assign v$OVERFLOW_19066_out0 = v$OVERFLOW_3821_out0;
assign v$OVERFLOW_19137_out0 = v$OVERFLOW_3820_out0;
assign v$OVERFLOW_19138_out0 = v$OVERFLOW_3821_out0;
assign v$_1348_out0 = { v$A15_13798_out0,v$A19_16512_out0 };
assign v$_1351_out0 = { v$A15_13801_out0,v$A19_16515_out0 };
assign v$_1955_out0 = { v$A22_18128_out0,v$A24_17570_out0 };
assign v$_1958_out0 = { v$A22_18131_out0,v$A24_17573_out0 };
assign v$_3065_out0 = { v$C14_341_out0,v$C15_13708_out0 };
assign v$_3068_out0 = { v$C14_344_out0,v$C15_13711_out0 };
assign v$ENDp_3410_out0 = v$A22_18128_out1;
assign v$ENDp_3413_out0 = v$A22_18131_out1;
assign v$ENDy_4272_out0 = v$A14_15942_out1;
assign v$ENDy_4275_out0 = v$A14_15945_out1;
assign v$ENDu_7314_out0 = v$A11_18485_out1;
assign v$ENDu_7317_out0 = v$A11_18488_out1;
assign v$_8194_out0 = { v$C16_15769_out0,v$C17_6343_out0 };
assign v$_8197_out0 = { v$C16_15772_out0,v$C17_6346_out0 };
assign v$_8642_out0 = { v$C18_18610_out0,v$C19_14422_out0 };
assign v$_8645_out0 = { v$C18_18613_out0,v$C19_14425_out0 };
assign v$G7_10067_out0 = v$G8_11975_out0 && v$P$CD_10956_out0;
assign v$G7_10086_out0 = v$G8_11994_out0 && v$P$CD_10975_out0;
assign v$G7_10190_out0 = v$G8_12098_out0 && v$P$CD_11079_out0;
assign v$G7_10209_out0 = v$G8_12117_out0 && v$P$CD_11098_out0;
assign v$IN_11584_out0 = v$MULTIPLIER$OUT_9712_out0;
assign v$IN_11585_out0 = v$MULTIPLIER$OUT_9712_out0;
assign v$IN_11586_out0 = v$MULTIPLIER$OUT_9713_out0;
assign v$IN_11587_out0 = v$MULTIPLIER$OUT_9713_out0;
assign {v$A1_12374_out1,v$A1_12374_out0 } = v$C1_7742_out0 + v$EXPONENT_16622_out0 + v$OVERFLOW_19137_out0;
assign {v$A1_12375_out1,v$A1_12375_out0 } = v$C1_7743_out0 + v$EXPONENT_16623_out0 + v$OVERFLOW_19138_out0;
assign v$_13878_out0 = { v$A14_15942_out0,v$A11_18485_out0 };
assign v$_13881_out0 = { v$A14_15945_out0,v$A11_18488_out0 };
assign {v$A1_16363_out1,v$A1_16363_out0 } = v$C1_14599_out0 + v$EXPONENT_14267_out0 + v$OVERFLOW_19065_out0;
assign {v$A1_16364_out1,v$A1_16364_out0 } = v$C1_14600_out0 + v$EXPONENT_14268_out0 + v$OVERFLOW_19066_out0;
assign v$ENDa_17184_out0 = v$A24_17570_out1;
assign v$ENDa_17187_out0 = v$A24_17573_out1;
assign v$ENDo_19305_out0 = v$A19_16512_out1;
assign v$ENDo_19308_out0 = v$A19_16515_out1;
assign v$OUT_170_out0 = v$A1_12374_out0;
assign v$OUT_171_out0 = v$A1_12375_out0;
assign v$G6_502_out0 = v$G4_11660_out0 || v$G7_10067_out0;
assign v$G6_521_out0 = v$G4_11679_out0 || v$G7_10086_out0;
assign v$G6_625_out0 = v$G4_11783_out0 || v$G7_10190_out0;
assign v$G6_644_out0 = v$G4_11802_out0 || v$G7_10209_out0;
assign v$_1396_out0 = { v$_10690_out0,v$_3065_out0 };
assign v$_1399_out0 = { v$_10693_out0,v$_3068_out0 };
assign v$NOT$USED_3098_out0 = v$A1_12374_out1;
assign v$NOT$USED_3099_out0 = v$A1_12375_out1;
assign v$NOT$USED_5689_out0 = v$A1_16363_out1;
assign v$NOT$USED_5690_out0 = v$A1_16364_out1;
assign v$_10812_out0 = { v$_8194_out0,v$_8642_out0 };
assign v$_10815_out0 = { v$_8197_out0,v$_8645_out0 };
assign v$IN_12204_out0 = v$IN_11584_out0;
assign v$IN_12205_out0 = v$IN_11585_out0;
assign v$IN_12206_out0 = v$IN_11586_out0;
assign v$IN_12207_out0 = v$IN_11587_out0;
assign v$OUT_15386_out0 = v$A1_16363_out0;
assign v$OUT_15387_out0 = v$A1_16364_out0;
assign v$_16867_out0 = { v$_13878_out0,v$_1348_out0 };
assign v$_16870_out0 = { v$_13881_out0,v$_1351_out0 };
assign v$COUTD_6980_out0 = v$G6_502_out0;
assign v$COUTD_6999_out0 = v$G6_521_out0;
assign v$COUTD_7103_out0 = v$G6_625_out0;
assign v$COUTD_7122_out0 = v$G6_644_out0;
assign v$IN_8605_out0 = v$IN_12204_out0;
assign v$IN_8606_out0 = v$IN_12205_out0;
assign v$IN_8607_out0 = v$IN_12206_out0;
assign v$IN_8608_out0 = v$IN_12207_out0;
assign v$IN_14140_out0 = v$IN_12204_out0;
assign v$IN_14142_out0 = v$IN_12205_out0;
assign v$IN_14144_out0 = v$IN_12206_out0;
assign v$IN_14146_out0 = v$IN_12207_out0;
assign v$_17996_out0 = { v$_18908_out0,v$_1396_out0 };
assign v$_17999_out0 = { v$_18911_out0,v$_1399_out0 };
assign v$IN_18864_out0 = v$IN_12204_out0;
assign v$IN_18865_out0 = v$IN_12205_out0;
assign v$IN_18866_out0 = v$IN_12206_out0;
assign v$IN_18867_out0 = v$IN_12207_out0;
assign v$IN_4348_out0 = v$IN_8605_out0;
assign v$IN_4349_out0 = v$IN_8606_out0;
assign v$IN_4350_out0 = v$IN_8607_out0;
assign v$IN_4351_out0 = v$IN_8608_out0;
assign v$_5083_out0 = { v$_8113_out0,v$_17996_out0 };
assign v$_5086_out0 = { v$_8116_out0,v$_17999_out0 };
assign v$IN_5380_out0 = v$IN_18864_out0;
assign v$IN_5390_out0 = v$IN_18865_out0;
assign v$IN_5411_out0 = v$IN_18866_out0;
assign v$IN_5421_out0 = v$IN_18867_out0;
assign v$SEL2_6634_out0 = v$IN_14140_out0[23:8];
assign v$SEL2_6635_out0 = v$IN_14142_out0[23:8];
assign v$SEL2_6636_out0 = v$IN_14144_out0[23:8];
assign v$SEL2_6637_out0 = v$IN_14146_out0[23:8];
assign v$C21_11259_out0 = v$COUTD_6999_out0;
assign v$C21_11262_out0 = v$COUTD_7122_out0;
assign v$C22_11489_out0 = v$COUTD_6980_out0;
assign v$C22_11492_out0 = v$COUTD_7103_out0;
assign v$SEL1_17306_out0 = v$IN_14140_out0[7:0];
assign v$SEL1_17308_out0 = v$IN_14142_out0[7:0];
assign v$SEL1_17310_out0 = v$IN_14144_out0[7:0];
assign v$SEL1_17312_out0 = v$IN_14146_out0[7:0];
assign v$IN_4039_out0 = v$IN_5380_out0;
assign v$IN_4042_out0 = v$IN_5390_out0;
assign v$IN_4048_out0 = v$IN_5411_out0;
assign v$IN_4051_out0 = v$IN_5421_out0;
assign v$SEL15_5102_out0 = v$IN_4348_out0[9:9];
assign v$SEL15_5103_out0 = v$IN_4349_out0[9:9];
assign v$SEL15_5104_out0 = v$IN_4350_out0[9:9];
assign v$SEL15_5105_out0 = v$IN_4351_out0[9:9];
assign v$C21_6609_out0 = v$C21_11259_out0;
assign v$C21_6612_out0 = v$C21_11262_out0;
assign v$SEL13_7205_out0 = v$IN_4348_out0[11:11];
assign v$SEL13_7206_out0 = v$IN_4349_out0[11:11];
assign v$SEL13_7207_out0 = v$IN_4350_out0[11:11];
assign v$SEL13_7208_out0 = v$IN_4351_out0[11:11];
assign v$SEL1_7378_out0 = v$IN_4348_out0[23:23];
assign v$SEL1_7379_out0 = v$IN_4349_out0[23:23];
assign v$SEL1_7380_out0 = v$IN_4350_out0[23:23];
assign v$SEL1_7381_out0 = v$IN_4351_out0[23:23];
assign v$SEL11_7539_out0 = v$IN_4348_out0[13:13];
assign v$SEL11_7540_out0 = v$IN_4349_out0[13:13];
assign v$SEL11_7541_out0 = v$IN_4350_out0[13:13];
assign v$SEL11_7542_out0 = v$IN_4351_out0[13:13];
assign v$SEL4_7639_out0 = v$IN_4348_out0[20:20];
assign v$SEL4_7640_out0 = v$IN_4349_out0[20:20];
assign v$SEL4_7641_out0 = v$IN_4350_out0[20:20];
assign v$SEL4_7642_out0 = v$IN_4351_out0[20:20];
assign v$SEL22_7712_out0 = v$IN_4348_out0[2:2];
assign v$SEL22_7713_out0 = v$IN_4349_out0[2:2];
assign v$SEL22_7714_out0 = v$IN_4350_out0[2:2];
assign v$SEL22_7715_out0 = v$IN_4351_out0[2:2];
assign v$SEL23_7945_out0 = v$IN_4348_out0[1:1];
assign v$SEL23_7946_out0 = v$IN_4349_out0[1:1];
assign v$SEL23_7947_out0 = v$IN_4350_out0[1:1];
assign v$SEL23_7948_out0 = v$IN_4351_out0[1:1];
assign v$SEL20_8483_out0 = v$IN_4348_out0[4:4];
assign v$SEL20_8484_out0 = v$IN_4349_out0[4:4];
assign v$SEL20_8485_out0 = v$IN_4350_out0[4:4];
assign v$SEL20_8486_out0 = v$IN_4351_out0[4:4];
assign v$C22_8715_out0 = v$C22_11489_out0;
assign v$C22_8718_out0 = v$C22_11492_out0;
assign v$SEL10_9883_out0 = v$IN_4348_out0[16:16];
assign v$SEL10_9884_out0 = v$IN_4349_out0[16:16];
assign v$SEL10_9885_out0 = v$IN_4350_out0[16:16];
assign v$SEL10_9886_out0 = v$IN_4351_out0[16:16];
assign {v$A23_9925_out1,v$A23_9925_out0 } = v$A23_5282_out0 + v$B23_1442_out0 + v$C22_11489_out0;
assign {v$A23_9928_out1,v$A23_9928_out0 } = v$A23_5285_out0 + v$B23_1445_out0 + v$C22_11492_out0;
assign v$SEL9_10717_out0 = v$IN_4348_out0[14:14];
assign v$SEL9_10718_out0 = v$IN_4349_out0[14:14];
assign v$SEL9_10719_out0 = v$IN_4350_out0[14:14];
assign v$SEL9_10720_out0 = v$IN_4351_out0[14:14];
assign v$SEL21_11560_out0 = v$IN_4348_out0[3:3];
assign v$SEL21_11561_out0 = v$IN_4349_out0[3:3];
assign v$SEL21_11562_out0 = v$IN_4350_out0[3:3];
assign v$SEL21_11563_out0 = v$IN_4351_out0[3:3];
assign v$SEL18_11908_out0 = v$IN_4348_out0[6:6];
assign v$SEL18_11909_out0 = v$IN_4349_out0[6:6];
assign v$SEL18_11910_out0 = v$IN_4350_out0[6:6];
assign v$SEL18_11911_out0 = v$IN_4351_out0[6:6];
assign v$SEL3_12298_out0 = v$IN_4348_out0[21:21];
assign v$SEL3_12299_out0 = v$IN_4349_out0[21:21];
assign v$SEL3_12300_out0 = v$IN_4350_out0[21:21];
assign v$SEL3_12301_out0 = v$IN_4351_out0[21:21];
assign v$SEL6_13066_out0 = v$IN_4348_out0[18:18];
assign v$SEL6_13067_out0 = v$IN_4349_out0[18:18];
assign v$SEL6_13068_out0 = v$IN_4350_out0[18:18];
assign v$SEL6_13069_out0 = v$IN_4351_out0[18:18];
assign v$SEL19_13385_out0 = v$IN_4348_out0[5:5];
assign v$SEL19_13386_out0 = v$IN_4349_out0[5:5];
assign v$SEL19_13387_out0 = v$IN_4350_out0[5:5];
assign v$SEL19_13388_out0 = v$IN_4351_out0[5:5];
assign v$SEL2_13906_out0 = v$IN_4348_out0[22:22];
assign v$SEL2_13907_out0 = v$IN_4349_out0[22:22];
assign v$SEL2_13908_out0 = v$IN_4350_out0[22:22];
assign v$SEL2_13909_out0 = v$IN_4351_out0[22:22];
assign v$IN_14141_out0 = v$SEL2_6634_out0;
assign v$IN_14143_out0 = v$SEL2_6635_out0;
assign v$IN_14145_out0 = v$SEL2_6636_out0;
assign v$IN_14147_out0 = v$SEL2_6637_out0;
assign v$SEL12_14433_out0 = v$IN_4348_out0[12:12];
assign v$SEL12_14434_out0 = v$IN_4349_out0[12:12];
assign v$SEL12_14435_out0 = v$IN_4350_out0[12:12];
assign v$SEL12_14436_out0 = v$IN_4351_out0[12:12];
assign v$SEL7_14936_out0 = v$IN_4348_out0[17:17];
assign v$SEL7_14937_out0 = v$IN_4349_out0[17:17];
assign v$SEL7_14938_out0 = v$IN_4350_out0[17:17];
assign v$SEL7_14939_out0 = v$IN_4351_out0[17:17];
assign v$IN_15468_out0 = v$SEL1_17306_out0;
assign v$IN_15469_out0 = v$SEL1_17308_out0;
assign v$IN_15473_out0 = v$SEL1_17310_out0;
assign v$IN_15474_out0 = v$SEL1_17312_out0;
assign v$SEL5_16038_out0 = v$IN_4348_out0[19:19];
assign v$SEL5_16039_out0 = v$IN_4349_out0[19:19];
assign v$SEL5_16040_out0 = v$IN_4350_out0[19:19];
assign v$SEL5_16041_out0 = v$IN_4351_out0[19:19];
assign v$SEL17_16683_out0 = v$IN_4348_out0[7:7];
assign v$SEL17_16684_out0 = v$IN_4349_out0[7:7];
assign v$SEL17_16685_out0 = v$IN_4350_out0[7:7];
assign v$SEL17_16686_out0 = v$IN_4351_out0[7:7];
assign v$SEL14_16964_out0 = v$IN_4348_out0[10:10];
assign v$SEL14_16965_out0 = v$IN_4349_out0[10:10];
assign v$SEL14_16966_out0 = v$IN_4350_out0[10:10];
assign v$SEL14_16967_out0 = v$IN_4351_out0[10:10];
assign v$SEL16_17505_out0 = v$IN_4348_out0[8:8];
assign v$SEL16_17506_out0 = v$IN_4349_out0[8:8];
assign v$SEL16_17507_out0 = v$IN_4350_out0[8:8];
assign v$SEL16_17508_out0 = v$IN_4351_out0[8:8];
assign v$SEL24_17529_out0 = v$IN_4348_out0[0:0];
assign v$SEL24_17530_out0 = v$IN_4349_out0[0:0];
assign v$SEL24_17531_out0 = v$IN_4350_out0[0:0];
assign v$SEL24_17532_out0 = v$IN_4351_out0[0:0];
assign v$SEL8_18285_out0 = v$IN_4348_out0[15:15];
assign v$SEL8_18286_out0 = v$IN_4349_out0[15:15];
assign v$SEL8_18287_out0 = v$IN_4350_out0[15:15];
assign v$SEL8_18288_out0 = v$IN_4351_out0[15:15];
assign {v$A21_19180_out1,v$A21_19180_out0 } = v$A22_4591_out0 + v$B22_11301_out0 + v$C21_11259_out0;
assign {v$A21_19183_out1,v$A21_19183_out0 } = v$A22_4594_out0 + v$B22_11304_out0 + v$C21_11262_out0;
assign v$_711_out0 = { v$C20_15593_out0,v$C21_6609_out0 };
assign v$_714_out0 = { v$C20_15596_out0,v$C21_6612_out0 };
assign v$_1734_out0 = { v$A21_19180_out0,v$A23_9925_out0 };
assign v$_1737_out0 = { v$A21_19183_out0,v$A23_9928_out0 };
assign v$SEL2_3238_out0 = v$IN_15468_out0[7:4];
assign v$SEL2_3239_out0 = v$IN_15469_out0[7:4];
assign v$SEL2_3243_out0 = v$IN_15473_out0[7:4];
assign v$SEL2_3244_out0 = v$IN_15474_out0[7:4];
assign v$ENDs_3436_out0 = v$A21_19180_out1;
assign v$ENDs_3439_out0 = v$A21_19183_out1;
assign v$SEL4_3592_out0 = v$IN_14141_out0[15:12];
assign v$SEL4_3593_out0 = v$IN_14143_out0[15:12];
assign v$SEL4_3594_out0 = v$IN_14145_out0[15:12];
assign v$SEL4_3595_out0 = v$IN_14147_out0[15:12];
assign v$SEL3_7683_out0 = v$IN_14141_out0[11:8];
assign v$SEL3_7684_out0 = v$IN_14143_out0[11:8];
assign v$SEL3_7685_out0 = v$IN_14145_out0[11:8];
assign v$SEL3_7686_out0 = v$IN_14147_out0[11:8];
assign v$SEL1_9061_out0 = v$IN_4039_out0[23:1];
assign v$SEL1_9071_out0 = v$IN_4042_out0[23:1];
assign v$SEL1_9092_out0 = v$IN_4048_out0[23:1];
assign v$SEL1_9102_out0 = v$IN_4051_out0[23:1];
assign v$ENDd_11331_out0 = v$A23_9925_out1;
assign v$ENDd_11334_out0 = v$A23_9928_out1;
assign v$SEL2_14439_out0 = v$IN_14141_out0[7:4];
assign v$SEL2_14440_out0 = v$IN_14143_out0[7:4];
assign v$SEL2_14441_out0 = v$IN_14145_out0[7:4];
assign v$SEL2_14442_out0 = v$IN_14147_out0[7:4];
assign v$SEL1_15989_out0 = v$IN_4039_out0[22:0];
assign v$SEL1_15999_out0 = v$IN_4042_out0[22:0];
assign v$SEL1_16020_out0 = v$IN_4048_out0[22:0];
assign v$SEL1_16030_out0 = v$IN_4051_out0[22:0];
assign v$_16304_out0 = { v$C22_8715_out0,v$C23_16759_out0 };
assign v$_16307_out0 = { v$C22_8718_out0,v$C23_16762_out0 };
assign v$SEL1_17082_out0 = v$IN_15468_out0[3:0];
assign v$SEL1_17083_out0 = v$IN_15469_out0[3:0];
assign v$SEL1_17087_out0 = v$IN_15473_out0[3:0];
assign v$SEL1_17088_out0 = v$IN_15474_out0[3:0];
assign v$SEL1_17307_out0 = v$IN_14141_out0[3:0];
assign v$SEL1_17309_out0 = v$IN_14143_out0[3:0];
assign v$SEL1_17311_out0 = v$IN_14145_out0[3:0];
assign v$SEL1_17313_out0 = v$IN_14147_out0[3:0];
assign v$MUX24_18661_out0 = v$EQ24_2732_out0 ? v$SEL24_17529_out0 : v$C1_16317_out0;
assign v$MUX24_18662_out0 = v$EQ24_2733_out0 ? v$SEL24_17530_out0 : v$C1_16318_out0;
assign v$MUX24_18663_out0 = v$EQ24_2734_out0 ? v$SEL24_17531_out0 : v$C1_16319_out0;
assign v$MUX24_18664_out0 = v$EQ24_2735_out0 ? v$SEL24_17532_out0 : v$C1_16320_out0;
assign v$_4421_out0 = { v$C2_119_out0,v$SEL1_15989_out0 };
assign v$_4431_out0 = { v$C2_129_out0,v$SEL1_15999_out0 };
assign v$_4452_out0 = { v$C2_150_out0,v$SEL1_16020_out0 };
assign v$_4462_out0 = { v$C2_160_out0,v$SEL1_16030_out0 };
assign v$_9322_out0 = { v$SEL1_9061_out0,v$C1_6257_out0 };
assign v$_9332_out0 = { v$SEL1_9071_out0,v$C1_6267_out0 };
assign v$_9353_out0 = { v$SEL1_9092_out0,v$C1_6288_out0 };
assign v$_9363_out0 = { v$SEL1_9102_out0,v$C1_6298_out0 };
assign v$_9866_out0 = { v$_1955_out0,v$_1734_out0 };
assign v$_9869_out0 = { v$_1958_out0,v$_1737_out0 };
assign v$_14315_out0 = { v$_711_out0,v$_16304_out0 };
assign v$_14318_out0 = { v$_714_out0,v$_16307_out0 };
assign v$IN_15683_out0 = v$SEL3_7683_out0;
assign v$IN_15684_out0 = v$SEL1_17307_out0;
assign v$IN_15685_out0 = v$SEL2_14439_out0;
assign v$IN_15686_out0 = v$SEL4_3592_out0;
assign v$IN_15687_out0 = v$SEL1_17082_out0;
assign v$IN_15688_out0 = v$SEL2_3238_out0;
assign v$IN_15689_out0 = v$SEL3_7684_out0;
assign v$IN_15690_out0 = v$SEL1_17309_out0;
assign v$IN_15691_out0 = v$SEL2_14440_out0;
assign v$IN_15692_out0 = v$SEL4_3593_out0;
assign v$IN_15693_out0 = v$SEL1_17083_out0;
assign v$IN_15694_out0 = v$SEL2_3239_out0;
assign v$IN_15701_out0 = v$SEL3_7685_out0;
assign v$IN_15702_out0 = v$SEL1_17311_out0;
assign v$IN_15703_out0 = v$SEL2_14441_out0;
assign v$IN_15704_out0 = v$SEL4_3594_out0;
assign v$IN_15705_out0 = v$SEL1_17087_out0;
assign v$IN_15706_out0 = v$SEL2_3243_out0;
assign v$IN_15707_out0 = v$SEL3_7686_out0;
assign v$IN_15708_out0 = v$SEL1_17313_out0;
assign v$IN_15709_out0 = v$SEL2_14442_out0;
assign v$IN_15710_out0 = v$SEL4_3595_out0;
assign v$IN_15711_out0 = v$SEL1_17088_out0;
assign v$IN_15712_out0 = v$SEL2_3244_out0;
assign v$MUX23_16833_out0 = v$EQ23_3415_out0 ? v$SEL23_7945_out0 : v$MUX24_18661_out0;
assign v$MUX23_16834_out0 = v$EQ23_3416_out0 ? v$SEL23_7946_out0 : v$MUX24_18662_out0;
assign v$MUX23_16835_out0 = v$EQ23_3417_out0 ? v$SEL23_7947_out0 : v$MUX24_18663_out0;
assign v$MUX23_16836_out0 = v$EQ23_3418_out0 ? v$SEL23_7948_out0 : v$MUX24_18664_out0;
assign v$SEL3_2505_out0 = v$IN_15683_out0[2:2];
assign v$SEL3_2506_out0 = v$IN_15684_out0[2:2];
assign v$SEL3_2507_out0 = v$IN_15685_out0[2:2];
assign v$SEL3_2508_out0 = v$IN_15686_out0[2:2];
assign v$SEL3_2509_out0 = v$IN_15687_out0[2:2];
assign v$SEL3_2510_out0 = v$IN_15688_out0[2:2];
assign v$SEL3_2511_out0 = v$IN_15689_out0[2:2];
assign v$SEL3_2512_out0 = v$IN_15690_out0[2:2];
assign v$SEL3_2513_out0 = v$IN_15691_out0[2:2];
assign v$SEL3_2514_out0 = v$IN_15692_out0[2:2];
assign v$SEL3_2515_out0 = v$IN_15693_out0[2:2];
assign v$SEL3_2516_out0 = v$IN_15694_out0[2:2];
assign v$SEL3_2523_out0 = v$IN_15701_out0[2:2];
assign v$SEL3_2524_out0 = v$IN_15702_out0[2:2];
assign v$SEL3_2525_out0 = v$IN_15703_out0[2:2];
assign v$SEL3_2526_out0 = v$IN_15704_out0[2:2];
assign v$SEL3_2527_out0 = v$IN_15705_out0[2:2];
assign v$SEL3_2528_out0 = v$IN_15706_out0[2:2];
assign v$SEL3_2529_out0 = v$IN_15707_out0[2:2];
assign v$SEL3_2530_out0 = v$IN_15708_out0[2:2];
assign v$SEL3_2531_out0 = v$IN_15709_out0[2:2];
assign v$SEL3_2532_out0 = v$IN_15710_out0[2:2];
assign v$SEL3_2533_out0 = v$IN_15711_out0[2:2];
assign v$SEL3_2534_out0 = v$IN_15712_out0[2:2];
assign v$MUX1_2558_out0 = v$LEFT$SHIT_3270_out0 ? v$_4421_out0 : v$_9322_out0;
assign v$MUX1_2568_out0 = v$LEFT$SHIT_3280_out0 ? v$_4431_out0 : v$_9332_out0;
assign v$MUX1_2589_out0 = v$LEFT$SHIT_3301_out0 ? v$_4452_out0 : v$_9353_out0;
assign v$MUX1_2599_out0 = v$LEFT$SHIT_3311_out0 ? v$_4462_out0 : v$_9363_out0;
assign v$_4249_out0 = { v$_10812_out0,v$_14315_out0 };
assign v$_4252_out0 = { v$_10815_out0,v$_14318_out0 };
assign v$SEL4_6362_out0 = v$IN_15683_out0[3:3];
assign v$SEL4_6363_out0 = v$IN_15684_out0[3:3];
assign v$SEL4_6364_out0 = v$IN_15685_out0[3:3];
assign v$SEL4_6365_out0 = v$IN_15686_out0[3:3];
assign v$SEL4_6366_out0 = v$IN_15687_out0[3:3];
assign v$SEL4_6367_out0 = v$IN_15688_out0[3:3];
assign v$SEL4_6368_out0 = v$IN_15689_out0[3:3];
assign v$SEL4_6369_out0 = v$IN_15690_out0[3:3];
assign v$SEL4_6370_out0 = v$IN_15691_out0[3:3];
assign v$SEL4_6371_out0 = v$IN_15692_out0[3:3];
assign v$SEL4_6372_out0 = v$IN_15693_out0[3:3];
assign v$SEL4_6373_out0 = v$IN_15694_out0[3:3];
assign v$SEL4_6380_out0 = v$IN_15701_out0[3:3];
assign v$SEL4_6381_out0 = v$IN_15702_out0[3:3];
assign v$SEL4_6382_out0 = v$IN_15703_out0[3:3];
assign v$SEL4_6383_out0 = v$IN_15704_out0[3:3];
assign v$SEL4_6384_out0 = v$IN_15705_out0[3:3];
assign v$SEL4_6385_out0 = v$IN_15706_out0[3:3];
assign v$SEL4_6386_out0 = v$IN_15707_out0[3:3];
assign v$SEL4_6387_out0 = v$IN_15708_out0[3:3];
assign v$SEL4_6388_out0 = v$IN_15709_out0[3:3];
assign v$SEL4_6389_out0 = v$IN_15710_out0[3:3];
assign v$SEL4_6390_out0 = v$IN_15711_out0[3:3];
assign v$SEL4_6391_out0 = v$IN_15712_out0[3:3];
assign v$_6894_out0 = { v$_16867_out0,v$_9866_out0 };
assign v$_6897_out0 = { v$_16870_out0,v$_9869_out0 };
assign v$SEL2_8005_out0 = v$IN_15683_out0[1:1];
assign v$SEL2_8006_out0 = v$IN_15684_out0[1:1];
assign v$SEL2_8007_out0 = v$IN_15685_out0[1:1];
assign v$SEL2_8008_out0 = v$IN_15686_out0[1:1];
assign v$SEL2_8009_out0 = v$IN_15687_out0[1:1];
assign v$SEL2_8010_out0 = v$IN_15688_out0[1:1];
assign v$SEL2_8011_out0 = v$IN_15689_out0[1:1];
assign v$SEL2_8012_out0 = v$IN_15690_out0[1:1];
assign v$SEL2_8013_out0 = v$IN_15691_out0[1:1];
assign v$SEL2_8014_out0 = v$IN_15692_out0[1:1];
assign v$SEL2_8015_out0 = v$IN_15693_out0[1:1];
assign v$SEL2_8016_out0 = v$IN_15694_out0[1:1];
assign v$SEL2_8023_out0 = v$IN_15701_out0[1:1];
assign v$SEL2_8024_out0 = v$IN_15702_out0[1:1];
assign v$SEL2_8025_out0 = v$IN_15703_out0[1:1];
assign v$SEL2_8026_out0 = v$IN_15704_out0[1:1];
assign v$SEL2_8027_out0 = v$IN_15705_out0[1:1];
assign v$SEL2_8028_out0 = v$IN_15706_out0[1:1];
assign v$SEL2_8029_out0 = v$IN_15707_out0[1:1];
assign v$SEL2_8030_out0 = v$IN_15708_out0[1:1];
assign v$SEL2_8031_out0 = v$IN_15709_out0[1:1];
assign v$SEL2_8032_out0 = v$IN_15710_out0[1:1];
assign v$SEL2_8033_out0 = v$IN_15711_out0[1:1];
assign v$SEL2_8034_out0 = v$IN_15712_out0[1:1];
assign v$SEL1_14050_out0 = v$IN_15683_out0[0:0];
assign v$SEL1_14051_out0 = v$IN_15684_out0[0:0];
assign v$SEL1_14052_out0 = v$IN_15685_out0[0:0];
assign v$SEL1_14053_out0 = v$IN_15686_out0[0:0];
assign v$SEL1_14054_out0 = v$IN_15687_out0[0:0];
assign v$SEL1_14055_out0 = v$IN_15688_out0[0:0];
assign v$SEL1_14056_out0 = v$IN_15689_out0[0:0];
assign v$SEL1_14057_out0 = v$IN_15690_out0[0:0];
assign v$SEL1_14058_out0 = v$IN_15691_out0[0:0];
assign v$SEL1_14059_out0 = v$IN_15692_out0[0:0];
assign v$SEL1_14060_out0 = v$IN_15693_out0[0:0];
assign v$SEL1_14061_out0 = v$IN_15694_out0[0:0];
assign v$SEL1_14068_out0 = v$IN_15701_out0[0:0];
assign v$SEL1_14069_out0 = v$IN_15702_out0[0:0];
assign v$SEL1_14070_out0 = v$IN_15703_out0[0:0];
assign v$SEL1_14071_out0 = v$IN_15704_out0[0:0];
assign v$SEL1_14072_out0 = v$IN_15705_out0[0:0];
assign v$SEL1_14073_out0 = v$IN_15706_out0[0:0];
assign v$SEL1_14074_out0 = v$IN_15707_out0[0:0];
assign v$SEL1_14075_out0 = v$IN_15708_out0[0:0];
assign v$SEL1_14076_out0 = v$IN_15709_out0[0:0];
assign v$SEL1_14077_out0 = v$IN_15710_out0[0:0];
assign v$SEL1_14078_out0 = v$IN_15711_out0[0:0];
assign v$SEL1_14079_out0 = v$IN_15712_out0[0:0];
assign v$MUX22_17090_out0 = v$EQ22_3060_out0 ? v$SEL22_7712_out0 : v$MUX23_16833_out0;
assign v$MUX22_17091_out0 = v$EQ22_3061_out0 ? v$SEL22_7713_out0 : v$MUX23_16834_out0;
assign v$MUX22_17092_out0 = v$EQ22_3062_out0 ? v$SEL22_7714_out0 : v$MUX23_16835_out0;
assign v$MUX22_17093_out0 = v$EQ22_3063_out0 ? v$SEL22_7715_out0 : v$MUX23_16836_out0;
assign v$G10_1549_out0 = !(v$SEL1_14050_out0 || v$SEL2_8005_out0);
assign v$G10_1550_out0 = !(v$SEL1_14051_out0 || v$SEL2_8006_out0);
assign v$G10_1551_out0 = !(v$SEL1_14052_out0 || v$SEL2_8007_out0);
assign v$G10_1552_out0 = !(v$SEL1_14053_out0 || v$SEL2_8008_out0);
assign v$G10_1553_out0 = !(v$SEL1_14054_out0 || v$SEL2_8009_out0);
assign v$G10_1554_out0 = !(v$SEL1_14055_out0 || v$SEL2_8010_out0);
assign v$G10_1555_out0 = !(v$SEL1_14056_out0 || v$SEL2_8011_out0);
assign v$G10_1556_out0 = !(v$SEL1_14057_out0 || v$SEL2_8012_out0);
assign v$G10_1557_out0 = !(v$SEL1_14058_out0 || v$SEL2_8013_out0);
assign v$G10_1558_out0 = !(v$SEL1_14059_out0 || v$SEL2_8014_out0);
assign v$G10_1559_out0 = !(v$SEL1_14060_out0 || v$SEL2_8015_out0);
assign v$G10_1560_out0 = !(v$SEL1_14061_out0 || v$SEL2_8016_out0);
assign v$G10_1567_out0 = !(v$SEL1_14068_out0 || v$SEL2_8023_out0);
assign v$G10_1568_out0 = !(v$SEL1_14069_out0 || v$SEL2_8024_out0);
assign v$G10_1569_out0 = !(v$SEL1_14070_out0 || v$SEL2_8025_out0);
assign v$G10_1570_out0 = !(v$SEL1_14071_out0 || v$SEL2_8026_out0);
assign v$G10_1571_out0 = !(v$SEL1_14072_out0 || v$SEL2_8027_out0);
assign v$G10_1572_out0 = !(v$SEL1_14073_out0 || v$SEL2_8028_out0);
assign v$G10_1573_out0 = !(v$SEL1_14074_out0 || v$SEL2_8029_out0);
assign v$G10_1574_out0 = !(v$SEL1_14075_out0 || v$SEL2_8030_out0);
assign v$G10_1575_out0 = !(v$SEL1_14076_out0 || v$SEL2_8031_out0);
assign v$G10_1576_out0 = !(v$SEL1_14077_out0 || v$SEL2_8032_out0);
assign v$G10_1577_out0 = !(v$SEL1_14078_out0 || v$SEL2_8033_out0);
assign v$G10_1578_out0 = !(v$SEL1_14079_out0 || v$SEL2_8034_out0);
assign v$G6_3762_out0 = ! v$SEL2_8005_out0;
assign v$G6_3763_out0 = ! v$SEL2_8006_out0;
assign v$G6_3764_out0 = ! v$SEL2_8007_out0;
assign v$G6_3765_out0 = ! v$SEL2_8008_out0;
assign v$G6_3766_out0 = ! v$SEL2_8009_out0;
assign v$G6_3767_out0 = ! v$SEL2_8010_out0;
assign v$G6_3768_out0 = ! v$SEL2_8011_out0;
assign v$G6_3769_out0 = ! v$SEL2_8012_out0;
assign v$G6_3770_out0 = ! v$SEL2_8013_out0;
assign v$G6_3771_out0 = ! v$SEL2_8014_out0;
assign v$G6_3772_out0 = ! v$SEL2_8015_out0;
assign v$G6_3773_out0 = ! v$SEL2_8016_out0;
assign v$G6_3780_out0 = ! v$SEL2_8023_out0;
assign v$G6_3781_out0 = ! v$SEL2_8024_out0;
assign v$G6_3782_out0 = ! v$SEL2_8025_out0;
assign v$G6_3783_out0 = ! v$SEL2_8026_out0;
assign v$G6_3784_out0 = ! v$SEL2_8027_out0;
assign v$G6_3785_out0 = ! v$SEL2_8028_out0;
assign v$G6_3786_out0 = ! v$SEL2_8029_out0;
assign v$G6_3787_out0 = ! v$SEL2_8030_out0;
assign v$G6_3788_out0 = ! v$SEL2_8031_out0;
assign v$G6_3789_out0 = ! v$SEL2_8032_out0;
assign v$G6_3790_out0 = ! v$SEL2_8033_out0;
assign v$G6_3791_out0 = ! v$SEL2_8034_out0;
assign v$_3940_out0 = { v$_5083_out0,v$_4249_out0 };
assign v$_3943_out0 = { v$_5086_out0,v$_4252_out0 };
assign v$MUX21_5118_out0 = v$EQ21_3547_out0 ? v$SEL21_11560_out0 : v$MUX22_17090_out0;
assign v$MUX21_5119_out0 = v$EQ21_3548_out0 ? v$SEL21_11561_out0 : v$MUX22_17091_out0;
assign v$MUX21_5120_out0 = v$EQ21_3549_out0 ? v$SEL21_11562_out0 : v$MUX22_17092_out0;
assign v$MUX21_5121_out0 = v$EQ21_3550_out0 ? v$SEL21_11563_out0 : v$MUX22_17093_out0;
assign v$G5_6125_out0 = ! v$SEL4_6362_out0;
assign v$G5_6126_out0 = ! v$SEL4_6363_out0;
assign v$G5_6127_out0 = ! v$SEL4_6364_out0;
assign v$G5_6128_out0 = ! v$SEL4_6365_out0;
assign v$G5_6129_out0 = ! v$SEL4_6366_out0;
assign v$G5_6130_out0 = ! v$SEL4_6367_out0;
assign v$G5_6131_out0 = ! v$SEL4_6368_out0;
assign v$G5_6132_out0 = ! v$SEL4_6369_out0;
assign v$G5_6133_out0 = ! v$SEL4_6370_out0;
assign v$G5_6134_out0 = ! v$SEL4_6371_out0;
assign v$G5_6135_out0 = ! v$SEL4_6372_out0;
assign v$G5_6136_out0 = ! v$SEL4_6373_out0;
assign v$G5_6143_out0 = ! v$SEL4_6380_out0;
assign v$G5_6144_out0 = ! v$SEL4_6381_out0;
assign v$G5_6145_out0 = ! v$SEL4_6382_out0;
assign v$G5_6146_out0 = ! v$SEL4_6383_out0;
assign v$G5_6147_out0 = ! v$SEL4_6384_out0;
assign v$G5_6148_out0 = ! v$SEL4_6385_out0;
assign v$G5_6149_out0 = ! v$SEL4_6386_out0;
assign v$G5_6150_out0 = ! v$SEL4_6387_out0;
assign v$G5_6151_out0 = ! v$SEL4_6388_out0;
assign v$G5_6152_out0 = ! v$SEL4_6389_out0;
assign v$G5_6153_out0 = ! v$SEL4_6390_out0;
assign v$G5_6154_out0 = ! v$SEL4_6391_out0;
assign v$G11_9195_out0 = !(v$SEL3_2505_out0 || v$SEL4_6362_out0);
assign v$G11_9196_out0 = !(v$SEL3_2506_out0 || v$SEL4_6363_out0);
assign v$G11_9197_out0 = !(v$SEL3_2507_out0 || v$SEL4_6364_out0);
assign v$G11_9198_out0 = !(v$SEL3_2508_out0 || v$SEL4_6365_out0);
assign v$G11_9199_out0 = !(v$SEL3_2509_out0 || v$SEL4_6366_out0);
assign v$G11_9200_out0 = !(v$SEL3_2510_out0 || v$SEL4_6367_out0);
assign v$G11_9201_out0 = !(v$SEL3_2511_out0 || v$SEL4_6368_out0);
assign v$G11_9202_out0 = !(v$SEL3_2512_out0 || v$SEL4_6369_out0);
assign v$G11_9203_out0 = !(v$SEL3_2513_out0 || v$SEL4_6370_out0);
assign v$G11_9204_out0 = !(v$SEL3_2514_out0 || v$SEL4_6371_out0);
assign v$G11_9205_out0 = !(v$SEL3_2515_out0 || v$SEL4_6372_out0);
assign v$G11_9206_out0 = !(v$SEL3_2516_out0 || v$SEL4_6373_out0);
assign v$G11_9213_out0 = !(v$SEL3_2523_out0 || v$SEL4_6380_out0);
assign v$G11_9214_out0 = !(v$SEL3_2524_out0 || v$SEL4_6381_out0);
assign v$G11_9215_out0 = !(v$SEL3_2525_out0 || v$SEL4_6382_out0);
assign v$G11_9216_out0 = !(v$SEL3_2526_out0 || v$SEL4_6383_out0);
assign v$G11_9217_out0 = !(v$SEL3_2527_out0 || v$SEL4_6384_out0);
assign v$G11_9218_out0 = !(v$SEL3_2528_out0 || v$SEL4_6385_out0);
assign v$G11_9219_out0 = !(v$SEL3_2529_out0 || v$SEL4_6386_out0);
assign v$G11_9220_out0 = !(v$SEL3_2530_out0 || v$SEL4_6387_out0);
assign v$G11_9221_out0 = !(v$SEL3_2531_out0 || v$SEL4_6388_out0);
assign v$G11_9222_out0 = !(v$SEL3_2532_out0 || v$SEL4_6389_out0);
assign v$G11_9223_out0 = !(v$SEL3_2533_out0 || v$SEL4_6390_out0);
assign v$G11_9224_out0 = !(v$SEL3_2534_out0 || v$SEL4_6391_out0);
assign v$_10328_out0 = { v$_18835_out0,v$_6894_out0 };
assign v$_10331_out0 = { v$_18838_out0,v$_6897_out0 };
assign v$G8_12573_out0 = ! v$SEL3_2505_out0;
assign v$G8_12574_out0 = ! v$SEL3_2506_out0;
assign v$G8_12575_out0 = ! v$SEL3_2507_out0;
assign v$G8_12576_out0 = ! v$SEL3_2508_out0;
assign v$G8_12577_out0 = ! v$SEL3_2509_out0;
assign v$G8_12578_out0 = ! v$SEL3_2510_out0;
assign v$G8_12579_out0 = ! v$SEL3_2511_out0;
assign v$G8_12580_out0 = ! v$SEL3_2512_out0;
assign v$G8_12581_out0 = ! v$SEL3_2513_out0;
assign v$G8_12582_out0 = ! v$SEL3_2514_out0;
assign v$G8_12583_out0 = ! v$SEL3_2515_out0;
assign v$G8_12584_out0 = ! v$SEL3_2516_out0;
assign v$G8_12591_out0 = ! v$SEL3_2523_out0;
assign v$G8_12592_out0 = ! v$SEL3_2524_out0;
assign v$G8_12593_out0 = ! v$SEL3_2525_out0;
assign v$G8_12594_out0 = ! v$SEL3_2526_out0;
assign v$G8_12595_out0 = ! v$SEL3_2527_out0;
assign v$G8_12596_out0 = ! v$SEL3_2528_out0;
assign v$G8_12597_out0 = ! v$SEL3_2529_out0;
assign v$G8_12598_out0 = ! v$SEL3_2530_out0;
assign v$G8_12599_out0 = ! v$SEL3_2531_out0;
assign v$G8_12600_out0 = ! v$SEL3_2532_out0;
assign v$G8_12601_out0 = ! v$SEL3_2533_out0;
assign v$G8_12602_out0 = ! v$SEL3_2534_out0;
assign v$SUM_9732_out0 = v$_10328_out0;
assign v$SUM_9735_out0 = v$_10331_out0;
assign v$MUX20_11892_out0 = v$EQ20_10370_out0 ? v$SEL20_8483_out0 : v$MUX21_5118_out0;
assign v$MUX20_11893_out0 = v$EQ20_10371_out0 ? v$SEL20_8484_out0 : v$MUX21_5119_out0;
assign v$MUX20_11894_out0 = v$EQ20_10372_out0 ? v$SEL20_8485_out0 : v$MUX21_5120_out0;
assign v$MUX20_11895_out0 = v$EQ20_10373_out0 ? v$SEL20_8486_out0 : v$MUX21_5121_out0;
assign v$G3_13250_out0 = v$G10_1549_out0 && v$G11_9195_out0;
assign v$G3_13251_out0 = v$G10_1550_out0 && v$G11_9196_out0;
assign v$G3_13252_out0 = v$G10_1551_out0 && v$G11_9197_out0;
assign v$G3_13253_out0 = v$G10_1552_out0 && v$G11_9198_out0;
assign v$G3_13254_out0 = v$G10_1553_out0 && v$G11_9199_out0;
assign v$G3_13255_out0 = v$G10_1554_out0 && v$G11_9200_out0;
assign v$G3_13256_out0 = v$G10_1555_out0 && v$G11_9201_out0;
assign v$G3_13257_out0 = v$G10_1556_out0 && v$G11_9202_out0;
assign v$G3_13258_out0 = v$G10_1557_out0 && v$G11_9203_out0;
assign v$G3_13259_out0 = v$G10_1558_out0 && v$G11_9204_out0;
assign v$G3_13260_out0 = v$G10_1559_out0 && v$G11_9205_out0;
assign v$G3_13261_out0 = v$G10_1560_out0 && v$G11_9206_out0;
assign v$G3_13268_out0 = v$G10_1567_out0 && v$G11_9213_out0;
assign v$G3_13269_out0 = v$G10_1568_out0 && v$G11_9214_out0;
assign v$G3_13270_out0 = v$G10_1569_out0 && v$G11_9215_out0;
assign v$G3_13271_out0 = v$G10_1570_out0 && v$G11_9216_out0;
assign v$G3_13272_out0 = v$G10_1571_out0 && v$G11_9217_out0;
assign v$G3_13273_out0 = v$G10_1572_out0 && v$G11_9218_out0;
assign v$G3_13274_out0 = v$G10_1573_out0 && v$G11_9219_out0;
assign v$G3_13275_out0 = v$G10_1574_out0 && v$G11_9220_out0;
assign v$G3_13276_out0 = v$G10_1575_out0 && v$G11_9221_out0;
assign v$G3_13277_out0 = v$G10_1576_out0 && v$G11_9222_out0;
assign v$G3_13278_out0 = v$G10_1577_out0 && v$G11_9223_out0;
assign v$G3_13279_out0 = v$G10_1578_out0 && v$G11_9224_out0;
assign v$SUM1_13398_out0 = v$_3940_out0;
assign v$SUM1_13401_out0 = v$_3943_out0;
assign v$G9_18217_out0 = v$G8_12573_out0 && v$G5_6125_out0;
assign v$G9_18218_out0 = v$G8_12574_out0 && v$G5_6126_out0;
assign v$G9_18219_out0 = v$G8_12575_out0 && v$G5_6127_out0;
assign v$G9_18220_out0 = v$G8_12576_out0 && v$G5_6128_out0;
assign v$G9_18221_out0 = v$G8_12577_out0 && v$G5_6129_out0;
assign v$G9_18222_out0 = v$G8_12578_out0 && v$G5_6130_out0;
assign v$G9_18223_out0 = v$G8_12579_out0 && v$G5_6131_out0;
assign v$G9_18224_out0 = v$G8_12580_out0 && v$G5_6132_out0;
assign v$G9_18225_out0 = v$G8_12581_out0 && v$G5_6133_out0;
assign v$G9_18226_out0 = v$G8_12582_out0 && v$G5_6134_out0;
assign v$G9_18227_out0 = v$G8_12583_out0 && v$G5_6135_out0;
assign v$G9_18228_out0 = v$G8_12584_out0 && v$G5_6136_out0;
assign v$G9_18235_out0 = v$G8_12591_out0 && v$G5_6143_out0;
assign v$G9_18236_out0 = v$G8_12592_out0 && v$G5_6144_out0;
assign v$G9_18237_out0 = v$G8_12593_out0 && v$G5_6145_out0;
assign v$G9_18238_out0 = v$G8_12594_out0 && v$G5_6146_out0;
assign v$G9_18239_out0 = v$G8_12595_out0 && v$G5_6147_out0;
assign v$G9_18240_out0 = v$G8_12596_out0 && v$G5_6148_out0;
assign v$G9_18241_out0 = v$G8_12597_out0 && v$G5_6149_out0;
assign v$G9_18242_out0 = v$G8_12598_out0 && v$G5_6150_out0;
assign v$G9_18243_out0 = v$G8_12599_out0 && v$G5_6151_out0;
assign v$G9_18244_out0 = v$G8_12600_out0 && v$G5_6152_out0;
assign v$G9_18245_out0 = v$G8_12601_out0 && v$G5_6153_out0;
assign v$G9_18246_out0 = v$G8_12602_out0 && v$G5_6154_out0;
assign v$G7_18747_out0 = v$G6_3762_out0 || v$SEL3_2505_out0;
assign v$G7_18748_out0 = v$G6_3763_out0 || v$SEL3_2506_out0;
assign v$G7_18749_out0 = v$G6_3764_out0 || v$SEL3_2507_out0;
assign v$G7_18750_out0 = v$G6_3765_out0 || v$SEL3_2508_out0;
assign v$G7_18751_out0 = v$G6_3766_out0 || v$SEL3_2509_out0;
assign v$G7_18752_out0 = v$G6_3767_out0 || v$SEL3_2510_out0;
assign v$G7_18753_out0 = v$G6_3768_out0 || v$SEL3_2511_out0;
assign v$G7_18754_out0 = v$G6_3769_out0 || v$SEL3_2512_out0;
assign v$G7_18755_out0 = v$G6_3770_out0 || v$SEL3_2513_out0;
assign v$G7_18756_out0 = v$G6_3771_out0 || v$SEL3_2514_out0;
assign v$G7_18757_out0 = v$G6_3772_out0 || v$SEL3_2515_out0;
assign v$G7_18758_out0 = v$G6_3773_out0 || v$SEL3_2516_out0;
assign v$G7_18765_out0 = v$G6_3780_out0 || v$SEL3_2523_out0;
assign v$G7_18766_out0 = v$G6_3781_out0 || v$SEL3_2524_out0;
assign v$G7_18767_out0 = v$G6_3782_out0 || v$SEL3_2525_out0;
assign v$G7_18768_out0 = v$G6_3783_out0 || v$SEL3_2526_out0;
assign v$G7_18769_out0 = v$G6_3784_out0 || v$SEL3_2527_out0;
assign v$G7_18770_out0 = v$G6_3785_out0 || v$SEL3_2528_out0;
assign v$G7_18771_out0 = v$G6_3786_out0 || v$SEL3_2529_out0;
assign v$G7_18772_out0 = v$G6_3787_out0 || v$SEL3_2530_out0;
assign v$G7_18773_out0 = v$G6_3788_out0 || v$SEL3_2531_out0;
assign v$G7_18774_out0 = v$G6_3789_out0 || v$SEL3_2532_out0;
assign v$G7_18775_out0 = v$G6_3790_out0 || v$SEL3_2533_out0;
assign v$G7_18776_out0 = v$G6_3791_out0 || v$SEL3_2534_out0;
assign v$SUM_2068_out0 = v$SUM_9732_out0;
assign v$SUM_2069_out0 = v$SUM_9735_out0;
assign v$MUX19_6614_out0 = v$EQ19_5682_out0 ? v$SEL19_13385_out0 : v$MUX20_11892_out0;
assign v$MUX19_6615_out0 = v$EQ19_5683_out0 ? v$SEL19_13386_out0 : v$MUX20_11893_out0;
assign v$MUX19_6616_out0 = v$EQ19_5684_out0 ? v$SEL19_13387_out0 : v$MUX20_11894_out0;
assign v$MUX19_6617_out0 = v$EQ19_5685_out0 ? v$SEL19_13388_out0 : v$MUX20_11895_out0;
assign v$END1_10352_out0 = v$SUM1_13398_out0;
assign v$END1_10353_out0 = v$SUM1_13401_out0;
assign v$Z_13153_out0 = v$G3_13250_out0;
assign v$Z_13154_out0 = v$G3_13251_out0;
assign v$Z_13155_out0 = v$G3_13252_out0;
assign v$Z_13156_out0 = v$G3_13253_out0;
assign v$Z_13157_out0 = v$G3_13254_out0;
assign v$Z_13158_out0 = v$G3_13255_out0;
assign v$Z_13159_out0 = v$G3_13256_out0;
assign v$Z_13160_out0 = v$G3_13257_out0;
assign v$Z_13161_out0 = v$G3_13258_out0;
assign v$Z_13162_out0 = v$G3_13259_out0;
assign v$Z_13163_out0 = v$G3_13260_out0;
assign v$Z_13164_out0 = v$G3_13261_out0;
assign v$Z_13171_out0 = v$G3_13268_out0;
assign v$Z_13172_out0 = v$G3_13269_out0;
assign v$Z_13173_out0 = v$G3_13270_out0;
assign v$Z_13174_out0 = v$G3_13271_out0;
assign v$Z_13175_out0 = v$G3_13272_out0;
assign v$Z_13176_out0 = v$G3_13273_out0;
assign v$Z_13177_out0 = v$G3_13274_out0;
assign v$Z_13178_out0 = v$G3_13275_out0;
assign v$Z_13179_out0 = v$G3_13276_out0;
assign v$Z_13180_out0 = v$G3_13277_out0;
assign v$Z_13181_out0 = v$G3_13278_out0;
assign v$Z_13182_out0 = v$G3_13279_out0;
assign v$SEL1_14967_out0 = v$SUM_9732_out0[23:1];
assign v$SEL1_14968_out0 = v$SUM_9735_out0[23:1];
assign v$G4_18164_out0 = v$G7_18747_out0 && v$G5_6125_out0;
assign v$G4_18165_out0 = v$G7_18748_out0 && v$G5_6126_out0;
assign v$G4_18166_out0 = v$G7_18749_out0 && v$G5_6127_out0;
assign v$G4_18167_out0 = v$G7_18750_out0 && v$G5_6128_out0;
assign v$G4_18168_out0 = v$G7_18751_out0 && v$G5_6129_out0;
assign v$G4_18169_out0 = v$G7_18752_out0 && v$G5_6130_out0;
assign v$G4_18170_out0 = v$G7_18753_out0 && v$G5_6131_out0;
assign v$G4_18171_out0 = v$G7_18754_out0 && v$G5_6132_out0;
assign v$G4_18172_out0 = v$G7_18755_out0 && v$G5_6133_out0;
assign v$G4_18173_out0 = v$G7_18756_out0 && v$G5_6134_out0;
assign v$G4_18174_out0 = v$G7_18757_out0 && v$G5_6135_out0;
assign v$G4_18175_out0 = v$G7_18758_out0 && v$G5_6136_out0;
assign v$G4_18182_out0 = v$G7_18765_out0 && v$G5_6143_out0;
assign v$G4_18183_out0 = v$G7_18766_out0 && v$G5_6144_out0;
assign v$G4_18184_out0 = v$G7_18767_out0 && v$G5_6145_out0;
assign v$G4_18185_out0 = v$G7_18768_out0 && v$G5_6146_out0;
assign v$G4_18186_out0 = v$G7_18769_out0 && v$G5_6147_out0;
assign v$G4_18187_out0 = v$G7_18770_out0 && v$G5_6148_out0;
assign v$G4_18188_out0 = v$G7_18771_out0 && v$G5_6149_out0;
assign v$G4_18189_out0 = v$G7_18772_out0 && v$G5_6150_out0;
assign v$G4_18190_out0 = v$G7_18773_out0 && v$G5_6151_out0;
assign v$G4_18191_out0 = v$G7_18774_out0 && v$G5_6152_out0;
assign v$G4_18192_out0 = v$G7_18775_out0 && v$G5_6153_out0;
assign v$G4_18193_out0 = v$G7_18776_out0 && v$G5_6154_out0;
assign v$Z2_183_out0 = v$Z_13157_out0;
assign v$Z2_184_out0 = v$Z_13163_out0;
assign v$Z2_188_out0 = v$Z_13175_out0;
assign v$Z2_189_out0 = v$Z_13181_out0;
assign v$_1665_out0 = { v$SEL1_14967_out0,v$C4_3935_out0 };
assign v$_1666_out0 = { v$SEL1_14968_out0,v$C4_3936_out0 };
assign v$MUX18_5072_out0 = v$EQ18_13375_out0 ? v$SEL18_11908_out0 : v$MUX19_6614_out0;
assign v$MUX18_5073_out0 = v$EQ18_13376_out0 ? v$SEL18_11909_out0 : v$MUX19_6615_out0;
assign v$MUX18_5074_out0 = v$EQ18_13377_out0 ? v$SEL18_11910_out0 : v$MUX19_6616_out0;
assign v$MUX18_5075_out0 = v$EQ18_13378_out0 ? v$SEL18_11911_out0 : v$MUX19_6617_out0;
assign v$XOR1_5640_out0 = v$SUM_2068_out0 ^ v$C9_15847_out0;
assign v$XOR1_5641_out0 = v$SUM_2069_out0 ^ v$C9_15848_out0;
assign v$Z1_6052_out0 = v$Z_13158_out0;
assign v$Z1_6053_out0 = v$Z_13164_out0;
assign v$Z1_6057_out0 = v$Z_13176_out0;
assign v$Z1_6058_out0 = v$Z_13182_out0;
assign v$_6538_out0 = { v$G4_18164_out0,v$G9_18217_out0 };
assign v$_6539_out0 = { v$G4_18165_out0,v$G9_18218_out0 };
assign v$_6540_out0 = { v$G4_18166_out0,v$G9_18219_out0 };
assign v$_6541_out0 = { v$G4_18167_out0,v$G9_18220_out0 };
assign v$_6542_out0 = { v$G4_18168_out0,v$G9_18221_out0 };
assign v$_6543_out0 = { v$G4_18169_out0,v$G9_18222_out0 };
assign v$_6544_out0 = { v$G4_18170_out0,v$G9_18223_out0 };
assign v$_6545_out0 = { v$G4_18171_out0,v$G9_18224_out0 };
assign v$_6546_out0 = { v$G4_18172_out0,v$G9_18225_out0 };
assign v$_6547_out0 = { v$G4_18173_out0,v$G9_18226_out0 };
assign v$_6548_out0 = { v$G4_18174_out0,v$G9_18227_out0 };
assign v$_6549_out0 = { v$G4_18175_out0,v$G9_18228_out0 };
assign v$_6556_out0 = { v$G4_18182_out0,v$G9_18235_out0 };
assign v$_6557_out0 = { v$G4_18183_out0,v$G9_18236_out0 };
assign v$_6558_out0 = { v$G4_18184_out0,v$G9_18237_out0 };
assign v$_6559_out0 = { v$G4_18185_out0,v$G9_18238_out0 };
assign v$_6560_out0 = { v$G4_18186_out0,v$G9_18239_out0 };
assign v$_6561_out0 = { v$G4_18187_out0,v$G9_18240_out0 };
assign v$_6562_out0 = { v$G4_18188_out0,v$G9_18241_out0 };
assign v$_6563_out0 = { v$G4_18189_out0,v$G9_18242_out0 };
assign v$_6564_out0 = { v$G4_18190_out0,v$G9_18243_out0 };
assign v$_6565_out0 = { v$G4_18191_out0,v$G9_18244_out0 };
assign v$_6566_out0 = { v$G4_18192_out0,v$G9_18245_out0 };
assign v$_6567_out0 = { v$G4_18193_out0,v$G9_18246_out0 };
assign v$Z2_6575_out0 = v$Z_13155_out0;
assign v$Z2_6577_out0 = v$Z_13161_out0;
assign v$Z2_6579_out0 = v$Z_13173_out0;
assign v$Z2_6581_out0 = v$Z_13179_out0;
assign v$Z4_8247_out0 = v$Z_13156_out0;
assign v$Z4_8248_out0 = v$Z_13162_out0;
assign v$Z4_8249_out0 = v$Z_13174_out0;
assign v$Z4_8250_out0 = v$Z_13180_out0;
assign v$Z1_17593_out0 = v$Z_13154_out0;
assign v$Z1_17595_out0 = v$Z_13160_out0;
assign v$Z1_17597_out0 = v$Z_13172_out0;
assign v$Z1_17599_out0 = v$Z_13178_out0;
assign v$Z3_18389_out0 = v$Z_13153_out0;
assign v$Z3_18390_out0 = v$Z_13159_out0;
assign v$Z3_18391_out0 = v$Z_13171_out0;
assign v$Z3_18392_out0 = v$Z_13177_out0;
assign v$MUX7_3505_out0 = v$OVERFLOW_15590_out0 ? v$_1665_out0 : v$SUM_2068_out0;
assign v$MUX7_3506_out0 = v$OVERFLOW_15591_out0 ? v$_1666_out0 : v$SUM_2069_out0;
assign v$G4_6334_out0 = ! v$Z4_8247_out0;
assign v$G4_6335_out0 = ! v$Z4_8248_out0;
assign v$G4_6336_out0 = ! v$Z4_8249_out0;
assign v$G4_6337_out0 = ! v$Z4_8250_out0;
assign v$G6_6435_out0 = ! v$Z2_6575_out0;
assign v$G6_6437_out0 = ! v$Z2_6577_out0;
assign v$G6_6439_out0 = ! v$Z2_6579_out0;
assign v$G6_6441_out0 = ! v$Z2_6581_out0;
assign v$Y_6737_out0 = v$_6538_out0;
assign v$Y_6738_out0 = v$_6539_out0;
assign v$Y_6739_out0 = v$_6540_out0;
assign v$Y_6740_out0 = v$_6541_out0;
assign v$Y_6741_out0 = v$_6542_out0;
assign v$Y_6742_out0 = v$_6543_out0;
assign v$Y_6743_out0 = v$_6544_out0;
assign v$Y_6744_out0 = v$_6545_out0;
assign v$Y_6745_out0 = v$_6546_out0;
assign v$Y_6746_out0 = v$_6547_out0;
assign v$Y_6747_out0 = v$_6548_out0;
assign v$Y_6748_out0 = v$_6549_out0;
assign v$Y_6755_out0 = v$_6556_out0;
assign v$Y_6756_out0 = v$_6557_out0;
assign v$Y_6757_out0 = v$_6558_out0;
assign v$Y_6758_out0 = v$_6559_out0;
assign v$Y_6759_out0 = v$_6560_out0;
assign v$Y_6760_out0 = v$_6561_out0;
assign v$Y_6761_out0 = v$_6562_out0;
assign v$Y_6762_out0 = v$_6563_out0;
assign v$Y_6763_out0 = v$_6564_out0;
assign v$Y_6764_out0 = v$_6565_out0;
assign v$Y_6765_out0 = v$_6566_out0;
assign v$Y_6766_out0 = v$_6567_out0;
assign v$A1_14170_out0 = v$XOR1_5640_out0;
assign v$A1_14173_out0 = v$XOR1_5641_out0;
assign v$G1_15194_out0 = v$Z1_6052_out0 && v$Z2_183_out0;
assign v$G1_15195_out0 = v$Z1_6053_out0 && v$Z2_184_out0;
assign v$G1_15199_out0 = v$Z1_6057_out0 && v$Z2_188_out0;
assign v$G1_15200_out0 = v$Z1_6058_out0 && v$Z2_189_out0;
assign v$G9_15798_out0 = v$Z1_17593_out0 && v$Z2_6575_out0;
assign v$G9_15800_out0 = v$Z1_17595_out0 && v$Z2_6577_out0;
assign v$G9_15802_out0 = v$Z1_17597_out0 && v$Z2_6579_out0;
assign v$G9_15804_out0 = v$Z1_17599_out0 && v$Z2_6581_out0;
assign v$MUX17_17156_out0 = v$EQ17_6155_out0 ? v$SEL17_16683_out0 : v$MUX18_5072_out0;
assign v$MUX17_17157_out0 = v$EQ17_6156_out0 ? v$SEL17_16684_out0 : v$MUX18_5073_out0;
assign v$MUX17_17158_out0 = v$EQ17_6157_out0 ? v$SEL17_16685_out0 : v$MUX18_5074_out0;
assign v$MUX17_17159_out0 = v$EQ17_6158_out0 ? v$SEL17_16686_out0 : v$MUX18_5075_out0;
assign v$G5_18148_out0 = ! v$Z3_18389_out0;
assign v$G5_18149_out0 = ! v$Z3_18390_out0;
assign v$G5_18150_out0 = ! v$Z3_18391_out0;
assign v$G5_18151_out0 = ! v$Z3_18392_out0;
assign v$_4136_out0 = { v$Y_6740_out0,v$C3_3527_out0 };
assign v$_4137_out0 = { v$Y_6746_out0,v$C3_3528_out0 };
assign v$_4138_out0 = { v$Y_6758_out0,v$C3_3529_out0 };
assign v$_4139_out0 = { v$Y_6764_out0,v$C3_3530_out0 };
assign v$_5310_out0 = { v$Y_6739_out0,v$C5_17520_out0 };
assign v$_5312_out0 = { v$Y_6745_out0,v$C5_17522_out0 };
assign v$_5314_out0 = { v$Y_6757_out0,v$C5_17524_out0 };
assign v$_5316_out0 = { v$Y_6763_out0,v$C5_17526_out0 };
assign v$_5708_out0 = { v$Y_6742_out0,v$C1_18269_out0 };
assign v$_5709_out0 = { v$Y_6748_out0,v$C1_18270_out0 };
assign v$_5713_out0 = { v$Y_6760_out0,v$C1_18274_out0 };
assign v$_5714_out0 = { v$Y_6766_out0,v$C1_18275_out0 };
assign v$_7860_out0 = v$A1_14170_out0[11:0];
assign v$_7860_out1 = v$A1_14170_out0[23:12];
assign v$_7863_out0 = v$A1_14173_out0[11:0];
assign v$_7863_out1 = v$A1_14173_out0[23:12];
assign v$_8456_out0 = { v$Y_6741_out0,v$C2_7954_out0 };
assign v$_8457_out0 = { v$Y_6747_out0,v$C2_7955_out0 };
assign v$_8461_out0 = { v$Y_6759_out0,v$C2_7959_out0 };
assign v$_8462_out0 = { v$Y_6765_out0,v$C2_7960_out0 };
assign v$_9130_out0 = { v$Y_6738_out0,v$C6_6772_out0 };
assign v$_9132_out0 = { v$Y_6744_out0,v$C6_6774_out0 };
assign v$_9134_out0 = { v$Y_6756_out0,v$C6_6776_out0 };
assign v$_9136_out0 = { v$Y_6762_out0,v$C6_6778_out0 };
assign v$_9231_out0 = { v$Y_6737_out0,v$C4_17134_out0 };
assign v$_9232_out0 = { v$Y_6743_out0,v$C4_17135_out0 };
assign v$_9233_out0 = { v$Y_6755_out0,v$C4_17136_out0 };
assign v$_9234_out0 = { v$Y_6761_out0,v$C4_17137_out0 };
assign v$G7_10275_out0 = v$G9_15798_out0 && v$Z3_18389_out0;
assign v$G7_10276_out0 = v$G9_15800_out0 && v$Z3_18390_out0;
assign v$G7_10277_out0 = v$G9_15802_out0 && v$Z3_18391_out0;
assign v$G7_10278_out0 = v$G9_15804_out0 && v$Z3_18392_out0;
assign v$Z_10790_out0 = v$G1_15194_out0;
assign v$Z_10791_out0 = v$G1_15195_out0;
assign v$Z_10795_out0 = v$G1_15199_out0;
assign v$Z_10796_out0 = v$G1_15200_out0;
assign v$SEL3_14851_out0 = v$MUX7_3505_out0[22:0];
assign v$SEL3_14852_out0 = v$MUX7_3506_out0[22:0];
assign v$MUX16_17383_out0 = v$EQ16_8597_out0 ? v$SEL16_17505_out0 : v$MUX17_17156_out0;
assign v$MUX16_17384_out0 = v$EQ16_8598_out0 ? v$SEL16_17506_out0 : v$MUX17_17157_out0;
assign v$MUX16_17385_out0 = v$EQ16_8599_out0 ? v$SEL16_17507_out0 : v$MUX17_17158_out0;
assign v$MUX16_17386_out0 = v$EQ16_8600_out0 ? v$SEL16_17508_out0 : v$MUX17_17159_out0;
assign v$MUX5_4213_out0 = v$G6_6435_out0 ? v$_5310_out0 : v$_9130_out0;
assign v$MUX5_4215_out0 = v$G6_6437_out0 ? v$_5312_out0 : v$_9132_out0;
assign v$MUX5_4217_out0 = v$G6_6439_out0 ? v$_5314_out0 : v$_9134_out0;
assign v$MUX5_4219_out0 = v$G6_6441_out0 ? v$_5316_out0 : v$_9136_out0;
assign v$LOWER$PART_6568_out0 = v$MUX16_17383_out0;
assign v$LOWER$PART_6569_out0 = v$MUX16_17384_out0;
assign v$LOWER$PART_6570_out0 = v$MUX16_17385_out0;
assign v$LOWER$PART_6571_out0 = v$MUX16_17386_out0;
assign v$MUX1_15300_out0 = v$Z1_6052_out0 ? v$_8456_out0 : v$_5708_out0;
assign v$MUX1_15301_out0 = v$Z1_6053_out0 ? v$_8457_out0 : v$_5709_out0;
assign v$MUX1_15305_out0 = v$Z1_6057_out0 ? v$_8461_out0 : v$_5713_out0;
assign v$MUX1_15306_out0 = v$Z1_6058_out0 ? v$_8462_out0 : v$_5714_out0;
assign v$_16723_out0 = v$_7860_out0[5:0];
assign v$_16723_out1 = v$_7860_out0[11:6];
assign v$_16726_out0 = v$_7863_out0[5:0];
assign v$_16726_out1 = v$_7863_out0[11:6];
assign v$G1_16754_out0 = v$G7_10275_out0 && v$Z4_8247_out0;
assign v$G1_16755_out0 = v$G7_10276_out0 && v$Z4_8248_out0;
assign v$G1_16756_out0 = v$G7_10277_out0 && v$Z4_8249_out0;
assign v$G1_16757_out0 = v$G7_10278_out0 && v$Z4_8250_out0;
assign v$Z1_17592_out0 = v$Z_10790_out0;
assign v$Z1_17594_out0 = v$Z_10791_out0;
assign v$Z1_17596_out0 = v$Z_10795_out0;
assign v$Z1_17598_out0 = v$Z_10796_out0;
assign v$_17622_out0 = v$_7860_out1[5:0];
assign v$_17622_out1 = v$_7860_out1[11:6];
assign v$_17625_out0 = v$_7863_out1[5:0];
assign v$_17625_out1 = v$_7863_out1[11:6];
assign v$MUX15_1479_out0 = v$EQ15_16574_out0 ? v$SEL15_5102_out0 : v$LOWER$PART_6568_out0;
assign v$MUX15_1480_out0 = v$EQ15_16575_out0 ? v$SEL15_5103_out0 : v$LOWER$PART_6569_out0;
assign v$MUX15_1481_out0 = v$EQ15_16576_out0 ? v$SEL15_5104_out0 : v$LOWER$PART_6570_out0;
assign v$MUX15_1482_out0 = v$EQ15_16577_out0 ? v$SEL15_5105_out0 : v$LOWER$PART_6571_out0;
assign v$_2024_out0 = v$_17622_out1[2:0];
assign v$_2024_out1 = v$_17622_out1[5:3];
assign v$_2027_out0 = v$_17625_out1[2:0];
assign v$_2027_out1 = v$_17625_out1[5:3];
assign v$Z_2748_out0 = v$G1_16754_out0;
assign v$Z_2750_out0 = v$G1_16755_out0;
assign v$Z_2752_out0 = v$G1_16756_out0;
assign v$Z_2754_out0 = v$G1_16757_out0;
assign v$MUX4_3084_out0 = v$G5_18148_out0 ? v$_9231_out0 : v$MUX5_4213_out0;
assign v$MUX4_3085_out0 = v$G5_18149_out0 ? v$_9232_out0 : v$MUX5_4215_out0;
assign v$MUX4_3086_out0 = v$G5_18150_out0 ? v$_9233_out0 : v$MUX5_4217_out0;
assign v$MUX4_3087_out0 = v$G5_18151_out0 ? v$_9234_out0 : v$MUX5_4219_out0;
assign v$Y_8077_out0 = v$MUX1_15300_out0;
assign v$Y_8078_out0 = v$MUX1_15301_out0;
assign v$Y_8082_out0 = v$MUX1_15305_out0;
assign v$Y_8083_out0 = v$MUX1_15306_out0;
assign v$_10474_out0 = v$_17622_out0[2:0];
assign v$_10474_out1 = v$_17622_out0[5:3];
assign v$_10477_out0 = v$_17625_out0[2:0];
assign v$_10477_out1 = v$_17625_out0[5:3];
assign v$_14355_out0 = v$_16723_out0[2:0];
assign v$_14355_out1 = v$_16723_out0[5:3];
assign v$_14358_out0 = v$_16726_out0[2:0];
assign v$_14358_out1 = v$_16726_out0[5:3];
assign v$_19027_out0 = v$_16723_out1[2:0];
assign v$_19027_out1 = v$_16723_out1[5:3];
assign v$_19030_out0 = v$_16726_out1[2:0];
assign v$_19030_out1 = v$_16726_out1[5:3];
assign v$_1462_out0 = v$_19027_out0[0:0];
assign v$_1462_out1 = v$_19027_out0[2:2];
assign v$_1465_out0 = v$_19030_out0[0:0];
assign v$_1465_out1 = v$_19030_out0[2:2];
assign v$_1515_out0 = v$_14355_out1[0:0];
assign v$_1515_out1 = v$_14355_out1[2:2];
assign v$_1518_out0 = v$_14358_out1[0:0];
assign v$_1518_out1 = v$_14358_out1[2:2];
assign v$_2014_out0 = v$_2024_out1[0:0];
assign v$_2014_out1 = v$_2024_out1[2:2];
assign v$_2017_out0 = v$_2027_out1[0:0];
assign v$_2017_out1 = v$_2027_out1[2:2];
assign v$MUX14_5134_out0 = v$EQ14_5642_out0 ? v$SEL14_16964_out0 : v$MUX15_1479_out0;
assign v$MUX14_5135_out0 = v$EQ14_5643_out0 ? v$SEL14_16965_out0 : v$MUX15_1480_out0;
assign v$MUX14_5136_out0 = v$EQ14_5644_out0 ? v$SEL14_16966_out0 : v$MUX15_1481_out0;
assign v$MUX14_5137_out0 = v$EQ14_5645_out0 ? v$SEL14_16967_out0 : v$MUX15_1482_out0;
assign v$Z2_6574_out0 = v$Z_2748_out0;
assign v$Z2_6576_out0 = v$Z_2750_out0;
assign v$Z2_6578_out0 = v$Z_2752_out0;
assign v$Z2_6580_out0 = v$Z_2754_out0;
assign v$_7355_out0 = v$_14355_out0[0:0];
assign v$_7355_out1 = v$_14355_out0[2:2];
assign v$_7358_out0 = v$_14358_out0[0:0];
assign v$_7358_out1 = v$_14358_out0[2:2];
assign v$_9129_out0 = { v$Y_8077_out0,v$C6_6771_out0 };
assign v$_9131_out0 = { v$Y_8078_out0,v$C6_6773_out0 };
assign v$_9133_out0 = { v$Y_8082_out0,v$C6_6775_out0 };
assign v$_9135_out0 = { v$Y_8083_out0,v$C6_6777_out0 };
assign v$_10898_out0 = v$_10474_out0[0:0];
assign v$_10898_out1 = v$_10474_out0[2:2];
assign v$_10901_out0 = v$_10477_out0[0:0];
assign v$_10901_out1 = v$_10477_out0[2:2];
assign v$_11413_out0 = v$_19027_out1[0:0];
assign v$_11413_out1 = v$_19027_out1[2:2];
assign v$_11416_out0 = v$_19030_out1[0:0];
assign v$_11416_out1 = v$_19030_out1[2:2];
assign v$_11596_out0 = v$_2024_out0[0:0];
assign v$_11596_out1 = v$_2024_out0[2:2];
assign v$_11599_out0 = v$_2027_out0[0:0];
assign v$_11599_out1 = v$_2027_out0[2:2];
assign v$_16742_out0 = v$_10474_out1[0:0];
assign v$_16742_out1 = v$_10474_out1[2:2];
assign v$_16745_out0 = v$_10477_out1[0:0];
assign v$_16745_out1 = v$_10477_out1[2:2];
assign v$MUX3_18114_out0 = v$G4_6334_out0 ? v$_4136_out0 : v$MUX4_3084_out0;
assign v$MUX3_18115_out0 = v$G4_6335_out0 ? v$_4137_out0 : v$MUX4_3085_out0;
assign v$MUX3_18116_out0 = v$G4_6336_out0 ? v$_4138_out0 : v$MUX4_3086_out0;
assign v$MUX3_18117_out0 = v$G4_6337_out0 ? v$_4139_out0 : v$MUX4_3087_out0;
assign v$A6_320_out0 = v$_1462_out0;
assign v$A6_323_out0 = v$_1465_out0;
assign v$A21_2792_out0 = v$_2014_out0;
assign v$A21_2795_out0 = v$_2017_out0;
assign v$A12_3355_out0 = v$_10898_out0;
assign v$A12_3358_out0 = v$_10901_out0;
assign v$A9_3643_out0 = v$_11413_out0;
assign v$A9_3646_out0 = v$_11416_out0;
assign v$A0_4468_out0 = v$_7355_out0;
assign v$A0_4471_out0 = v$_7358_out0;
assign v$_6228_out0 = v$_16742_out1[0:0];
assign v$_6228_out1 = v$_16742_out1[1:1];
assign v$_6231_out0 = v$_16745_out1[0:0];
assign v$_6231_out1 = v$_16745_out1[1:1];
assign v$G6_6434_out0 = ! v$Z2_6574_out0;
assign v$G6_6436_out0 = ! v$Z2_6576_out0;
assign v$G6_6438_out0 = ! v$Z2_6578_out0;
assign v$G6_6440_out0 = ! v$Z2_6580_out0;
assign v$_7676_out0 = v$_1515_out1[0:0];
assign v$_7676_out1 = v$_1515_out1[1:1];
assign v$_7679_out0 = v$_1518_out1[0:0];
assign v$_7679_out1 = v$_1518_out1[1:1];
assign v$OUT_9282_out0 = v$MUX3_18114_out0;
assign v$OUT_9284_out0 = v$MUX3_18115_out0;
assign v$OUT_9286_out0 = v$MUX3_18116_out0;
assign v$OUT_9288_out0 = v$MUX3_18117_out0;
assign v$_10739_out0 = v$_2014_out1[0:0];
assign v$_10739_out1 = v$_2014_out1[1:1];
assign v$_10742_out0 = v$_2017_out1[0:0];
assign v$_10742_out1 = v$_2017_out1[1:1];
assign v$_12178_out0 = v$_7355_out1[0:0];
assign v$_12178_out1 = v$_7355_out1[1:1];
assign v$_12181_out0 = v$_7358_out1[0:0];
assign v$_12181_out1 = v$_7358_out1[1:1];
assign v$MUX13_14263_out0 = v$EQ13_9893_out0 ? v$SEL13_7205_out0 : v$MUX14_5134_out0;
assign v$MUX13_14264_out0 = v$EQ13_9894_out0 ? v$SEL13_7206_out0 : v$MUX14_5135_out0;
assign v$MUX13_14265_out0 = v$EQ13_9895_out0 ? v$SEL13_7207_out0 : v$MUX14_5136_out0;
assign v$MUX13_14266_out0 = v$EQ13_9896_out0 ? v$SEL13_7208_out0 : v$MUX14_5137_out0;
assign v$A3_15209_out0 = v$_1515_out0;
assign v$A3_15212_out0 = v$_1518_out0;
assign v$G9_15797_out0 = v$Z1_17592_out0 && v$Z2_6574_out0;
assign v$G9_15799_out0 = v$Z1_17594_out0 && v$Z2_6576_out0;
assign v$G9_15801_out0 = v$Z1_17596_out0 && v$Z2_6578_out0;
assign v$G9_15803_out0 = v$Z1_17598_out0 && v$Z2_6580_out0;
assign v$_16339_out0 = v$_1462_out1[0:0];
assign v$_16339_out1 = v$_1462_out1[1:1];
assign v$_16342_out0 = v$_1465_out1[0:0];
assign v$_16342_out1 = v$_1465_out1[1:1];
assign v$_16791_out0 = v$_10898_out1[0:0];
assign v$_16791_out1 = v$_10898_out1[1:1];
assign v$_16794_out0 = v$_10901_out1[0:0];
assign v$_16794_out1 = v$_10901_out1[1:1];
assign v$_17322_out0 = v$_11596_out1[0:0];
assign v$_17322_out1 = v$_11596_out1[1:1];
assign v$_17325_out0 = v$_11599_out1[0:0];
assign v$_17325_out1 = v$_11599_out1[1:1];
assign v$A15_17957_out0 = v$_16742_out0;
assign v$A15_17960_out0 = v$_16745_out0;
assign v$A18_18300_out0 = v$_11596_out0;
assign v$A18_18303_out0 = v$_11599_out0;
assign v$_18366_out0 = v$_11413_out1[0:0];
assign v$_18366_out1 = v$_11413_out1[1:1];
assign v$_18369_out0 = v$_11416_out1[0:0];
assign v$_18369_out1 = v$_11416_out1[1:1];
assign v$A14_738_out0 = v$_16791_out1;
assign v$A14_741_out0 = v$_16794_out1;
assign v$A19_1363_out0 = v$_17322_out0;
assign v$A19_1366_out0 = v$_17325_out0;
assign v$A10_1703_out0 = v$_18366_out0;
assign v$A10_1706_out0 = v$_18369_out0;
assign v$A1_1869_out0 = v$_12178_out0;
assign v$A1_1872_out0 = v$_12181_out0;
assign v$Z_2747_out0 = v$G9_15797_out0;
assign v$Z_2749_out0 = v$G9_15799_out0;
assign v$Z_2751_out0 = v$G9_15801_out0;
assign v$Z_2753_out0 = v$G9_15803_out0;
assign v$A22_4590_out0 = v$_10739_out0;
assign v$A22_4593_out0 = v$_10742_out0;
assign v$A20_4603_out0 = v$_17322_out1;
assign v$A20_4606_out0 = v$_17325_out1;
assign v$A23_5281_out0 = v$_10739_out1;
assign v$A23_5284_out0 = v$_10742_out1;
assign v$_5309_out0 = { v$OUT_9282_out0,v$C5_17519_out0 };
assign v$_5311_out0 = { v$OUT_9284_out0,v$C5_17521_out0 };
assign v$_5313_out0 = { v$OUT_9286_out0,v$C5_17523_out0 };
assign v$_5315_out0 = { v$OUT_9288_out0,v$C5_17525_out0 };
assign v$A5_6901_out0 = v$_7676_out1;
assign v$A5_6904_out0 = v$_7679_out1;
assign v$A_7391_out0 = v$A6_320_out0;
assign v$A_7392_out0 = v$A3_15209_out0;
assign v$A_7393_out0 = v$A21_2792_out0;
assign v$A_7394_out0 = v$A9_3643_out0;
assign v$A_7395_out0 = v$A15_17957_out0;
assign v$A_7399_out0 = v$A12_3355_out0;
assign v$A_7403_out0 = v$A0_4468_out0;
assign v$A_7408_out0 = v$A18_18300_out0;
assign v$A_7463_out0 = v$A6_323_out0;
assign v$A_7464_out0 = v$A3_15212_out0;
assign v$A_7465_out0 = v$A21_2795_out0;
assign v$A_7466_out0 = v$A9_3646_out0;
assign v$A_7467_out0 = v$A15_17960_out0;
assign v$A_7471_out0 = v$A12_3358_out0;
assign v$A_7475_out0 = v$A0_4471_out0;
assign v$A_7480_out0 = v$A18_18303_out0;
assign v$A11_10386_out0 = v$_18366_out1;
assign v$A11_10389_out0 = v$_18369_out1;
assign {v$A1A_12224_out1,v$A1A_12224_out0 } = v$A0_4468_out0 + v$B0_3421_out0 + v$C1_4633_out0;
assign {v$A1A_12227_out1,v$A1A_12227_out0 } = v$A0_4471_out0 + v$B0_3424_out0 + v$C1_4636_out0;
assign v$A16_14191_out0 = v$_6228_out0;
assign v$A16_14194_out0 = v$_6231_out0;
assign v$A13_14445_out0 = v$_16791_out0;
assign v$A13_14448_out0 = v$_16794_out0;
assign v$A7_15891_out0 = v$_16339_out0;
assign v$A7_15894_out0 = v$_16342_out0;
assign v$A17_17342_out0 = v$_6228_out1;
assign v$A17_17345_out0 = v$_6231_out1;
assign v$A4_18138_out0 = v$_7676_out0;
assign v$A4_18141_out0 = v$_7679_out0;
assign v$MUX12_18419_out0 = v$EQ12_14427_out0 ? v$SEL12_14433_out0 : v$MUX13_14263_out0;
assign v$MUX12_18420_out0 = v$EQ12_14428_out0 ? v$SEL12_14434_out0 : v$MUX13_14264_out0;
assign v$MUX12_18421_out0 = v$EQ12_14429_out0 ? v$SEL12_14435_out0 : v$MUX13_14265_out0;
assign v$MUX12_18422_out0 = v$EQ12_14430_out0 ? v$SEL12_14436_out0 : v$MUX13_14266_out0;
assign v$A8_18697_out0 = v$_16339_out1;
assign v$A8_18700_out0 = v$_16342_out1;
assign v$A2_18868_out0 = v$_12178_out1;
assign v$A2_18871_out0 = v$_12181_out1;
assign v$MUX5_4212_out0 = v$G6_6434_out0 ? v$_5309_out0 : v$_9129_out0;
assign v$MUX5_4214_out0 = v$G6_6436_out0 ? v$_5311_out0 : v$_9131_out0;
assign v$MUX5_4216_out0 = v$G6_6438_out0 ? v$_5313_out0 : v$_9133_out0;
assign v$MUX5_4218_out0 = v$G6_6440_out0 ? v$_5315_out0 : v$_9135_out0;
assign v$G2_5478_out0 = ((v$A_7391_out0 && !v$B_2896_out0) || (!v$A_7391_out0) && v$B_2896_out0);
assign v$G2_5479_out0 = ((v$A_7392_out0 && !v$B_2897_out0) || (!v$A_7392_out0) && v$B_2897_out0);
assign v$G2_5480_out0 = ((v$A_7393_out0 && !v$B_2898_out0) || (!v$A_7393_out0) && v$B_2898_out0);
assign v$G2_5481_out0 = ((v$A_7394_out0 && !v$B_2899_out0) || (!v$A_7394_out0) && v$B_2899_out0);
assign v$G2_5482_out0 = ((v$A_7395_out0 && !v$B_2900_out0) || (!v$A_7395_out0) && v$B_2900_out0);
assign v$G2_5486_out0 = ((v$A_7399_out0 && !v$B_2904_out0) || (!v$A_7399_out0) && v$B_2904_out0);
assign v$G2_5490_out0 = ((v$A_7403_out0 && !v$B_2908_out0) || (!v$A_7403_out0) && v$B_2908_out0);
assign v$G2_5495_out0 = ((v$A_7408_out0 && !v$B_2913_out0) || (!v$A_7408_out0) && v$B_2913_out0);
assign v$G2_5550_out0 = ((v$A_7463_out0 && !v$B_2968_out0) || (!v$A_7463_out0) && v$B_2968_out0);
assign v$G2_5551_out0 = ((v$A_7464_out0 && !v$B_2969_out0) || (!v$A_7464_out0) && v$B_2969_out0);
assign v$G2_5552_out0 = ((v$A_7465_out0 && !v$B_2970_out0) || (!v$A_7465_out0) && v$B_2970_out0);
assign v$G2_5553_out0 = ((v$A_7466_out0 && !v$B_2971_out0) || (!v$A_7466_out0) && v$B_2971_out0);
assign v$G2_5554_out0 = ((v$A_7467_out0 && !v$B_2972_out0) || (!v$A_7467_out0) && v$B_2972_out0);
assign v$G2_5558_out0 = ((v$A_7471_out0 && !v$B_2976_out0) || (!v$A_7471_out0) && v$B_2976_out0);
assign v$G2_5562_out0 = ((v$A_7475_out0 && !v$B_2980_out0) || (!v$A_7475_out0) && v$B_2980_out0);
assign v$G2_5567_out0 = ((v$A_7480_out0 && !v$B_2985_out0) || (!v$A_7480_out0) && v$B_2985_out0);
assign v$A_7396_out0 = v$A7_15891_out0;
assign v$A_7397_out0 = v$A1_1869_out0;
assign v$A_7398_out0 = v$A14_738_out0;
assign v$A_7400_out0 = v$A8_18697_out0;
assign v$A_7401_out0 = v$A17_17342_out0;
assign v$A_7402_out0 = v$A23_5281_out0;
assign v$A_7404_out0 = v$A13_14445_out0;
assign v$A_7405_out0 = v$A4_18138_out0;
assign v$A_7406_out0 = v$A19_1363_out0;
assign v$A_7407_out0 = v$A22_4590_out0;
assign v$A_7409_out0 = v$A10_1703_out0;
assign v$A_7410_out0 = v$A20_4603_out0;
assign v$A_7411_out0 = v$A2_18868_out0;
assign v$A_7412_out0 = v$A11_10386_out0;
assign v$A_7413_out0 = v$A5_6901_out0;
assign v$A_7414_out0 = v$A16_14191_out0;
assign v$A_7468_out0 = v$A7_15894_out0;
assign v$A_7469_out0 = v$A1_1872_out0;
assign v$A_7470_out0 = v$A14_741_out0;
assign v$A_7472_out0 = v$A8_18700_out0;
assign v$A_7473_out0 = v$A17_17345_out0;
assign v$A_7474_out0 = v$A23_5284_out0;
assign v$A_7476_out0 = v$A13_14448_out0;
assign v$A_7477_out0 = v$A4_18141_out0;
assign v$A_7478_out0 = v$A19_1366_out0;
assign v$A_7479_out0 = v$A22_4593_out0;
assign v$A_7481_out0 = v$A10_1706_out0;
assign v$A_7482_out0 = v$A20_4606_out0;
assign v$A_7483_out0 = v$A2_18871_out0;
assign v$A_7484_out0 = v$A11_10389_out0;
assign v$A_7485_out0 = v$A5_6904_out0;
assign v$A_7486_out0 = v$A16_14194_out0;
assign v$G1_12902_out0 = v$A_7391_out0 && v$B_2896_out0;
assign v$G1_12903_out0 = v$A_7392_out0 && v$B_2897_out0;
assign v$G1_12904_out0 = v$A_7393_out0 && v$B_2898_out0;
assign v$G1_12905_out0 = v$A_7394_out0 && v$B_2899_out0;
assign v$G1_12906_out0 = v$A_7395_out0 && v$B_2900_out0;
assign v$G1_12910_out0 = v$A_7399_out0 && v$B_2904_out0;
assign v$G1_12914_out0 = v$A_7403_out0 && v$B_2908_out0;
assign v$G1_12919_out0 = v$A_7408_out0 && v$B_2913_out0;
assign v$G1_12974_out0 = v$A_7463_out0 && v$B_2968_out0;
assign v$G1_12975_out0 = v$A_7464_out0 && v$B_2969_out0;
assign v$G1_12976_out0 = v$A_7465_out0 && v$B_2970_out0;
assign v$G1_12977_out0 = v$A_7466_out0 && v$B_2971_out0;
assign v$G1_12978_out0 = v$A_7467_out0 && v$B_2972_out0;
assign v$G1_12982_out0 = v$A_7471_out0 && v$B_2976_out0;
assign v$G1_12986_out0 = v$A_7475_out0 && v$B_2980_out0;
assign v$G1_12991_out0 = v$A_7480_out0 && v$B_2985_out0;
assign v$Z_16411_out0 = v$Z_2747_out0;
assign v$Z_16412_out0 = v$Z_2749_out0;
assign v$Z_16413_out0 = v$Z_2751_out0;
assign v$Z_16414_out0 = v$Z_2753_out0;
assign v$MUX11_18547_out0 = v$EQ11_6408_out0 ? v$SEL11_7539_out0 : v$MUX12_18419_out0;
assign v$MUX11_18548_out0 = v$EQ11_6409_out0 ? v$SEL11_7540_out0 : v$MUX12_18420_out0;
assign v$MUX11_18549_out0 = v$EQ11_6410_out0 ? v$SEL11_7541_out0 : v$MUX12_18421_out0;
assign v$MUX11_18550_out0 = v$EQ11_6411_out0 ? v$SEL11_7542_out0 : v$MUX12_18422_out0;
assign v$END_18875_out0 = v$A1A_12224_out1;
assign v$END_18878_out0 = v$A1A_12227_out1;
assign v$MUX8_3154_out0 = v$EQ9_14361_out0 ? v$SEL9_10717_out0 : v$MUX11_18547_out0;
assign v$MUX8_3155_out0 = v$EQ9_14362_out0 ? v$SEL9_10718_out0 : v$MUX11_18548_out0;
assign v$MUX8_3156_out0 = v$EQ9_14363_out0 ? v$SEL9_10719_out0 : v$MUX11_18549_out0;
assign v$MUX8_3157_out0 = v$EQ9_14364_out0 ? v$SEL9_10720_out0 : v$MUX11_18550_out0;
assign v$G2_5483_out0 = ((v$A_7396_out0 && !v$B_2901_out0) || (!v$A_7396_out0) && v$B_2901_out0);
assign v$G2_5484_out0 = ((v$A_7397_out0 && !v$B_2902_out0) || (!v$A_7397_out0) && v$B_2902_out0);
assign v$G2_5485_out0 = ((v$A_7398_out0 && !v$B_2903_out0) || (!v$A_7398_out0) && v$B_2903_out0);
assign v$G2_5487_out0 = ((v$A_7400_out0 && !v$B_2905_out0) || (!v$A_7400_out0) && v$B_2905_out0);
assign v$G2_5488_out0 = ((v$A_7401_out0 && !v$B_2906_out0) || (!v$A_7401_out0) && v$B_2906_out0);
assign v$G2_5489_out0 = ((v$A_7402_out0 && !v$B_2907_out0) || (!v$A_7402_out0) && v$B_2907_out0);
assign v$G2_5491_out0 = ((v$A_7404_out0 && !v$B_2909_out0) || (!v$A_7404_out0) && v$B_2909_out0);
assign v$G2_5492_out0 = ((v$A_7405_out0 && !v$B_2910_out0) || (!v$A_7405_out0) && v$B_2910_out0);
assign v$G2_5493_out0 = ((v$A_7406_out0 && !v$B_2911_out0) || (!v$A_7406_out0) && v$B_2911_out0);
assign v$G2_5494_out0 = ((v$A_7407_out0 && !v$B_2912_out0) || (!v$A_7407_out0) && v$B_2912_out0);
assign v$G2_5496_out0 = ((v$A_7409_out0 && !v$B_2914_out0) || (!v$A_7409_out0) && v$B_2914_out0);
assign v$G2_5497_out0 = ((v$A_7410_out0 && !v$B_2915_out0) || (!v$A_7410_out0) && v$B_2915_out0);
assign v$G2_5498_out0 = ((v$A_7411_out0 && !v$B_2916_out0) || (!v$A_7411_out0) && v$B_2916_out0);
assign v$G2_5499_out0 = ((v$A_7412_out0 && !v$B_2917_out0) || (!v$A_7412_out0) && v$B_2917_out0);
assign v$G2_5500_out0 = ((v$A_7413_out0 && !v$B_2918_out0) || (!v$A_7413_out0) && v$B_2918_out0);
assign v$G2_5501_out0 = ((v$A_7414_out0 && !v$B_2919_out0) || (!v$A_7414_out0) && v$B_2919_out0);
assign v$G2_5555_out0 = ((v$A_7468_out0 && !v$B_2973_out0) || (!v$A_7468_out0) && v$B_2973_out0);
assign v$G2_5556_out0 = ((v$A_7469_out0 && !v$B_2974_out0) || (!v$A_7469_out0) && v$B_2974_out0);
assign v$G2_5557_out0 = ((v$A_7470_out0 && !v$B_2975_out0) || (!v$A_7470_out0) && v$B_2975_out0);
assign v$G2_5559_out0 = ((v$A_7472_out0 && !v$B_2977_out0) || (!v$A_7472_out0) && v$B_2977_out0);
assign v$G2_5560_out0 = ((v$A_7473_out0 && !v$B_2978_out0) || (!v$A_7473_out0) && v$B_2978_out0);
assign v$G2_5561_out0 = ((v$A_7474_out0 && !v$B_2979_out0) || (!v$A_7474_out0) && v$B_2979_out0);
assign v$G2_5563_out0 = ((v$A_7476_out0 && !v$B_2981_out0) || (!v$A_7476_out0) && v$B_2981_out0);
assign v$G2_5564_out0 = ((v$A_7477_out0 && !v$B_2982_out0) || (!v$A_7477_out0) && v$B_2982_out0);
assign v$G2_5565_out0 = ((v$A_7478_out0 && !v$B_2983_out0) || (!v$A_7478_out0) && v$B_2983_out0);
assign v$G2_5566_out0 = ((v$A_7479_out0 && !v$B_2984_out0) || (!v$A_7479_out0) && v$B_2984_out0);
assign v$G2_5568_out0 = ((v$A_7481_out0 && !v$B_2986_out0) || (!v$A_7481_out0) && v$B_2986_out0);
assign v$G2_5569_out0 = ((v$A_7482_out0 && !v$B_2987_out0) || (!v$A_7482_out0) && v$B_2987_out0);
assign v$G2_5570_out0 = ((v$A_7483_out0 && !v$B_2988_out0) || (!v$A_7483_out0) && v$B_2988_out0);
assign v$G2_5571_out0 = ((v$A_7484_out0 && !v$B_2989_out0) || (!v$A_7484_out0) && v$B_2989_out0);
assign v$G2_5572_out0 = ((v$A_7485_out0 && !v$B_2990_out0) || (!v$A_7485_out0) && v$B_2990_out0);
assign v$G2_5573_out0 = ((v$A_7486_out0 && !v$B_2991_out0) || (!v$A_7486_out0) && v$B_2991_out0);
assign v$OUT_9281_out0 = v$MUX5_4212_out0;
assign v$OUT_9283_out0 = v$MUX5_4214_out0;
assign v$OUT_9285_out0 = v$MUX5_4216_out0;
assign v$OUT_9287_out0 = v$MUX5_4218_out0;
assign v$G_10482_out0 = v$G1_12902_out0;
assign v$G_10483_out0 = v$G1_12903_out0;
assign v$G_10484_out0 = v$G1_12904_out0;
assign v$G_10485_out0 = v$G1_12905_out0;
assign v$G_10486_out0 = v$G1_12906_out0;
assign v$G_10490_out0 = v$G1_12910_out0;
assign v$G_10494_out0 = v$G1_12914_out0;
assign v$G_10499_out0 = v$G1_12919_out0;
assign v$G_10554_out0 = v$G1_12974_out0;
assign v$G_10555_out0 = v$G1_12975_out0;
assign v$G_10556_out0 = v$G1_12976_out0;
assign v$G_10557_out0 = v$G1_12977_out0;
assign v$G_10558_out0 = v$G1_12978_out0;
assign v$G_10562_out0 = v$G1_12982_out0;
assign v$G_10566_out0 = v$G1_12986_out0;
assign v$G_10571_out0 = v$G1_12991_out0;
assign v$G1_12907_out0 = v$A_7396_out0 && v$B_2901_out0;
assign v$G1_12908_out0 = v$A_7397_out0 && v$B_2902_out0;
assign v$G1_12909_out0 = v$A_7398_out0 && v$B_2903_out0;
assign v$G1_12911_out0 = v$A_7400_out0 && v$B_2905_out0;
assign v$G1_12912_out0 = v$A_7401_out0 && v$B_2906_out0;
assign v$G1_12913_out0 = v$A_7402_out0 && v$B_2907_out0;
assign v$G1_12915_out0 = v$A_7404_out0 && v$B_2909_out0;
assign v$G1_12916_out0 = v$A_7405_out0 && v$B_2910_out0;
assign v$G1_12917_out0 = v$A_7406_out0 && v$B_2911_out0;
assign v$G1_12918_out0 = v$A_7407_out0 && v$B_2912_out0;
assign v$G1_12920_out0 = v$A_7409_out0 && v$B_2914_out0;
assign v$G1_12921_out0 = v$A_7410_out0 && v$B_2915_out0;
assign v$G1_12922_out0 = v$A_7411_out0 && v$B_2916_out0;
assign v$G1_12923_out0 = v$A_7412_out0 && v$B_2917_out0;
assign v$G1_12924_out0 = v$A_7413_out0 && v$B_2918_out0;
assign v$G1_12925_out0 = v$A_7414_out0 && v$B_2919_out0;
assign v$G1_12979_out0 = v$A_7468_out0 && v$B_2973_out0;
assign v$G1_12980_out0 = v$A_7469_out0 && v$B_2974_out0;
assign v$G1_12981_out0 = v$A_7470_out0 && v$B_2975_out0;
assign v$G1_12983_out0 = v$A_7472_out0 && v$B_2977_out0;
assign v$G1_12984_out0 = v$A_7473_out0 && v$B_2978_out0;
assign v$G1_12985_out0 = v$A_7474_out0 && v$B_2979_out0;
assign v$G1_12987_out0 = v$A_7476_out0 && v$B_2981_out0;
assign v$G1_12988_out0 = v$A_7477_out0 && v$B_2982_out0;
assign v$G1_12989_out0 = v$A_7478_out0 && v$B_2983_out0;
assign v$G1_12990_out0 = v$A_7479_out0 && v$B_2984_out0;
assign v$G1_12992_out0 = v$A_7481_out0 && v$B_2986_out0;
assign v$G1_12993_out0 = v$A_7482_out0 && v$B_2987_out0;
assign v$G1_12994_out0 = v$A_7483_out0 && v$B_2988_out0;
assign v$G1_12995_out0 = v$A_7484_out0 && v$B_2989_out0;
assign v$G1_12996_out0 = v$A_7485_out0 && v$B_2990_out0;
assign v$G1_12997_out0 = v$A_7486_out0 && v$B_2991_out0;
assign v$P_14453_out0 = v$G2_5478_out0;
assign v$P_14454_out0 = v$G2_5479_out0;
assign v$P_14455_out0 = v$G2_5480_out0;
assign v$P_14456_out0 = v$G2_5481_out0;
assign v$P_14457_out0 = v$G2_5482_out0;
assign v$P_14461_out0 = v$G2_5486_out0;
assign v$P_14465_out0 = v$G2_5490_out0;
assign v$P_14470_out0 = v$G2_5495_out0;
assign v$P_14525_out0 = v$G2_5550_out0;
assign v$P_14526_out0 = v$G2_5551_out0;
assign v$P_14527_out0 = v$G2_5552_out0;
assign v$P_14528_out0 = v$G2_5553_out0;
assign v$P_14529_out0 = v$G2_5554_out0;
assign v$P_14533_out0 = v$G2_5558_out0;
assign v$P_14537_out0 = v$G2_5562_out0;
assign v$P_14542_out0 = v$G2_5567_out0;
assign v$P12_243_out0 = v$P_14461_out0;
assign v$P12_246_out0 = v$P_14533_out0;
assign v$P21_4981_out0 = v$P_14455_out0;
assign v$P21_4984_out0 = v$P_14527_out0;
assign v$P0_5023_out0 = v$P_14465_out0;
assign v$P0_5026_out0 = v$P_14537_out0;
assign v$P15_7183_out0 = v$P_14457_out0;
assign v$P15_7186_out0 = v$P_14529_out0;
assign v$G12_7327_out0 = v$G_10490_out0;
assign v$G12_7330_out0 = v$G_10562_out0;
assign v$P6_8418_out0 = v$P_14453_out0;
assign v$P6_8421_out0 = v$P_14525_out0;
assign v$G9_9255_out0 = v$G_10485_out0;
assign v$G9_9258_out0 = v$G_10557_out0;
assign v$AMOUNT$OF$SHIFT_9833_out0 = v$OUT_9281_out0;
assign v$AMOUNT$OF$SHIFT_9834_out0 = v$OUT_9283_out0;
assign v$AMOUNT$OF$SHIFT_9835_out0 = v$OUT_9285_out0;
assign v$AMOUNT$OF$SHIFT_9836_out0 = v$OUT_9287_out0;
assign v$G_10487_out0 = v$G1_12907_out0;
assign v$G_10488_out0 = v$G1_12908_out0;
assign v$G_10489_out0 = v$G1_12909_out0;
assign v$G_10491_out0 = v$G1_12911_out0;
assign v$G_10492_out0 = v$G1_12912_out0;
assign v$G_10493_out0 = v$G1_12913_out0;
assign v$G_10495_out0 = v$G1_12915_out0;
assign v$G_10496_out0 = v$G1_12916_out0;
assign v$G_10497_out0 = v$G1_12917_out0;
assign v$G_10498_out0 = v$G1_12918_out0;
assign v$G_10500_out0 = v$G1_12920_out0;
assign v$G_10501_out0 = v$G1_12921_out0;
assign v$G_10502_out0 = v$G1_12922_out0;
assign v$G_10503_out0 = v$G1_12923_out0;
assign v$G_10504_out0 = v$G1_12924_out0;
assign v$G_10505_out0 = v$G1_12925_out0;
assign v$G_10559_out0 = v$G1_12979_out0;
assign v$G_10560_out0 = v$G1_12980_out0;
assign v$G_10561_out0 = v$G1_12981_out0;
assign v$G_10563_out0 = v$G1_12983_out0;
assign v$G_10564_out0 = v$G1_12984_out0;
assign v$G_10565_out0 = v$G1_12985_out0;
assign v$G_10567_out0 = v$G1_12987_out0;
assign v$G_10568_out0 = v$G1_12988_out0;
assign v$G_10569_out0 = v$G1_12989_out0;
assign v$G_10570_out0 = v$G1_12990_out0;
assign v$G_10572_out0 = v$G1_12992_out0;
assign v$G_10573_out0 = v$G1_12993_out0;
assign v$G_10574_out0 = v$G1_12994_out0;
assign v$G_10575_out0 = v$G1_12995_out0;
assign v$G_10576_out0 = v$G1_12996_out0;
assign v$G_10577_out0 = v$G1_12997_out0;
assign v$G15_11541_out0 = v$G_10486_out0;
assign v$G15_11544_out0 = v$G_10558_out0;
assign v$G3_11602_out0 = v$G_10483_out0;
assign v$G3_11605_out0 = v$G_10555_out0;
assign v$P18_12290_out0 = v$P_14470_out0;
assign v$P18_12293_out0 = v$P_14542_out0;
assign v$G18_13508_out0 = v$G_10499_out0;
assign v$G18_13511_out0 = v$G_10571_out0;
assign v$P_14458_out0 = v$G2_5483_out0;
assign v$P_14459_out0 = v$G2_5484_out0;
assign v$P_14460_out0 = v$G2_5485_out0;
assign v$P_14462_out0 = v$G2_5487_out0;
assign v$P_14463_out0 = v$G2_5488_out0;
assign v$P_14464_out0 = v$G2_5489_out0;
assign v$P_14466_out0 = v$G2_5491_out0;
assign v$P_14467_out0 = v$G2_5492_out0;
assign v$P_14468_out0 = v$G2_5493_out0;
assign v$P_14469_out0 = v$G2_5494_out0;
assign v$P_14471_out0 = v$G2_5496_out0;
assign v$P_14472_out0 = v$G2_5497_out0;
assign v$P_14473_out0 = v$G2_5498_out0;
assign v$P_14474_out0 = v$G2_5499_out0;
assign v$P_14475_out0 = v$G2_5500_out0;
assign v$P_14476_out0 = v$G2_5501_out0;
assign v$P_14530_out0 = v$G2_5555_out0;
assign v$P_14531_out0 = v$G2_5556_out0;
assign v$P_14532_out0 = v$G2_5557_out0;
assign v$P_14534_out0 = v$G2_5559_out0;
assign v$P_14535_out0 = v$G2_5560_out0;
assign v$P_14536_out0 = v$G2_5561_out0;
assign v$P_14538_out0 = v$G2_5563_out0;
assign v$P_14539_out0 = v$G2_5564_out0;
assign v$P_14540_out0 = v$G2_5565_out0;
assign v$P_14541_out0 = v$G2_5566_out0;
assign v$P_14543_out0 = v$G2_5568_out0;
assign v$P_14544_out0 = v$G2_5569_out0;
assign v$P_14545_out0 = v$G2_5570_out0;
assign v$P_14546_out0 = v$G2_5571_out0;
assign v$P_14547_out0 = v$G2_5572_out0;
assign v$P_14548_out0 = v$G2_5573_out0;
assign v$G21_14626_out0 = v$G_10484_out0;
assign v$G21_14629_out0 = v$G_10556_out0;
assign v$P3_15921_out0 = v$P_14454_out0;
assign v$P3_15924_out0 = v$P_14526_out0;
assign v$MUX10_16266_out0 = v$EQ10_6169_out0 ? v$SEL8_18285_out0 : v$MUX8_3154_out0;
assign v$MUX10_16267_out0 = v$EQ10_6170_out0 ? v$SEL8_18286_out0 : v$MUX8_3155_out0;
assign v$MUX10_16268_out0 = v$EQ10_6171_out0 ? v$SEL8_18287_out0 : v$MUX8_3156_out0;
assign v$MUX10_16269_out0 = v$EQ10_6172_out0 ? v$SEL8_18288_out0 : v$MUX8_3157_out0;
assign v$G0_16548_out0 = v$G_10494_out0;
assign v$G0_16551_out0 = v$G_10566_out0;
assign v$G6_16970_out0 = v$G_10482_out0;
assign v$G6_16973_out0 = v$G_10554_out0;
assign v$P9_19053_out0 = v$P_14456_out0;
assign v$P9_19056_out0 = v$P_14528_out0;
assign v$P5_228_out0 = v$P_14475_out0;
assign v$P5_231_out0 = v$P_14547_out0;
assign v$P10_360_out0 = v$P_14471_out0;
assign v$P10_363_out0 = v$P_14543_out0;
assign v$G$CD_1027_out0 = v$G6_16970_out0;
assign v$G$CD_1028_out0 = v$G3_11602_out0;
assign v$G$CD_1029_out0 = v$G12_7327_out0;
assign v$G$CD_1030_out0 = v$G9_9255_out0;
assign v$G$CD_1033_out0 = v$G18_13508_out0;
assign v$G$CD_1044_out0 = v$G15_11541_out0;
assign v$G$CD_1045_out0 = v$G21_14626_out0;
assign v$G$CD_1150_out0 = v$G6_16973_out0;
assign v$G$CD_1151_out0 = v$G3_11605_out0;
assign v$G$CD_1152_out0 = v$G12_7330_out0;
assign v$G$CD_1153_out0 = v$G9_9258_out0;
assign v$G$CD_1156_out0 = v$G18_13511_out0;
assign v$G$CD_1167_out0 = v$G15_11544_out0;
assign v$G$CD_1168_out0 = v$G21_14629_out0;
assign v$G7_1849_out0 = v$G_10487_out0;
assign v$G7_1852_out0 = v$G_10559_out0;
assign v$P8_1861_out0 = v$P_14462_out0;
assign v$P8_1864_out0 = v$P_14534_out0;
assign v$G10_1993_out0 = v$G_10500_out0;
assign v$G10_1996_out0 = v$G_10572_out0;
assign v$SEL4_2005_out0 = v$AMOUNT$OF$SHIFT_9833_out0[3:3];
assign v$SEL4_2006_out0 = v$AMOUNT$OF$SHIFT_9834_out0[3:3];
assign v$SEL4_2007_out0 = v$AMOUNT$OF$SHIFT_9835_out0[3:3];
assign v$SEL4_2008_out0 = v$AMOUNT$OF$SHIFT_9836_out0[3:3];
assign v$G19_2044_out0 = v$G_10497_out0;
assign v$G19_2047_out0 = v$G_10569_out0;
assign v$P$AB_2168_out0 = v$P0_5023_out0;
assign v$P$AB_2171_out0 = v$P18_12290_out0;
assign v$P$AB_2172_out0 = v$P21_4981_out0;
assign v$P$AB_2184_out0 = v$P12_243_out0;
assign v$P$AB_2186_out0 = v$P15_7183_out0;
assign v$P$AB_2189_out0 = v$P6_8418_out0;
assign v$P$AB_2195_out0 = v$P3_15921_out0;
assign v$P$AB_2200_out0 = v$P9_19053_out0;
assign v$P$AB_2291_out0 = v$P0_5026_out0;
assign v$P$AB_2294_out0 = v$P18_12293_out0;
assign v$P$AB_2295_out0 = v$P21_4984_out0;
assign v$P$AB_2307_out0 = v$P12_246_out0;
assign v$P$AB_2309_out0 = v$P15_7186_out0;
assign v$P$AB_2312_out0 = v$P6_8421_out0;
assign v$P$AB_2318_out0 = v$P3_15924_out0;
assign v$P$AB_2323_out0 = v$P9_19056_out0;
assign v$P2_2424_out0 = v$P_14473_out0;
assign v$P2_2427_out0 = v$P_14545_out0;
assign v$G8_2770_out0 = v$G_10491_out0;
assign v$G8_2773_out0 = v$G_10563_out0;
assign v$G13_3052_out0 = v$G_10495_out0;
assign v$G13_3055_out0 = v$G_10567_out0;
assign v$P1_3168_out0 = v$P_14459_out0;
assign v$P1_3171_out0 = v$P_14531_out0;
assign v$P13_3245_out0 = v$P_14466_out0;
assign v$P13_3248_out0 = v$P_14538_out0;
assign v$P14_3369_out0 = v$P_14460_out0;
assign v$P14_3372_out0 = v$P_14532_out0;
assign v$P22_4945_out0 = v$P_14469_out0;
assign v$P22_4948_out0 = v$P_14541_out0;
assign v$G1_5269_out0 = v$G_10488_out0;
assign v$G1_5272_out0 = v$G_10560_out0;
assign v$G4_6019_out0 = v$G_10496_out0;
assign v$G4_6022_out0 = v$G_10568_out0;
assign v$P23_6626_out0 = v$P_14464_out0;
assign v$P23_6629_out0 = v$P_14536_out0;
assign v$P16_7243_out0 = v$P_14476_out0;
assign v$P16_7246_out0 = v$P_14548_out0;
assign v$G20_8533_out0 = v$G_10501_out0;
assign v$G20_8536_out0 = v$G_10573_out0;
assign v$MUX9_8553_out0 = v$EQ8_15018_out0 ? v$SEL10_9883_out0 : v$MUX10_16266_out0;
assign v$MUX9_8554_out0 = v$EQ8_15019_out0 ? v$SEL10_9884_out0 : v$MUX10_16267_out0;
assign v$MUX9_8555_out0 = v$EQ8_15020_out0 ? v$SEL10_9885_out0 : v$MUX10_16268_out0;
assign v$MUX9_8556_out0 = v$EQ8_15021_out0 ? v$SEL10_9886_out0 : v$MUX10_16269_out0;
assign v$G$AB_9468_out0 = v$G0_16548_out0;
assign v$G$AB_9471_out0 = v$G18_13508_out0;
assign v$G$AB_9472_out0 = v$G21_14626_out0;
assign v$G$AB_9484_out0 = v$G12_7327_out0;
assign v$G$AB_9486_out0 = v$G15_11541_out0;
assign v$G$AB_9489_out0 = v$G6_16970_out0;
assign v$G$AB_9495_out0 = v$G3_11602_out0;
assign v$G$AB_9500_out0 = v$G9_9255_out0;
assign v$G$AB_9591_out0 = v$G0_16551_out0;
assign v$G$AB_9594_out0 = v$G18_13511_out0;
assign v$G$AB_9595_out0 = v$G21_14629_out0;
assign v$G$AB_9607_out0 = v$G12_7330_out0;
assign v$G$AB_9609_out0 = v$G15_11544_out0;
assign v$G$AB_9612_out0 = v$G6_16973_out0;
assign v$G$AB_9618_out0 = v$G3_11605_out0;
assign v$G$AB_9623_out0 = v$G9_9258_out0;
assign v$G17_9714_out0 = v$G_10492_out0;
assign v$G17_9717_out0 = v$G_10564_out0;
assign v$P11_9992_out0 = v$P_14474_out0;
assign v$P11_9995_out0 = v$P_14546_out0;
assign v$P$CD_10916_out0 = v$P6_8418_out0;
assign v$P$CD_10917_out0 = v$P3_15921_out0;
assign v$P$CD_10918_out0 = v$P12_243_out0;
assign v$P$CD_10919_out0 = v$P9_19053_out0;
assign v$P$CD_10922_out0 = v$P18_12290_out0;
assign v$P$CD_10933_out0 = v$P15_7183_out0;
assign v$P$CD_10934_out0 = v$P21_4981_out0;
assign v$P$CD_11039_out0 = v$P6_8421_out0;
assign v$P$CD_11040_out0 = v$P3_15924_out0;
assign v$P$CD_11041_out0 = v$P12_246_out0;
assign v$P$CD_11042_out0 = v$P9_19056_out0;
assign v$P$CD_11045_out0 = v$P18_12293_out0;
assign v$P$CD_11056_out0 = v$P15_7186_out0;
assign v$P$CD_11057_out0 = v$P21_4984_out0;
assign v$P20_11152_out0 = v$P_14472_out0;
assign v$P20_11155_out0 = v$P_14544_out0;
assign v$G5_11170_out0 = v$G_10504_out0;
assign v$G5_11173_out0 = v$G_10576_out0;
assign v$G11_11575_out0 = v$G_10503_out0;
assign v$G11_11578_out0 = v$G_10575_out0;
assign v$SEL5_12232_out0 = v$AMOUNT$OF$SHIFT_9833_out0[4:4];
assign v$SEL5_12233_out0 = v$AMOUNT$OF$SHIFT_9834_out0[4:4];
assign v$SEL5_12234_out0 = v$AMOUNT$OF$SHIFT_9835_out0[4:4];
assign v$SEL5_12235_out0 = v$AMOUNT$OF$SHIFT_9836_out0[4:4];
assign v$P17_12328_out0 = v$P_14463_out0;
assign v$P17_12331_out0 = v$P_14535_out0;
assign v$P7_12338_out0 = v$P_14458_out0;
assign v$P7_12341_out0 = v$P_14530_out0;
assign v$G22_13104_out0 = v$G_10498_out0;
assign v$G22_13107_out0 = v$G_10570_out0;
assign v$SEL1_13940_out0 = v$AMOUNT$OF$SHIFT_9833_out0[0:0];
assign v$SEL1_13941_out0 = v$AMOUNT$OF$SHIFT_9834_out0[0:0];
assign v$SEL1_13942_out0 = v$AMOUNT$OF$SHIFT_9835_out0[0:0];
assign v$SEL1_13943_out0 = v$AMOUNT$OF$SHIFT_9836_out0[0:0];
assign v$P4_14214_out0 = v$P_14467_out0;
assign v$P4_14217_out0 = v$P_14539_out0;
assign v$SEL3_14614_out0 = v$AMOUNT$OF$SHIFT_9833_out0[2:2];
assign v$SEL3_14615_out0 = v$AMOUNT$OF$SHIFT_9834_out0[2:2];
assign v$SEL3_14616_out0 = v$AMOUNT$OF$SHIFT_9835_out0[2:2];
assign v$SEL3_14617_out0 = v$AMOUNT$OF$SHIFT_9836_out0[2:2];
assign v$G23_14920_out0 = v$G_10493_out0;
assign v$G23_14923_out0 = v$G_10565_out0;
assign v$GATE2_16355_out0 = v$CIN_16717_out0 && v$P0_5023_out0;
assign v$GATE2_16358_out0 = v$CIN_16720_out0 && v$P0_5026_out0;
assign v$G2_16568_out0 = v$G_10502_out0;
assign v$G2_16571_out0 = v$G_10574_out0;
assign v$P19_16932_out0 = v$P_14468_out0;
assign v$P19_16935_out0 = v$P_14540_out0;
assign v$G16_17071_out0 = v$G_10505_out0;
assign v$G16_17074_out0 = v$G_10577_out0;
assign v$G14_18593_out0 = v$G_10489_out0;
assign v$G14_18596_out0 = v$G_10561_out0;
assign v$SEL2_19113_out0 = v$AMOUNT$OF$SHIFT_9833_out0[1:1];
assign v$SEL2_19114_out0 = v$AMOUNT$OF$SHIFT_9834_out0[1:1];
assign v$SEL2_19115_out0 = v$AMOUNT$OF$SHIFT_9835_out0[1:1];
assign v$SEL2_19116_out0 = v$AMOUNT$OF$SHIFT_9836_out0[1:1];
assign v$GATE1_720_out0 = v$GATE2_16355_out0 || v$G0_16548_out0;
assign v$GATE1_723_out0 = v$GATE2_16358_out0 || v$G0_16551_out0;
assign v$G$CD_1018_out0 = v$G14_18593_out0;
assign v$G$CD_1019_out0 = v$G8_2770_out0;
assign v$G$CD_1021_out0 = v$G1_5269_out0;
assign v$G$CD_1024_out0 = v$G19_2044_out0;
assign v$G$CD_1025_out0 = v$G22_13104_out0;
assign v$G$CD_1032_out0 = v$G23_14920_out0;
assign v$G$CD_1034_out0 = v$G2_16568_out0;
assign v$G$CD_1035_out0 = v$G5_11170_out0;
assign v$G$CD_1037_out0 = v$G13_3052_out0;
assign v$G$CD_1038_out0 = v$G17_9714_out0;
assign v$G$CD_1039_out0 = v$G16_17071_out0;
assign v$G$CD_1042_out0 = v$G7_1849_out0;
assign v$G$CD_1048_out0 = v$G4_6019_out0;
assign v$G$CD_1052_out0 = v$G20_8533_out0;
assign v$G$CD_1053_out0 = v$G10_1993_out0;
assign v$G$CD_1057_out0 = v$G11_11575_out0;
assign v$G$CD_1141_out0 = v$G14_18596_out0;
assign v$G$CD_1142_out0 = v$G8_2773_out0;
assign v$G$CD_1144_out0 = v$G1_5272_out0;
assign v$G$CD_1147_out0 = v$G19_2047_out0;
assign v$G$CD_1148_out0 = v$G22_13107_out0;
assign v$G$CD_1155_out0 = v$G23_14923_out0;
assign v$G$CD_1157_out0 = v$G2_16571_out0;
assign v$G$CD_1158_out0 = v$G5_11173_out0;
assign v$G$CD_1160_out0 = v$G13_3055_out0;
assign v$G$CD_1161_out0 = v$G17_9717_out0;
assign v$G$CD_1162_out0 = v$G16_17074_out0;
assign v$G$CD_1165_out0 = v$G7_1852_out0;
assign v$G$CD_1171_out0 = v$G4_6022_out0;
assign v$G$CD_1175_out0 = v$G20_8536_out0;
assign v$G$CD_1176_out0 = v$G10_1996_out0;
assign v$G$CD_1180_out0 = v$G11_11578_out0;
assign v$MUX7_1378_out0 = v$EQ7_4242_out0 ? v$SEL7_14936_out0 : v$MUX9_8553_out0;
assign v$MUX7_1379_out0 = v$EQ7_4243_out0 ? v$SEL7_14937_out0 : v$MUX9_8554_out0;
assign v$MUX7_1380_out0 = v$EQ7_4244_out0 ? v$SEL7_14938_out0 : v$MUX9_8555_out0;
assign v$MUX7_1381_out0 = v$EQ7_4245_out0 ? v$SEL7_14939_out0 : v$MUX9_8556_out0;
assign v$EN_1499_out0 = v$SEL4_2005_out0;
assign v$EN_1502_out0 = v$SEL4_2006_out0;
assign v$EN_1509_out0 = v$SEL4_2007_out0;
assign v$EN_1512_out0 = v$SEL4_2008_out0;
assign v$EN_4054_out0 = v$SEL1_13940_out0;
assign v$EN_4055_out0 = v$SEL1_13941_out0;
assign v$EN_4057_out0 = v$SEL1_13942_out0;
assign v$EN_4058_out0 = v$SEL1_13943_out0;
assign v$EN_4966_out0 = v$SEL3_14614_out0;
assign v$EN_4968_out0 = v$SEL3_14615_out0;
assign v$EN_4972_out0 = v$SEL3_14616_out0;
assign v$EN_4974_out0 = v$SEL3_14617_out0;
assign v$EN_5430_out0 = v$SEL5_12232_out0;
assign v$EN_5432_out0 = v$SEL5_12233_out0;
assign v$EN_5436_out0 = v$SEL5_12234_out0;
assign v$EN_5438_out0 = v$SEL5_12235_out0;
assign v$EN_8202_out0 = v$SEL2_19113_out0;
assign v$EN_8204_out0 = v$SEL2_19114_out0;
assign v$EN_8208_out0 = v$SEL2_19115_out0;
assign v$EN_8210_out0 = v$SEL2_19116_out0;
assign v$P$CD_10907_out0 = v$P14_3369_out0;
assign v$P$CD_10908_out0 = v$P8_1861_out0;
assign v$P$CD_10910_out0 = v$P1_3168_out0;
assign v$P$CD_10913_out0 = v$P19_16932_out0;
assign v$P$CD_10914_out0 = v$P22_4945_out0;
assign v$P$CD_10921_out0 = v$P23_6626_out0;
assign v$P$CD_10923_out0 = v$P2_2424_out0;
assign v$P$CD_10924_out0 = v$P5_228_out0;
assign v$P$CD_10926_out0 = v$P13_3245_out0;
assign v$P$CD_10927_out0 = v$P17_12328_out0;
assign v$P$CD_10928_out0 = v$P16_7243_out0;
assign v$P$CD_10931_out0 = v$P7_12338_out0;
assign v$P$CD_10937_out0 = v$P4_14214_out0;
assign v$P$CD_10941_out0 = v$P20_11152_out0;
assign v$P$CD_10942_out0 = v$P10_360_out0;
assign v$P$CD_10946_out0 = v$P11_9992_out0;
assign v$P$CD_11030_out0 = v$P14_3372_out0;
assign v$P$CD_11031_out0 = v$P8_1864_out0;
assign v$P$CD_11033_out0 = v$P1_3171_out0;
assign v$P$CD_11036_out0 = v$P19_16935_out0;
assign v$P$CD_11037_out0 = v$P22_4948_out0;
assign v$P$CD_11044_out0 = v$P23_6629_out0;
assign v$P$CD_11046_out0 = v$P2_2427_out0;
assign v$P$CD_11047_out0 = v$P5_231_out0;
assign v$P$CD_11049_out0 = v$P13_3248_out0;
assign v$P$CD_11050_out0 = v$P17_12331_out0;
assign v$P$CD_11051_out0 = v$P16_7246_out0;
assign v$P$CD_11054_out0 = v$P7_12341_out0;
assign v$P$CD_11060_out0 = v$P4_14217_out0;
assign v$P$CD_11064_out0 = v$P20_11155_out0;
assign v$P$CD_11065_out0 = v$P10_363_out0;
assign v$P$CD_11069_out0 = v$P11_9995_out0;
assign v$G8_11929_out0 = v$CINA_8774_out0 && v$P$AB_2168_out0;
assign v$G8_11932_out0 = v$CINA_8777_out0 && v$P$AB_2171_out0;
assign v$G8_11933_out0 = v$CINA_8778_out0 && v$P$AB_2172_out0;
assign v$G8_11945_out0 = v$CINA_8790_out0 && v$P$AB_2184_out0;
assign v$G8_11947_out0 = v$CINA_8792_out0 && v$P$AB_2186_out0;
assign v$G8_11950_out0 = v$CINA_8795_out0 && v$P$AB_2189_out0;
assign v$G8_11956_out0 = v$CINA_8801_out0 && v$P$AB_2195_out0;
assign v$G8_11961_out0 = v$CINA_8806_out0 && v$P$AB_2200_out0;
assign v$G8_12052_out0 = v$CINA_8897_out0 && v$P$AB_2291_out0;
assign v$G8_12055_out0 = v$CINA_8900_out0 && v$P$AB_2294_out0;
assign v$G8_12056_out0 = v$CINA_8901_out0 && v$P$AB_2295_out0;
assign v$G8_12068_out0 = v$CINA_8913_out0 && v$P$AB_2307_out0;
assign v$G8_12070_out0 = v$CINA_8915_out0 && v$P$AB_2309_out0;
assign v$G8_12073_out0 = v$CINA_8918_out0 && v$P$AB_2312_out0;
assign v$G8_12079_out0 = v$CINA_8924_out0 && v$P$AB_2318_out0;
assign v$G8_12084_out0 = v$CINA_8929_out0 && v$P$AB_2323_out0;
assign v$G5_4693_out0 = v$G$AB_9468_out0 && v$P$CD_10910_out0;
assign v$G5_4696_out0 = v$G$AB_9471_out0 && v$P$CD_10913_out0;
assign v$G5_4697_out0 = v$G$AB_9472_out0 && v$P$CD_10914_out0;
assign v$G5_4709_out0 = v$G$AB_9484_out0 && v$P$CD_10926_out0;
assign v$G5_4711_out0 = v$G$AB_9486_out0 && v$P$CD_10928_out0;
assign v$G5_4714_out0 = v$G$AB_9489_out0 && v$P$CD_10931_out0;
assign v$G5_4720_out0 = v$G$AB_9495_out0 && v$P$CD_10937_out0;
assign v$G5_4725_out0 = v$G$AB_9500_out0 && v$P$CD_10942_out0;
assign v$G5_4816_out0 = v$G$AB_9591_out0 && v$P$CD_11033_out0;
assign v$G5_4819_out0 = v$G$AB_9594_out0 && v$P$CD_11036_out0;
assign v$G5_4820_out0 = v$G$AB_9595_out0 && v$P$CD_11037_out0;
assign v$G5_4832_out0 = v$G$AB_9607_out0 && v$P$CD_11049_out0;
assign v$G5_4834_out0 = v$G$AB_9609_out0 && v$P$CD_11051_out0;
assign v$G5_4837_out0 = v$G$AB_9612_out0 && v$P$CD_11054_out0;
assign v$G5_4843_out0 = v$G$AB_9618_out0 && v$P$CD_11060_out0;
assign v$G5_4848_out0 = v$G$AB_9623_out0 && v$P$CD_11065_out0;
assign v$G1_5767_out0 = v$P$AB_2168_out0 && v$P$CD_10910_out0;
assign v$G1_5770_out0 = v$P$AB_2171_out0 && v$P$CD_10913_out0;
assign v$G1_5771_out0 = v$P$AB_2172_out0 && v$P$CD_10914_out0;
assign v$G1_5783_out0 = v$P$AB_2184_out0 && v$P$CD_10926_out0;
assign v$G1_5785_out0 = v$P$AB_2186_out0 && v$P$CD_10928_out0;
assign v$G1_5788_out0 = v$P$AB_2189_out0 && v$P$CD_10931_out0;
assign v$G1_5794_out0 = v$P$AB_2195_out0 && v$P$CD_10937_out0;
assign v$G1_5799_out0 = v$P$AB_2200_out0 && v$P$CD_10942_out0;
assign v$G1_5890_out0 = v$P$AB_2291_out0 && v$P$CD_11033_out0;
assign v$G1_5893_out0 = v$P$AB_2294_out0 && v$P$CD_11036_out0;
assign v$G1_5894_out0 = v$P$AB_2295_out0 && v$P$CD_11037_out0;
assign v$G1_5906_out0 = v$P$AB_2307_out0 && v$P$CD_11049_out0;
assign v$G1_5908_out0 = v$P$AB_2309_out0 && v$P$CD_11051_out0;
assign v$G1_5911_out0 = v$P$AB_2312_out0 && v$P$CD_11054_out0;
assign v$G1_5917_out0 = v$P$AB_2318_out0 && v$P$CD_11060_out0;
assign v$G1_5922_out0 = v$P$AB_2323_out0 && v$P$CD_11065_out0;
assign v$G7_10021_out0 = v$G8_11929_out0 && v$P$CD_10910_out0;
assign v$G7_10024_out0 = v$G8_11932_out0 && v$P$CD_10913_out0;
assign v$G7_10025_out0 = v$G8_11933_out0 && v$P$CD_10914_out0;
assign v$G7_10037_out0 = v$G8_11945_out0 && v$P$CD_10926_out0;
assign v$G7_10039_out0 = v$G8_11947_out0 && v$P$CD_10928_out0;
assign v$G7_10042_out0 = v$G8_11950_out0 && v$P$CD_10931_out0;
assign v$G7_10048_out0 = v$G8_11956_out0 && v$P$CD_10937_out0;
assign v$G7_10053_out0 = v$G8_11961_out0 && v$P$CD_10942_out0;
assign v$G7_10144_out0 = v$G8_12052_out0 && v$P$CD_11033_out0;
assign v$G7_10147_out0 = v$G8_12055_out0 && v$P$CD_11036_out0;
assign v$G7_10148_out0 = v$G8_12056_out0 && v$P$CD_11037_out0;
assign v$G7_10160_out0 = v$G8_12068_out0 && v$P$CD_11049_out0;
assign v$G7_10162_out0 = v$G8_12070_out0 && v$P$CD_11051_out0;
assign v$G7_10165_out0 = v$G8_12073_out0 && v$P$CD_11054_out0;
assign v$G7_10171_out0 = v$G8_12079_out0 && v$P$CD_11060_out0;
assign v$G7_10176_out0 = v$G8_12084_out0 && v$P$CD_11065_out0;
assign v$C0_11188_out0 = v$GATE1_720_out0;
assign v$C0_11191_out0 = v$GATE1_723_out0;
assign v$MUX2_15434_out0 = v$EN_4054_out0 ? v$MUX1_2558_out0 : v$IN_4039_out0;
assign v$MUX2_15435_out0 = v$EN_4055_out0 ? v$MUX1_2568_out0 : v$IN_4042_out0;
assign v$MUX2_15437_out0 = v$EN_4057_out0 ? v$MUX1_2589_out0 : v$IN_4048_out0;
assign v$MUX2_15438_out0 = v$EN_4058_out0 ? v$MUX1_2599_out0 : v$IN_4051_out0;
assign v$MUX6_16898_out0 = v$EQ6_5666_out0 ? v$SEL6_13066_out0 : v$MUX7_1378_out0;
assign v$MUX6_16899_out0 = v$EQ6_5667_out0 ? v$SEL6_13067_out0 : v$MUX7_1379_out0;
assign v$MUX6_16900_out0 = v$EQ6_5668_out0 ? v$SEL6_13068_out0 : v$MUX7_1380_out0;
assign v$MUX6_16901_out0 = v$EQ6_5669_out0 ? v$SEL6_13069_out0 : v$MUX7_1381_out0;
assign v$P$AD_754_out0 = v$G1_5767_out0;
assign v$P$AD_757_out0 = v$G1_5770_out0;
assign v$P$AD_758_out0 = v$G1_5771_out0;
assign v$P$AD_770_out0 = v$G1_5783_out0;
assign v$P$AD_772_out0 = v$G1_5785_out0;
assign v$P$AD_775_out0 = v$G1_5788_out0;
assign v$P$AD_781_out0 = v$G1_5794_out0;
assign v$P$AD_786_out0 = v$G1_5799_out0;
assign v$P$AD_877_out0 = v$G1_5890_out0;
assign v$P$AD_880_out0 = v$G1_5893_out0;
assign v$P$AD_881_out0 = v$G1_5894_out0;
assign v$P$AD_893_out0 = v$G1_5906_out0;
assign v$P$AD_895_out0 = v$G1_5908_out0;
assign v$P$AD_898_out0 = v$G1_5911_out0;
assign v$P$AD_904_out0 = v$G1_5917_out0;
assign v$P$AD_909_out0 = v$G1_5922_out0;
assign {v$A2A_1788_out1,v$A2A_1788_out0 } = v$A1_1869_out0 + v$B1_8426_out0 + v$C0_11188_out0;
assign {v$A2A_1791_out1,v$A2A_1791_out0 } = v$A1_1872_out0 + v$B1_8429_out0 + v$C0_11191_out0;
assign v$MUX5_7209_out0 = v$EQ5_3537_out0 ? v$SEL5_16038_out0 : v$MUX6_16898_out0;
assign v$MUX5_7210_out0 = v$EQ5_3538_out0 ? v$SEL5_16039_out0 : v$MUX6_16899_out0;
assign v$MUX5_7211_out0 = v$EQ5_3539_out0 ? v$SEL5_16040_out0 : v$MUX6_16900_out0;
assign v$MUX5_7212_out0 = v$EQ5_3540_out0 ? v$SEL5_16041_out0 : v$MUX6_16901_out0;
assign v$C0_9745_out0 = v$C0_11188_out0;
assign v$C0_9748_out0 = v$C0_11191_out0;
assign v$G4_11614_out0 = v$G5_4693_out0 || v$G$CD_1021_out0;
assign v$G4_11617_out0 = v$G5_4696_out0 || v$G$CD_1024_out0;
assign v$G4_11618_out0 = v$G5_4697_out0 || v$G$CD_1025_out0;
assign v$G4_11630_out0 = v$G5_4709_out0 || v$G$CD_1037_out0;
assign v$G4_11632_out0 = v$G5_4711_out0 || v$G$CD_1039_out0;
assign v$G4_11635_out0 = v$G5_4714_out0 || v$G$CD_1042_out0;
assign v$G4_11641_out0 = v$G5_4720_out0 || v$G$CD_1048_out0;
assign v$G4_11646_out0 = v$G5_4725_out0 || v$G$CD_1053_out0;
assign v$G4_11737_out0 = v$G5_4816_out0 || v$G$CD_1144_out0;
assign v$G4_11740_out0 = v$G5_4819_out0 || v$G$CD_1147_out0;
assign v$G4_11741_out0 = v$G5_4820_out0 || v$G$CD_1148_out0;
assign v$G4_11753_out0 = v$G5_4832_out0 || v$G$CD_1160_out0;
assign v$G4_11755_out0 = v$G5_4834_out0 || v$G$CD_1162_out0;
assign v$G4_11758_out0 = v$G5_4837_out0 || v$G$CD_1165_out0;
assign v$G4_11764_out0 = v$G5_4843_out0 || v$G$CD_1171_out0;
assign v$G4_11769_out0 = v$G5_4848_out0 || v$G$CD_1176_out0;
assign v$OUT_15530_out0 = v$MUX2_15434_out0;
assign v$OUT_15540_out0 = v$MUX2_15435_out0;
assign v$OUT_15561_out0 = v$MUX2_15437_out0;
assign v$OUT_15571_out0 = v$MUX2_15438_out0;
assign v$G6_456_out0 = v$G4_11614_out0 || v$G7_10021_out0;
assign v$G6_459_out0 = v$G4_11617_out0 || v$G7_10024_out0;
assign v$G6_460_out0 = v$G4_11618_out0 || v$G7_10025_out0;
assign v$G6_472_out0 = v$G4_11630_out0 || v$G7_10037_out0;
assign v$G6_474_out0 = v$G4_11632_out0 || v$G7_10039_out0;
assign v$G6_477_out0 = v$G4_11635_out0 || v$G7_10042_out0;
assign v$G6_483_out0 = v$G4_11641_out0 || v$G7_10048_out0;
assign v$G6_488_out0 = v$G4_11646_out0 || v$G7_10053_out0;
assign v$G6_579_out0 = v$G4_11737_out0 || v$G7_10144_out0;
assign v$G6_582_out0 = v$G4_11740_out0 || v$G7_10147_out0;
assign v$G6_583_out0 = v$G4_11741_out0 || v$G7_10148_out0;
assign v$G6_595_out0 = v$G4_11753_out0 || v$G7_10160_out0;
assign v$G6_597_out0 = v$G4_11755_out0 || v$G7_10162_out0;
assign v$G6_600_out0 = v$G4_11758_out0 || v$G7_10165_out0;
assign v$G6_606_out0 = v$G4_11764_out0 || v$G7_10171_out0;
assign v$G6_611_out0 = v$G4_11769_out0 || v$G7_10176_out0;
assign v$END1_1697_out0 = v$A2A_1788_out1;
assign v$END1_1700_out0 = v$A2A_1791_out1;
assign v$P$AB_2165_out0 = v$P$AD_770_out0;
assign v$P$AB_2166_out0 = v$P$AD_775_out0;
assign v$P$AB_2179_out0 = v$P$AD_758_out0;
assign v$P$AB_2181_out0 = v$P$AD_754_out0;
assign v$P$AB_2182_out0 = v$P$AD_781_out0;
assign v$P$AB_2185_out0 = v$P$AD_772_out0;
assign v$P$AB_2199_out0 = v$P$AD_757_out0;
assign v$P$AB_2204_out0 = v$P$AD_786_out0;
assign v$P$AB_2288_out0 = v$P$AD_893_out0;
assign v$P$AB_2289_out0 = v$P$AD_898_out0;
assign v$P$AB_2302_out0 = v$P$AD_881_out0;
assign v$P$AB_2304_out0 = v$P$AD_877_out0;
assign v$P$AB_2305_out0 = v$P$AD_904_out0;
assign v$P$AB_2308_out0 = v$P$AD_895_out0;
assign v$P$AB_2322_out0 = v$P$AD_880_out0;
assign v$P$AB_2327_out0 = v$P$AD_909_out0;
assign v$IN_5384_out0 = v$OUT_15530_out0;
assign v$IN_5394_out0 = v$OUT_15540_out0;
assign v$IN_5415_out0 = v$OUT_15561_out0;
assign v$IN_5425_out0 = v$OUT_15571_out0;
assign v$MUX4_8124_out0 = v$EQ4_19209_out0 ? v$SEL4_7639_out0 : v$MUX5_7209_out0;
assign v$MUX4_8125_out0 = v$EQ4_19210_out0 ? v$SEL4_7640_out0 : v$MUX5_7210_out0;
assign v$MUX4_8126_out0 = v$EQ4_19211_out0 ? v$SEL4_7641_out0 : v$MUX5_7211_out0;
assign v$MUX4_8127_out0 = v$EQ4_19212_out0 ? v$SEL4_7642_out0 : v$MUX5_7212_out0;
assign v$P$CD_10911_out0 = v$P$AD_781_out0;
assign v$P$CD_10915_out0 = v$P$AD_758_out0;
assign v$P$CD_10936_out0 = v$P$AD_772_out0;
assign v$P$CD_10939_out0 = v$P$AD_770_out0;
assign v$P$CD_10940_out0 = v$P$AD_786_out0;
assign v$P$CD_10944_out0 = v$P$AD_757_out0;
assign v$P$CD_10945_out0 = v$P$AD_775_out0;
assign v$P$CD_11034_out0 = v$P$AD_904_out0;
assign v$P$CD_11038_out0 = v$P$AD_881_out0;
assign v$P$CD_11059_out0 = v$P$AD_895_out0;
assign v$P$CD_11062_out0 = v$P$AD_893_out0;
assign v$P$CD_11063_out0 = v$P$AD_909_out0;
assign v$P$CD_11067_out0 = v$P$AD_880_out0;
assign v$P$CD_11068_out0 = v$P$AD_898_out0;
assign v$_14021_out0 = { v$A1A_12224_out0,v$A2A_1788_out0 };
assign v$_14024_out0 = { v$A1A_12227_out0,v$A2A_1791_out0 };
assign v$G$AD_17688_out0 = v$G4_11614_out0;
assign v$G$AD_17691_out0 = v$G4_11617_out0;
assign v$G$AD_17692_out0 = v$G4_11618_out0;
assign v$G$AD_17704_out0 = v$G4_11630_out0;
assign v$G$AD_17706_out0 = v$G4_11632_out0;
assign v$G$AD_17709_out0 = v$G4_11635_out0;
assign v$G$AD_17715_out0 = v$G4_11641_out0;
assign v$G$AD_17720_out0 = v$G4_11646_out0;
assign v$G$AD_17811_out0 = v$G4_11737_out0;
assign v$G$AD_17814_out0 = v$G4_11740_out0;
assign v$G$AD_17815_out0 = v$G4_11741_out0;
assign v$G$AD_17827_out0 = v$G4_11753_out0;
assign v$G$AD_17829_out0 = v$G4_11755_out0;
assign v$G$AD_17832_out0 = v$G4_11758_out0;
assign v$G$AD_17838_out0 = v$G4_11764_out0;
assign v$G$AD_17843_out0 = v$G4_11769_out0;
assign v$G$CD_1022_out0 = v$G$AD_17715_out0;
assign v$G$CD_1026_out0 = v$G$AD_17692_out0;
assign v$G$CD_1047_out0 = v$G$AD_17706_out0;
assign v$G$CD_1050_out0 = v$G$AD_17704_out0;
assign v$G$CD_1051_out0 = v$G$AD_17720_out0;
assign v$G$CD_1055_out0 = v$G$AD_17691_out0;
assign v$G$CD_1056_out0 = v$G$AD_17709_out0;
assign v$G$CD_1145_out0 = v$G$AD_17838_out0;
assign v$G$CD_1149_out0 = v$G$AD_17815_out0;
assign v$G$CD_1170_out0 = v$G$AD_17829_out0;
assign v$G$CD_1173_out0 = v$G$AD_17827_out0;
assign v$G$CD_1174_out0 = v$G$AD_17843_out0;
assign v$G$CD_1178_out0 = v$G$AD_17814_out0;
assign v$G$CD_1179_out0 = v$G$AD_17832_out0;
assign v$G1_5764_out0 = v$P$AB_2165_out0 && v$P$CD_10907_out0;
assign v$G1_5765_out0 = v$P$AB_2166_out0 && v$P$CD_10908_out0;
assign v$G1_5778_out0 = v$P$AB_2179_out0 && v$P$CD_10921_out0;
assign v$G1_5780_out0 = v$P$AB_2181_out0 && v$P$CD_10923_out0;
assign v$G1_5781_out0 = v$P$AB_2182_out0 && v$P$CD_10924_out0;
assign v$G1_5784_out0 = v$P$AB_2185_out0 && v$P$CD_10927_out0;
assign v$G1_5798_out0 = v$P$AB_2199_out0 && v$P$CD_10941_out0;
assign v$G1_5803_out0 = v$P$AB_2204_out0 && v$P$CD_10946_out0;
assign v$G1_5887_out0 = v$P$AB_2288_out0 && v$P$CD_11030_out0;
assign v$G1_5888_out0 = v$P$AB_2289_out0 && v$P$CD_11031_out0;
assign v$G1_5901_out0 = v$P$AB_2302_out0 && v$P$CD_11044_out0;
assign v$G1_5903_out0 = v$P$AB_2304_out0 && v$P$CD_11046_out0;
assign v$G1_5904_out0 = v$P$AB_2305_out0 && v$P$CD_11047_out0;
assign v$G1_5907_out0 = v$P$AB_2308_out0 && v$P$CD_11050_out0;
assign v$G1_5921_out0 = v$P$AB_2322_out0 && v$P$CD_11064_out0;
assign v$G1_5926_out0 = v$P$AB_2327_out0 && v$P$CD_11069_out0;
assign v$COUTD_6934_out0 = v$G6_456_out0;
assign v$COUTD_6937_out0 = v$G6_459_out0;
assign v$COUTD_6938_out0 = v$G6_460_out0;
assign v$COUTD_6950_out0 = v$G6_472_out0;
assign v$COUTD_6952_out0 = v$G6_474_out0;
assign v$COUTD_6955_out0 = v$G6_477_out0;
assign v$COUTD_6961_out0 = v$G6_483_out0;
assign v$COUTD_6966_out0 = v$G6_488_out0;
assign v$COUTD_7057_out0 = v$G6_579_out0;
assign v$COUTD_7060_out0 = v$G6_582_out0;
assign v$COUTD_7061_out0 = v$G6_583_out0;
assign v$COUTD_7073_out0 = v$G6_595_out0;
assign v$COUTD_7075_out0 = v$G6_597_out0;
assign v$COUTD_7078_out0 = v$G6_600_out0;
assign v$COUTD_7084_out0 = v$G6_606_out0;
assign v$COUTD_7089_out0 = v$G6_611_out0;
assign v$MUX3_7928_out0 = v$EQ3_1977_out0 ? v$SEL3_12298_out0 : v$MUX4_8124_out0;
assign v$MUX3_7929_out0 = v$EQ3_1978_out0 ? v$SEL3_12299_out0 : v$MUX4_8125_out0;
assign v$MUX3_7930_out0 = v$EQ3_1979_out0 ? v$SEL3_12300_out0 : v$MUX4_8126_out0;
assign v$MUX3_7931_out0 = v$EQ3_1980_out0 ? v$SEL3_12301_out0 : v$MUX4_8127_out0;
assign v$G$AB_9465_out0 = v$G$AD_17704_out0;
assign v$G$AB_9466_out0 = v$G$AD_17709_out0;
assign v$G$AB_9479_out0 = v$G$AD_17692_out0;
assign v$G$AB_9481_out0 = v$G$AD_17688_out0;
assign v$G$AB_9482_out0 = v$G$AD_17715_out0;
assign v$G$AB_9485_out0 = v$G$AD_17706_out0;
assign v$G$AB_9499_out0 = v$G$AD_17691_out0;
assign v$G$AB_9504_out0 = v$G$AD_17720_out0;
assign v$G$AB_9588_out0 = v$G$AD_17827_out0;
assign v$G$AB_9589_out0 = v$G$AD_17832_out0;
assign v$G$AB_9602_out0 = v$G$AD_17815_out0;
assign v$G$AB_9604_out0 = v$G$AD_17811_out0;
assign v$G$AB_9605_out0 = v$G$AD_17838_out0;
assign v$G$AB_9608_out0 = v$G$AD_17829_out0;
assign v$G$AB_9622_out0 = v$G$AD_17814_out0;
assign v$G$AB_9627_out0 = v$G$AD_17843_out0;
assign v$IN_12355_out0 = v$IN_5384_out0;
assign v$IN_12357_out0 = v$IN_5394_out0;
assign v$IN_12361_out0 = v$IN_5415_out0;
assign v$IN_12363_out0 = v$IN_5425_out0;
assign v$P$AD_751_out0 = v$G1_5764_out0;
assign v$P$AD_752_out0 = v$G1_5765_out0;
assign v$P$AD_765_out0 = v$G1_5778_out0;
assign v$P$AD_767_out0 = v$G1_5780_out0;
assign v$P$AD_768_out0 = v$G1_5781_out0;
assign v$P$AD_771_out0 = v$G1_5784_out0;
assign v$P$AD_785_out0 = v$G1_5798_out0;
assign v$P$AD_790_out0 = v$G1_5803_out0;
assign v$P$AD_874_out0 = v$G1_5887_out0;
assign v$P$AD_875_out0 = v$G1_5888_out0;
assign v$P$AD_888_out0 = v$G1_5901_out0;
assign v$P$AD_890_out0 = v$G1_5903_out0;
assign v$P$AD_891_out0 = v$G1_5904_out0;
assign v$P$AD_894_out0 = v$G1_5907_out0;
assign v$P$AD_908_out0 = v$G1_5921_out0;
assign v$P$AD_913_out0 = v$G1_5926_out0;
assign v$G5_4690_out0 = v$G$AB_9465_out0 && v$P$CD_10907_out0;
assign v$G5_4691_out0 = v$G$AB_9466_out0 && v$P$CD_10908_out0;
assign v$G5_4704_out0 = v$G$AB_9479_out0 && v$P$CD_10921_out0;
assign v$G5_4706_out0 = v$G$AB_9481_out0 && v$P$CD_10923_out0;
assign v$G5_4707_out0 = v$G$AB_9482_out0 && v$P$CD_10924_out0;
assign v$G5_4710_out0 = v$G$AB_9485_out0 && v$P$CD_10927_out0;
assign v$G5_4724_out0 = v$G$AB_9499_out0 && v$P$CD_10941_out0;
assign v$G5_4729_out0 = v$G$AB_9504_out0 && v$P$CD_10946_out0;
assign v$G5_4813_out0 = v$G$AB_9588_out0 && v$P$CD_11030_out0;
assign v$G5_4814_out0 = v$G$AB_9589_out0 && v$P$CD_11031_out0;
assign v$G5_4827_out0 = v$G$AB_9602_out0 && v$P$CD_11044_out0;
assign v$G5_4829_out0 = v$G$AB_9604_out0 && v$P$CD_11046_out0;
assign v$G5_4830_out0 = v$G$AB_9605_out0 && v$P$CD_11047_out0;
assign v$G5_4833_out0 = v$G$AB_9608_out0 && v$P$CD_11050_out0;
assign v$G5_4847_out0 = v$G$AB_9622_out0 && v$P$CD_11064_out0;
assign v$G5_4852_out0 = v$G$AB_9627_out0 && v$P$CD_11069_out0;
assign v$CINA_8771_out0 = v$COUTD_6950_out0;
assign v$CINA_8772_out0 = v$COUTD_6955_out0;
assign v$CINA_8785_out0 = v$COUTD_6938_out0;
assign v$CINA_8787_out0 = v$COUTD_6934_out0;
assign v$CINA_8788_out0 = v$COUTD_6961_out0;
assign v$CINA_8791_out0 = v$COUTD_6952_out0;
assign v$CINA_8805_out0 = v$COUTD_6937_out0;
assign v$CINA_8810_out0 = v$COUTD_6966_out0;
assign v$CINA_8894_out0 = v$COUTD_7073_out0;
assign v$CINA_8895_out0 = v$COUTD_7078_out0;
assign v$CINA_8908_out0 = v$COUTD_7061_out0;
assign v$CINA_8910_out0 = v$COUTD_7057_out0;
assign v$CINA_8911_out0 = v$COUTD_7084_out0;
assign v$CINA_8914_out0 = v$COUTD_7075_out0;
assign v$CINA_8928_out0 = v$COUTD_7060_out0;
assign v$CINA_8933_out0 = v$COUTD_7089_out0;
assign v$SEL1_9065_out0 = v$IN_12355_out0[23:2];
assign v$SEL1_9075_out0 = v$IN_12357_out0[23:2];
assign v$SEL1_9096_out0 = v$IN_12361_out0[23:2];
assign v$SEL1_9106_out0 = v$IN_12363_out0[23:2];
assign v$MUX2_14185_out0 = v$EQ2_14810_out0 ? v$SEL2_13906_out0 : v$MUX3_7928_out0;
assign v$MUX2_14186_out0 = v$EQ2_14811_out0 ? v$SEL2_13907_out0 : v$MUX3_7929_out0;
assign v$MUX2_14187_out0 = v$EQ2_14812_out0 ? v$SEL2_13908_out0 : v$MUX3_7930_out0;
assign v$MUX2_14188_out0 = v$EQ2_14813_out0 ? v$SEL2_13909_out0 : v$MUX3_7931_out0;
assign v$SEL1_15993_out0 = v$IN_12355_out0[21:0];
assign v$SEL1_16003_out0 = v$IN_12357_out0[21:0];
assign v$SEL1_16024_out0 = v$IN_12361_out0[21:0];
assign v$SEL1_16034_out0 = v$IN_12363_out0[21:0];
assign v$C1_17401_out0 = v$COUTD_6934_out0;
assign v$C1_17404_out0 = v$COUTD_7057_out0;
assign v$P$AB_2164_out0 = v$P$AD_752_out0;
assign v$P$AB_2169_out0 = v$P$AD_767_out0;
assign v$P$AB_2175_out0 = v$P$AD_767_out0;
assign v$P$AB_2178_out0 = v$P$AD_785_out0;
assign v$P$AB_2183_out0 = v$P$AD_751_out0;
assign v$P$AB_2196_out0 = v$P$AD_767_out0;
assign v$P$AB_2287_out0 = v$P$AD_875_out0;
assign v$P$AB_2292_out0 = v$P$AD_890_out0;
assign v$P$AB_2298_out0 = v$P$AD_890_out0;
assign v$P$AB_2301_out0 = v$P$AD_908_out0;
assign v$P$AB_2306_out0 = v$P$AD_874_out0;
assign v$P$AB_2319_out0 = v$P$AD_890_out0;
assign v$MUX1_3078_out0 = v$EQ1_13999_out0 ? v$SEL1_7378_out0 : v$MUX2_14185_out0;
assign v$MUX1_3079_out0 = v$EQ1_14000_out0 ? v$SEL1_7379_out0 : v$MUX2_14186_out0;
assign v$MUX1_3080_out0 = v$EQ1_14001_out0 ? v$SEL1_7380_out0 : v$MUX2_14187_out0;
assign v$MUX1_3081_out0 = v$EQ1_14002_out0 ? v$SEL1_7381_out0 : v$MUX2_14188_out0;
assign v$_4425_out0 = { v$C2_123_out0,v$SEL1_15993_out0 };
assign v$_4435_out0 = { v$C2_133_out0,v$SEL1_16003_out0 };
assign v$_4456_out0 = { v$C2_154_out0,v$SEL1_16024_out0 };
assign v$_4466_out0 = { v$C2_164_out0,v$SEL1_16034_out0 };
assign v$_9326_out0 = { v$SEL1_9065_out0,v$C1_6261_out0 };
assign v$_9336_out0 = { v$SEL1_9075_out0,v$C1_6271_out0 };
assign v$_9357_out0 = { v$SEL1_9096_out0,v$C1_6292_out0 };
assign v$_9367_out0 = { v$SEL1_9106_out0,v$C1_6302_out0 };
assign v$P$CD_10906_out0 = v$P$AD_790_out0;
assign v$P$CD_10912_out0 = v$P$AD_752_out0;
assign v$P$CD_10920_out0 = v$P$AD_765_out0;
assign v$P$CD_10925_out0 = v$P$AD_771_out0;
assign v$P$CD_10929_out0 = v$P$AD_785_out0;
assign v$P$CD_10930_out0 = v$P$AD_751_out0;
assign v$P$CD_10938_out0 = v$P$AD_768_out0;
assign v$P$CD_11029_out0 = v$P$AD_913_out0;
assign v$P$CD_11035_out0 = v$P$AD_875_out0;
assign v$P$CD_11043_out0 = v$P$AD_888_out0;
assign v$P$CD_11048_out0 = v$P$AD_894_out0;
assign v$P$CD_11052_out0 = v$P$AD_908_out0;
assign v$P$CD_11053_out0 = v$P$AD_874_out0;
assign v$P$CD_11061_out0 = v$P$AD_891_out0;
assign v$G4_11611_out0 = v$G5_4690_out0 || v$G$CD_1018_out0;
assign v$G4_11612_out0 = v$G5_4691_out0 || v$G$CD_1019_out0;
assign v$G4_11625_out0 = v$G5_4704_out0 || v$G$CD_1032_out0;
assign v$G4_11627_out0 = v$G5_4706_out0 || v$G$CD_1034_out0;
assign v$G4_11628_out0 = v$G5_4707_out0 || v$G$CD_1035_out0;
assign v$G4_11631_out0 = v$G5_4710_out0 || v$G$CD_1038_out0;
assign v$G4_11645_out0 = v$G5_4724_out0 || v$G$CD_1052_out0;
assign v$G4_11650_out0 = v$G5_4729_out0 || v$G$CD_1057_out0;
assign v$G4_11734_out0 = v$G5_4813_out0 || v$G$CD_1141_out0;
assign v$G4_11735_out0 = v$G5_4814_out0 || v$G$CD_1142_out0;
assign v$G4_11748_out0 = v$G5_4827_out0 || v$G$CD_1155_out0;
assign v$G4_11750_out0 = v$G5_4829_out0 || v$G$CD_1157_out0;
assign v$G4_11751_out0 = v$G5_4830_out0 || v$G$CD_1158_out0;
assign v$G4_11754_out0 = v$G5_4833_out0 || v$G$CD_1161_out0;
assign v$G4_11768_out0 = v$G5_4847_out0 || v$G$CD_1175_out0;
assign v$G4_11773_out0 = v$G5_4852_out0 || v$G$CD_1180_out0;
assign v$G8_11926_out0 = v$CINA_8771_out0 && v$P$AB_2165_out0;
assign v$G8_11927_out0 = v$CINA_8772_out0 && v$P$AB_2166_out0;
assign v$G8_11940_out0 = v$CINA_8785_out0 && v$P$AB_2179_out0;
assign v$G8_11942_out0 = v$CINA_8787_out0 && v$P$AB_2181_out0;
assign v$G8_11943_out0 = v$CINA_8788_out0 && v$P$AB_2182_out0;
assign v$G8_11946_out0 = v$CINA_8791_out0 && v$P$AB_2185_out0;
assign v$G8_11960_out0 = v$CINA_8805_out0 && v$P$AB_2199_out0;
assign v$G8_11965_out0 = v$CINA_8810_out0 && v$P$AB_2204_out0;
assign v$G8_12049_out0 = v$CINA_8894_out0 && v$P$AB_2288_out0;
assign v$G8_12050_out0 = v$CINA_8895_out0 && v$P$AB_2289_out0;
assign v$G8_12063_out0 = v$CINA_8908_out0 && v$P$AB_2302_out0;
assign v$G8_12065_out0 = v$CINA_8910_out0 && v$P$AB_2304_out0;
assign v$G8_12066_out0 = v$CINA_8911_out0 && v$P$AB_2305_out0;
assign v$G8_12069_out0 = v$CINA_8914_out0 && v$P$AB_2308_out0;
assign v$G8_12083_out0 = v$CINA_8928_out0 && v$P$AB_2322_out0;
assign v$G8_12088_out0 = v$CINA_8933_out0 && v$P$AB_2327_out0;
assign v$C1_12421_out0 = v$C1_17401_out0;
assign v$C1_12424_out0 = v$C1_17404_out0;
assign {v$A3A_12525_out1,v$A3A_12525_out0 } = v$A2_18868_out0 + v$B2_3326_out0 + v$C1_17401_out0;
assign {v$A3A_12528_out1,v$A3A_12528_out0 } = v$A2_18871_out0 + v$B2_3329_out0 + v$C1_17404_out0;
assign v$MUX1_2562_out0 = v$LEFT$SHIT_3274_out0 ? v$_4425_out0 : v$_9326_out0;
assign v$MUX1_2572_out0 = v$LEFT$SHIT_3284_out0 ? v$_4435_out0 : v$_9336_out0;
assign v$MUX1_2593_out0 = v$LEFT$SHIT_3305_out0 ? v$_4456_out0 : v$_9357_out0;
assign v$MUX1_2603_out0 = v$LEFT$SHIT_3315_out0 ? v$_4466_out0 : v$_9367_out0;
assign v$END2_5449_out0 = v$A3A_12525_out1;
assign v$END2_5452_out0 = v$A3A_12528_out1;
assign v$G1_5763_out0 = v$P$AB_2164_out0 && v$P$CD_10906_out0;
assign v$G1_5768_out0 = v$P$AB_2169_out0 && v$P$CD_10911_out0;
assign v$G1_5774_out0 = v$P$AB_2175_out0 && v$P$CD_10917_out0;
assign v$G1_5777_out0 = v$P$AB_2178_out0 && v$P$CD_10920_out0;
assign v$G1_5782_out0 = v$P$AB_2183_out0 && v$P$CD_10925_out0;
assign v$G1_5795_out0 = v$P$AB_2196_out0 && v$P$CD_10938_out0;
assign v$G1_5886_out0 = v$P$AB_2287_out0 && v$P$CD_11029_out0;
assign v$G1_5891_out0 = v$P$AB_2292_out0 && v$P$CD_11034_out0;
assign v$G1_5897_out0 = v$P$AB_2298_out0 && v$P$CD_11040_out0;
assign v$G1_5900_out0 = v$P$AB_2301_out0 && v$P$CD_11043_out0;
assign v$G1_5905_out0 = v$P$AB_2306_out0 && v$P$CD_11048_out0;
assign v$G1_5918_out0 = v$P$AB_2319_out0 && v$P$CD_11061_out0;
assign v$MUX25_8708_out0 = v$G2_12476_out0 ? v$C2_15778_out0 : v$MUX1_3078_out0;
assign v$MUX25_8709_out0 = v$G2_12477_out0 ? v$C2_15779_out0 : v$MUX1_3079_out0;
assign v$MUX25_8710_out0 = v$G2_12478_out0 ? v$C2_15780_out0 : v$MUX1_3080_out0;
assign v$MUX25_8711_out0 = v$G2_12479_out0 ? v$C2_15781_out0 : v$MUX1_3081_out0;
assign v$_9235_out0 = { v$C0_9745_out0,v$C1_12421_out0 };
assign v$_9238_out0 = { v$C0_9748_out0,v$C1_12424_out0 };
assign v$G7_10018_out0 = v$G8_11926_out0 && v$P$CD_10907_out0;
assign v$G7_10019_out0 = v$G8_11927_out0 && v$P$CD_10908_out0;
assign v$G7_10032_out0 = v$G8_11940_out0 && v$P$CD_10921_out0;
assign v$G7_10034_out0 = v$G8_11942_out0 && v$P$CD_10923_out0;
assign v$G7_10035_out0 = v$G8_11943_out0 && v$P$CD_10924_out0;
assign v$G7_10038_out0 = v$G8_11946_out0 && v$P$CD_10927_out0;
assign v$G7_10052_out0 = v$G8_11960_out0 && v$P$CD_10941_out0;
assign v$G7_10057_out0 = v$G8_11965_out0 && v$P$CD_10946_out0;
assign v$G7_10141_out0 = v$G8_12049_out0 && v$P$CD_11030_out0;
assign v$G7_10142_out0 = v$G8_12050_out0 && v$P$CD_11031_out0;
assign v$G7_10155_out0 = v$G8_12063_out0 && v$P$CD_11044_out0;
assign v$G7_10157_out0 = v$G8_12065_out0 && v$P$CD_11046_out0;
assign v$G7_10158_out0 = v$G8_12066_out0 && v$P$CD_11047_out0;
assign v$G7_10161_out0 = v$G8_12069_out0 && v$P$CD_11050_out0;
assign v$G7_10175_out0 = v$G8_12083_out0 && v$P$CD_11064_out0;
assign v$G7_10180_out0 = v$G8_12088_out0 && v$P$CD_11069_out0;
assign v$G$AD_17685_out0 = v$G4_11611_out0;
assign v$G$AD_17686_out0 = v$G4_11612_out0;
assign v$G$AD_17699_out0 = v$G4_11625_out0;
assign v$G$AD_17701_out0 = v$G4_11627_out0;
assign v$G$AD_17702_out0 = v$G4_11628_out0;
assign v$G$AD_17705_out0 = v$G4_11631_out0;
assign v$G$AD_17719_out0 = v$G4_11645_out0;
assign v$G$AD_17724_out0 = v$G4_11650_out0;
assign v$G$AD_17808_out0 = v$G4_11734_out0;
assign v$G$AD_17809_out0 = v$G4_11735_out0;
assign v$G$AD_17822_out0 = v$G4_11748_out0;
assign v$G$AD_17824_out0 = v$G4_11750_out0;
assign v$G$AD_17825_out0 = v$G4_11751_out0;
assign v$G$AD_17828_out0 = v$G4_11754_out0;
assign v$G$AD_17842_out0 = v$G4_11768_out0;
assign v$G$AD_17847_out0 = v$G4_11773_out0;
assign v$G6_453_out0 = v$G4_11611_out0 || v$G7_10018_out0;
assign v$G6_454_out0 = v$G4_11612_out0 || v$G7_10019_out0;
assign v$G6_467_out0 = v$G4_11625_out0 || v$G7_10032_out0;
assign v$G6_469_out0 = v$G4_11627_out0 || v$G7_10034_out0;
assign v$G6_470_out0 = v$G4_11628_out0 || v$G7_10035_out0;
assign v$G6_473_out0 = v$G4_11631_out0 || v$G7_10038_out0;
assign v$G6_487_out0 = v$G4_11645_out0 || v$G7_10052_out0;
assign v$G6_492_out0 = v$G4_11650_out0 || v$G7_10057_out0;
assign v$G6_576_out0 = v$G4_11734_out0 || v$G7_10141_out0;
assign v$G6_577_out0 = v$G4_11735_out0 || v$G7_10142_out0;
assign v$G6_590_out0 = v$G4_11748_out0 || v$G7_10155_out0;
assign v$G6_592_out0 = v$G4_11750_out0 || v$G7_10157_out0;
assign v$G6_593_out0 = v$G4_11751_out0 || v$G7_10158_out0;
assign v$G6_596_out0 = v$G4_11754_out0 || v$G7_10161_out0;
assign v$G6_610_out0 = v$G4_11768_out0 || v$G7_10175_out0;
assign v$G6_615_out0 = v$G4_11773_out0 || v$G7_10180_out0;
assign v$P$AD_750_out0 = v$G1_5763_out0;
assign v$P$AD_755_out0 = v$G1_5768_out0;
assign v$P$AD_761_out0 = v$G1_5774_out0;
assign v$P$AD_764_out0 = v$G1_5777_out0;
assign v$P$AD_769_out0 = v$G1_5782_out0;
assign v$P$AD_782_out0 = v$G1_5795_out0;
assign v$P$AD_873_out0 = v$G1_5886_out0;
assign v$P$AD_878_out0 = v$G1_5891_out0;
assign v$P$AD_884_out0 = v$G1_5897_out0;
assign v$P$AD_887_out0 = v$G1_5900_out0;
assign v$P$AD_892_out0 = v$G1_5905_out0;
assign v$P$AD_905_out0 = v$G1_5918_out0;
assign v$G$CD_1017_out0 = v$G$AD_17724_out0;
assign v$G$CD_1023_out0 = v$G$AD_17686_out0;
assign v$G$CD_1031_out0 = v$G$AD_17699_out0;
assign v$G$CD_1036_out0 = v$G$AD_17705_out0;
assign v$G$CD_1040_out0 = v$G$AD_17719_out0;
assign v$G$CD_1041_out0 = v$G$AD_17685_out0;
assign v$G$CD_1049_out0 = v$G$AD_17702_out0;
assign v$G$CD_1140_out0 = v$G$AD_17847_out0;
assign v$G$CD_1146_out0 = v$G$AD_17809_out0;
assign v$G$CD_1154_out0 = v$G$AD_17822_out0;
assign v$G$CD_1159_out0 = v$G$AD_17828_out0;
assign v$G$CD_1163_out0 = v$G$AD_17842_out0;
assign v$G$CD_1164_out0 = v$G$AD_17808_out0;
assign v$G$CD_1172_out0 = v$G$AD_17825_out0;
assign v$MUX2_2673_out0 = v$EN_8202_out0 ? v$MUX1_2562_out0 : v$IN_12355_out0;
assign v$MUX2_2675_out0 = v$EN_8204_out0 ? v$MUX1_2572_out0 : v$IN_12357_out0;
assign v$MUX2_2679_out0 = v$EN_8208_out0 ? v$MUX1_2593_out0 : v$IN_12361_out0;
assign v$MUX2_2681_out0 = v$EN_8210_out0 ? v$MUX1_2603_out0 : v$IN_12363_out0;
assign v$G$AB_9464_out0 = v$G$AD_17686_out0;
assign v$G$AB_9469_out0 = v$G$AD_17701_out0;
assign v$G$AB_9475_out0 = v$G$AD_17701_out0;
assign v$G$AB_9478_out0 = v$G$AD_17719_out0;
assign v$G$AB_9483_out0 = v$G$AD_17685_out0;
assign v$G$AB_9496_out0 = v$G$AD_17701_out0;
assign v$G$AB_9587_out0 = v$G$AD_17809_out0;
assign v$G$AB_9592_out0 = v$G$AD_17824_out0;
assign v$G$AB_9598_out0 = v$G$AD_17824_out0;
assign v$G$AB_9601_out0 = v$G$AD_17842_out0;
assign v$G$AB_9606_out0 = v$G$AD_17808_out0;
assign v$G$AB_9619_out0 = v$G$AD_17824_out0;
assign v$OUT_9851_out0 = v$MUX25_8708_out0;
assign v$OUT_9852_out0 = v$MUX25_8709_out0;
assign v$OUT_9853_out0 = v$MUX25_8710_out0;
assign v$OUT_9854_out0 = v$MUX25_8711_out0;
assign v$P$AB_2170_out0 = v$P$AD_782_out0;
assign v$P$AB_2174_out0 = v$P$AD_782_out0;
assign v$P$AB_2193_out0 = v$P$AD_782_out0;
assign v$P$AB_2201_out0 = v$P$AD_769_out0;
assign v$P$AB_2203_out0 = v$P$AD_782_out0;
assign v$P$AB_2293_out0 = v$P$AD_905_out0;
assign v$P$AB_2297_out0 = v$P$AD_905_out0;
assign v$P$AB_2316_out0 = v$P$AD_905_out0;
assign v$P$AB_2324_out0 = v$P$AD_892_out0;
assign v$P$AB_2326_out0 = v$P$AD_905_out0;
assign {v$A1_2859_out1,v$A1_2859_out0 } = v$LARGER$EXP_10729_out0 + v$SMALLER$EXP_3150_out0 + v$OUT_9851_out0;
assign {v$A1_2860_out1,v$A1_2860_out0 } = v$LARGER$EXP_10730_out0 + v$SMALLER$EXP_3151_out0 + v$OUT_9852_out0;
assign {v$A1_2861_out1,v$A1_2861_out0 } = v$LARGER$EXP_10731_out0 + v$SMALLER$EXP_3152_out0 + v$OUT_9853_out0;
assign {v$A1_2862_out1,v$A1_2862_out0 } = v$LARGER$EXP_10732_out0 + v$SMALLER$EXP_3153_out0 + v$OUT_9854_out0;
assign v$G5_4689_out0 = v$G$AB_9464_out0 && v$P$CD_10906_out0;
assign v$G5_4694_out0 = v$G$AB_9469_out0 && v$P$CD_10911_out0;
assign v$G5_4700_out0 = v$G$AB_9475_out0 && v$P$CD_10917_out0;
assign v$G5_4703_out0 = v$G$AB_9478_out0 && v$P$CD_10920_out0;
assign v$G5_4708_out0 = v$G$AB_9483_out0 && v$P$CD_10925_out0;
assign v$G5_4721_out0 = v$G$AB_9496_out0 && v$P$CD_10938_out0;
assign v$G5_4812_out0 = v$G$AB_9587_out0 && v$P$CD_11029_out0;
assign v$G5_4817_out0 = v$G$AB_9592_out0 && v$P$CD_11034_out0;
assign v$G5_4823_out0 = v$G$AB_9598_out0 && v$P$CD_11040_out0;
assign v$G5_4826_out0 = v$G$AB_9601_out0 && v$P$CD_11043_out0;
assign v$G5_4831_out0 = v$G$AB_9606_out0 && v$P$CD_11048_out0;
assign v$G5_4844_out0 = v$G$AB_9619_out0 && v$P$CD_11061_out0;
assign v$COUTD_6931_out0 = v$G6_453_out0;
assign v$COUTD_6932_out0 = v$G6_454_out0;
assign v$COUTD_6945_out0 = v$G6_467_out0;
assign v$COUTD_6947_out0 = v$G6_469_out0;
assign v$COUTD_6948_out0 = v$G6_470_out0;
assign v$COUTD_6951_out0 = v$G6_473_out0;
assign v$COUTD_6965_out0 = v$G6_487_out0;
assign v$COUTD_6970_out0 = v$G6_492_out0;
assign v$COUTD_7054_out0 = v$G6_576_out0;
assign v$COUTD_7055_out0 = v$G6_577_out0;
assign v$COUTD_7068_out0 = v$G6_590_out0;
assign v$COUTD_7070_out0 = v$G6_592_out0;
assign v$COUTD_7071_out0 = v$G6_593_out0;
assign v$COUTD_7074_out0 = v$G6_596_out0;
assign v$COUTD_7088_out0 = v$G6_610_out0;
assign v$COUTD_7093_out0 = v$G6_615_out0;
assign v$P$CD_10909_out0 = v$P$AD_769_out0;
assign v$P$CD_10935_out0 = v$P$AD_750_out0;
assign v$P$CD_10943_out0 = v$P$AD_764_out0;
assign v$P$CD_11032_out0 = v$P$AD_892_out0;
assign v$P$CD_11058_out0 = v$P$AD_873_out0;
assign v$P$CD_11066_out0 = v$P$AD_887_out0;
assign v$END11_12655_out0 = v$P$AD_761_out0;
assign v$END11_12658_out0 = v$P$AD_884_out0;
assign v$OUT_15534_out0 = v$MUX2_2673_out0;
assign v$OUT_15544_out0 = v$MUX2_2675_out0;
assign v$OUT_15565_out0 = v$MUX2_2679_out0;
assign v$OUT_15575_out0 = v$MUX2_2681_out0;
assign v$END13_18673_out0 = v$P$AD_755_out0;
assign v$END13_18676_out0 = v$P$AD_878_out0;
assign v$END1_1450_out0 = v$COUTD_6970_out0;
assign v$END1_1453_out0 = v$COUTD_7093_out0;
assign v$C2_2884_out0 = v$COUTD_6947_out0;
assign v$C2_2887_out0 = v$COUTD_7070_out0;
assign v$END_3541_out0 = v$COUTD_6948_out0;
assign v$END_3544_out0 = v$COUTD_7071_out0;
assign v$END3_3655_out0 = v$COUTD_6945_out0;
assign v$END3_3658_out0 = v$COUTD_7068_out0;
assign v$IN_5382_out0 = v$OUT_15534_out0;
assign v$IN_5392_out0 = v$OUT_15544_out0;
assign v$IN_5413_out0 = v$OUT_15565_out0;
assign v$IN_5423_out0 = v$OUT_15575_out0;
assign v$G1_5769_out0 = v$P$AB_2170_out0 && v$P$CD_10912_out0;
assign v$G1_5773_out0 = v$P$AB_2174_out0 && v$P$CD_10916_out0;
assign v$G1_5792_out0 = v$P$AB_2193_out0 && v$P$CD_10935_out0;
assign v$G1_5800_out0 = v$P$AB_2201_out0 && v$P$CD_10943_out0;
assign v$G1_5802_out0 = v$P$AB_2203_out0 && v$P$CD_10945_out0;
assign v$G1_5892_out0 = v$P$AB_2293_out0 && v$P$CD_11035_out0;
assign v$G1_5896_out0 = v$P$AB_2297_out0 && v$P$CD_11039_out0;
assign v$G1_5915_out0 = v$P$AB_2316_out0 && v$P$CD_11058_out0;
assign v$G1_5923_out0 = v$P$AB_2324_out0 && v$P$CD_11066_out0;
assign v$G1_5925_out0 = v$P$AB_2326_out0 && v$P$CD_11068_out0;
assign v$END2_8068_out0 = v$COUTD_6951_out0;
assign v$END2_8071_out0 = v$COUTD_7074_out0;
assign v$CINA_8770_out0 = v$COUTD_6932_out0;
assign v$CINA_8775_out0 = v$COUTD_6947_out0;
assign v$CINA_8781_out0 = v$COUTD_6947_out0;
assign v$CINA_8784_out0 = v$COUTD_6965_out0;
assign v$CINA_8789_out0 = v$COUTD_6931_out0;
assign v$CINA_8802_out0 = v$COUTD_6947_out0;
assign v$CINA_8893_out0 = v$COUTD_7055_out0;
assign v$CINA_8898_out0 = v$COUTD_7070_out0;
assign v$CINA_8904_out0 = v$COUTD_7070_out0;
assign v$CINA_8907_out0 = v$COUTD_7088_out0;
assign v$CINA_8912_out0 = v$COUTD_7054_out0;
assign v$CINA_8925_out0 = v$COUTD_7070_out0;
assign v$END45_9383_out0 = v$COUTD_6965_out0;
assign v$END45_9386_out0 = v$COUTD_7088_out0;
assign {v$A2_10470_out1,v$A2_10470_out0 } = v$A1_2859_out0 + v$C1_6236_out0 + v$C2_16894_out0;
assign {v$A2_10471_out1,v$A2_10471_out0 } = v$A1_2860_out0 + v$C1_6237_out0 + v$C2_16895_out0;
assign {v$A2_10472_out1,v$A2_10472_out0 } = v$A1_2861_out0 + v$C1_6238_out0 + v$C2_16896_out0;
assign {v$A2_10473_out1,v$A2_10473_out0 } = v$A1_2862_out0 + v$C1_6239_out0 + v$C2_16897_out0;
assign v$G4_11610_out0 = v$G5_4689_out0 || v$G$CD_1017_out0;
assign v$G4_11615_out0 = v$G5_4694_out0 || v$G$CD_1022_out0;
assign v$G4_11621_out0 = v$G5_4700_out0 || v$G$CD_1028_out0;
assign v$G4_11624_out0 = v$G5_4703_out0 || v$G$CD_1031_out0;
assign v$G4_11629_out0 = v$G5_4708_out0 || v$G$CD_1036_out0;
assign v$G4_11642_out0 = v$G5_4721_out0 || v$G$CD_1049_out0;
assign v$G4_11733_out0 = v$G5_4812_out0 || v$G$CD_1140_out0;
assign v$G4_11738_out0 = v$G5_4817_out0 || v$G$CD_1145_out0;
assign v$G4_11744_out0 = v$G5_4823_out0 || v$G$CD_1151_out0;
assign v$G4_11747_out0 = v$G5_4826_out0 || v$G$CD_1154_out0;
assign v$G4_11752_out0 = v$G5_4831_out0 || v$G$CD_1159_out0;
assign v$G4_11765_out0 = v$G5_4844_out0 || v$G$CD_1172_out0;
assign v$NOT$USED$CARRY_19386_out0 = v$A1_2859_out1;
assign v$NOT$USED$CARRY_19387_out0 = v$A1_2860_out1;
assign v$NOT$USED$CARRY_19388_out0 = v$A1_2861_out1;
assign v$NOT$USED$CARRY_19389_out0 = v$A1_2862_out1;
assign v$P$AD_756_out0 = v$G1_5769_out0;
assign v$P$AD_760_out0 = v$G1_5773_out0;
assign v$P$AD_779_out0 = v$G1_5792_out0;
assign v$P$AD_787_out0 = v$G1_5800_out0;
assign v$P$AD_789_out0 = v$G1_5802_out0;
assign v$P$AD_879_out0 = v$G1_5892_out0;
assign v$P$AD_883_out0 = v$G1_5896_out0;
assign v$P$AD_902_out0 = v$G1_5915_out0;
assign v$P$AD_910_out0 = v$G1_5923_out0;
assign v$P$AD_912_out0 = v$G1_5925_out0;
assign v$G8_11925_out0 = v$CINA_8770_out0 && v$P$AB_2164_out0;
assign v$G8_11930_out0 = v$CINA_8775_out0 && v$P$AB_2169_out0;
assign v$G8_11936_out0 = v$CINA_8781_out0 && v$P$AB_2175_out0;
assign v$G8_11939_out0 = v$CINA_8784_out0 && v$P$AB_2178_out0;
assign v$G8_11944_out0 = v$CINA_8789_out0 && v$P$AB_2183_out0;
assign v$G8_11957_out0 = v$CINA_8802_out0 && v$P$AB_2196_out0;
assign v$G8_12048_out0 = v$CINA_8893_out0 && v$P$AB_2287_out0;
assign v$G8_12053_out0 = v$CINA_8898_out0 && v$P$AB_2292_out0;
assign v$G8_12059_out0 = v$CINA_8904_out0 && v$P$AB_2298_out0;
assign v$G8_12062_out0 = v$CINA_8907_out0 && v$P$AB_2301_out0;
assign v$G8_12067_out0 = v$CINA_8912_out0 && v$P$AB_2306_out0;
assign v$G8_12080_out0 = v$CINA_8925_out0 && v$P$AB_2319_out0;
assign {v$A4A_13731_out1,v$A4A_13731_out0 } = v$A3_15209_out0 + v$B3_9845_out0 + v$C2_2884_out0;
assign {v$A4A_13734_out1,v$A4A_13734_out0 } = v$A3_15212_out0 + v$B3_9848_out0 + v$C2_2887_out0;
assign v$IN_16199_out0 = v$IN_5382_out0;
assign v$IN_16201_out0 = v$IN_5392_out0;
assign v$IN_16205_out0 = v$IN_5413_out0;
assign v$IN_16207_out0 = v$IN_5423_out0;
assign v$NOT$USED_16558_out0 = v$A2_10470_out1;
assign v$NOT$USED_16559_out0 = v$A2_10471_out1;
assign v$NOT$USED_16560_out0 = v$A2_10472_out1;
assign v$NOT$USED_16561_out0 = v$A2_10473_out1;
assign v$G$AD_17684_out0 = v$G4_11610_out0;
assign v$G$AD_17689_out0 = v$G4_11615_out0;
assign v$G$AD_17695_out0 = v$G4_11621_out0;
assign v$G$AD_17698_out0 = v$G4_11624_out0;
assign v$G$AD_17703_out0 = v$G4_11629_out0;
assign v$G$AD_17716_out0 = v$G4_11642_out0;
assign v$G$AD_17807_out0 = v$G4_11733_out0;
assign v$G$AD_17812_out0 = v$G4_11738_out0;
assign v$G$AD_17818_out0 = v$G4_11744_out0;
assign v$G$AD_17821_out0 = v$G4_11747_out0;
assign v$G$AD_17826_out0 = v$G4_11752_out0;
assign v$G$AD_17839_out0 = v$G4_11765_out0;
assign v$C2_18777_out0 = v$C2_2884_out0;
assign v$C2_18780_out0 = v$C2_2887_out0;
assign v$G$CD_1020_out0 = v$G$AD_17703_out0;
assign v$G$CD_1046_out0 = v$G$AD_17684_out0;
assign v$G$CD_1054_out0 = v$G$AD_17698_out0;
assign v$G$CD_1143_out0 = v$G$AD_17826_out0;
assign v$G$CD_1169_out0 = v$G$AD_17807_out0;
assign v$G$CD_1177_out0 = v$G$AD_17821_out0;
assign v$END10_1295_out0 = v$G$AD_17695_out0;
assign v$END10_1298_out0 = v$G$AD_17818_out0;
assign v$P$AB_2167_out0 = v$P$AD_779_out0;
assign v$P$AB_2176_out0 = v$P$AD_779_out0;
assign v$P$AB_2177_out0 = v$P$AD_756_out0;
assign v$P$AB_2188_out0 = v$P$AD_779_out0;
assign v$P$AB_2190_out0 = v$P$AD_779_out0;
assign v$P$AB_2197_out0 = v$P$AD_779_out0;
assign v$P$AB_2198_out0 = v$P$AD_756_out0;
assign v$P$AB_2290_out0 = v$P$AD_902_out0;
assign v$P$AB_2299_out0 = v$P$AD_902_out0;
assign v$P$AB_2300_out0 = v$P$AD_879_out0;
assign v$P$AB_2311_out0 = v$P$AD_902_out0;
assign v$P$AB_2313_out0 = v$P$AD_902_out0;
assign v$P$AB_2320_out0 = v$P$AD_902_out0;
assign v$P$AB_2321_out0 = v$P$AD_879_out0;
assign v$END15_7696_out0 = v$P$AD_760_out0;
assign v$END15_7699_out0 = v$P$AD_883_out0;
assign v$END17_7965_out0 = v$P$AD_789_out0;
assign v$END17_7968_out0 = v$P$AD_912_out0;
assign v$END3_8257_out0 = v$A4A_13731_out1;
assign v$END3_8260_out0 = v$A4A_13734_out1;
assign v$SEL1_9063_out0 = v$IN_16199_out0[23:4];
assign v$SEL1_9073_out0 = v$IN_16201_out0[23:4];
assign v$SEL1_9094_out0 = v$IN_16205_out0[23:4];
assign v$SEL1_9104_out0 = v$IN_16207_out0[23:4];
assign v$G$AB_9470_out0 = v$G$AD_17716_out0;
assign v$G$AB_9474_out0 = v$G$AD_17716_out0;
assign v$G$AB_9493_out0 = v$G$AD_17716_out0;
assign v$G$AB_9501_out0 = v$G$AD_17703_out0;
assign v$G$AB_9503_out0 = v$G$AD_17716_out0;
assign v$G$AB_9593_out0 = v$G$AD_17839_out0;
assign v$G$AB_9597_out0 = v$G$AD_17839_out0;
assign v$G$AB_9616_out0 = v$G$AD_17839_out0;
assign v$G$AB_9624_out0 = v$G$AD_17826_out0;
assign v$G$AB_9626_out0 = v$G$AD_17839_out0;
assign v$G7_10017_out0 = v$G8_11925_out0 && v$P$CD_10906_out0;
assign v$G7_10022_out0 = v$G8_11930_out0 && v$P$CD_10911_out0;
assign v$G7_10028_out0 = v$G8_11936_out0 && v$P$CD_10917_out0;
assign v$G7_10031_out0 = v$G8_11939_out0 && v$P$CD_10920_out0;
assign v$G7_10036_out0 = v$G8_11944_out0 && v$P$CD_10925_out0;
assign v$G7_10049_out0 = v$G8_11957_out0 && v$P$CD_10938_out0;
assign v$G7_10140_out0 = v$G8_12048_out0 && v$P$CD_11029_out0;
assign v$G7_10145_out0 = v$G8_12053_out0 && v$P$CD_11034_out0;
assign v$G7_10151_out0 = v$G8_12059_out0 && v$P$CD_11040_out0;
assign v$G7_10154_out0 = v$G8_12062_out0 && v$P$CD_11043_out0;
assign v$G7_10159_out0 = v$G8_12067_out0 && v$P$CD_11048_out0;
assign v$G7_10172_out0 = v$G8_12080_out0 && v$P$CD_11061_out0;
assign v$P$CD_10932_out0 = v$P$AD_787_out0;
assign v$P$CD_11055_out0 = v$P$AD_910_out0;
assign v$END12_11274_out0 = v$G$AD_17689_out0;
assign v$END12_11277_out0 = v$G$AD_17812_out0;
assign v$END19_12218_out0 = v$P$AD_756_out0;
assign v$END19_12221_out0 = v$P$AD_879_out0;
assign v$SEL1_15991_out0 = v$IN_16199_out0[19:0];
assign v$SEL1_16001_out0 = v$IN_16201_out0[19:0];
assign v$SEL1_16022_out0 = v$IN_16205_out0[19:0];
assign v$SEL1_16032_out0 = v$IN_16207_out0[19:0];
assign v$_19274_out0 = { v$A3A_12525_out0,v$A4A_13731_out0 };
assign v$_19277_out0 = { v$A3A_12528_out0,v$A4A_13734_out0 };
assign v$G6_452_out0 = v$G4_11610_out0 || v$G7_10017_out0;
assign v$G6_457_out0 = v$G4_11615_out0 || v$G7_10022_out0;
assign v$G6_463_out0 = v$G4_11621_out0 || v$G7_10028_out0;
assign v$G6_466_out0 = v$G4_11624_out0 || v$G7_10031_out0;
assign v$G6_471_out0 = v$G4_11629_out0 || v$G7_10036_out0;
assign v$G6_484_out0 = v$G4_11642_out0 || v$G7_10049_out0;
assign v$G6_575_out0 = v$G4_11733_out0 || v$G7_10140_out0;
assign v$G6_580_out0 = v$G4_11738_out0 || v$G7_10145_out0;
assign v$G6_586_out0 = v$G4_11744_out0 || v$G7_10151_out0;
assign v$G6_589_out0 = v$G4_11747_out0 || v$G7_10154_out0;
assign v$G6_594_out0 = v$G4_11752_out0 || v$G7_10159_out0;
assign v$G6_607_out0 = v$G4_11765_out0 || v$G7_10172_out0;
assign v$_4423_out0 = { v$C2_121_out0,v$SEL1_15991_out0 };
assign v$_4433_out0 = { v$C2_131_out0,v$SEL1_16001_out0 };
assign v$_4454_out0 = { v$C2_152_out0,v$SEL1_16022_out0 };
assign v$_4464_out0 = { v$C2_162_out0,v$SEL1_16032_out0 };
assign v$G5_4695_out0 = v$G$AB_9470_out0 && v$P$CD_10912_out0;
assign v$G5_4699_out0 = v$G$AB_9474_out0 && v$P$CD_10916_out0;
assign v$G5_4718_out0 = v$G$AB_9493_out0 && v$P$CD_10935_out0;
assign v$G5_4726_out0 = v$G$AB_9501_out0 && v$P$CD_10943_out0;
assign v$G5_4728_out0 = v$G$AB_9503_out0 && v$P$CD_10945_out0;
assign v$G5_4818_out0 = v$G$AB_9593_out0 && v$P$CD_11035_out0;
assign v$G5_4822_out0 = v$G$AB_9597_out0 && v$P$CD_11039_out0;
assign v$G5_4841_out0 = v$G$AB_9616_out0 && v$P$CD_11058_out0;
assign v$G5_4849_out0 = v$G$AB_9624_out0 && v$P$CD_11066_out0;
assign v$G5_4851_out0 = v$G$AB_9626_out0 && v$P$CD_11068_out0;
assign v$G1_5766_out0 = v$P$AB_2167_out0 && v$P$CD_10909_out0;
assign v$G1_5775_out0 = v$P$AB_2176_out0 && v$P$CD_10918_out0;
assign v$G1_5776_out0 = v$P$AB_2177_out0 && v$P$CD_10919_out0;
assign v$G1_5787_out0 = v$P$AB_2188_out0 && v$P$CD_10930_out0;
assign v$G1_5789_out0 = v$P$AB_2190_out0 && v$P$CD_10932_out0;
assign v$G1_5796_out0 = v$P$AB_2197_out0 && v$P$CD_10939_out0;
assign v$G1_5797_out0 = v$P$AB_2198_out0 && v$P$CD_10940_out0;
assign v$G1_5889_out0 = v$P$AB_2290_out0 && v$P$CD_11032_out0;
assign v$G1_5898_out0 = v$P$AB_2299_out0 && v$P$CD_11041_out0;
assign v$G1_5899_out0 = v$P$AB_2300_out0 && v$P$CD_11042_out0;
assign v$G1_5910_out0 = v$P$AB_2311_out0 && v$P$CD_11053_out0;
assign v$G1_5912_out0 = v$P$AB_2313_out0 && v$P$CD_11055_out0;
assign v$G1_5919_out0 = v$P$AB_2320_out0 && v$P$CD_11062_out0;
assign v$G1_5920_out0 = v$P$AB_2321_out0 && v$P$CD_11063_out0;
assign v$_9324_out0 = { v$SEL1_9063_out0,v$C1_6259_out0 };
assign v$_9334_out0 = { v$SEL1_9073_out0,v$C1_6269_out0 };
assign v$_9355_out0 = { v$SEL1_9094_out0,v$C1_6290_out0 };
assign v$_9365_out0 = { v$SEL1_9104_out0,v$C1_6300_out0 };
assign v$_10817_out0 = { v$_14021_out0,v$_19274_out0 };
assign v$_10820_out0 = { v$_14024_out0,v$_19277_out0 };
assign v$P$AD_753_out0 = v$G1_5766_out0;
assign v$P$AD_762_out0 = v$G1_5775_out0;
assign v$P$AD_763_out0 = v$G1_5776_out0;
assign v$P$AD_774_out0 = v$G1_5787_out0;
assign v$P$AD_776_out0 = v$G1_5789_out0;
assign v$P$AD_783_out0 = v$G1_5796_out0;
assign v$P$AD_784_out0 = v$G1_5797_out0;
assign v$P$AD_876_out0 = v$G1_5889_out0;
assign v$P$AD_885_out0 = v$G1_5898_out0;
assign v$P$AD_886_out0 = v$G1_5899_out0;
assign v$P$AD_897_out0 = v$G1_5910_out0;
assign v$P$AD_899_out0 = v$G1_5912_out0;
assign v$P$AD_906_out0 = v$G1_5919_out0;
assign v$P$AD_907_out0 = v$G1_5920_out0;
assign v$MUX1_2560_out0 = v$LEFT$SHIT_3272_out0 ? v$_4423_out0 : v$_9324_out0;
assign v$MUX1_2570_out0 = v$LEFT$SHIT_3282_out0 ? v$_4433_out0 : v$_9334_out0;
assign v$MUX1_2591_out0 = v$LEFT$SHIT_3303_out0 ? v$_4454_out0 : v$_9355_out0;
assign v$MUX1_2601_out0 = v$LEFT$SHIT_3313_out0 ? v$_4464_out0 : v$_9365_out0;
assign v$COUTD_6930_out0 = v$G6_452_out0;
assign v$COUTD_6935_out0 = v$G6_457_out0;
assign v$COUTD_6941_out0 = v$G6_463_out0;
assign v$COUTD_6944_out0 = v$G6_466_out0;
assign v$COUTD_6949_out0 = v$G6_471_out0;
assign v$COUTD_6962_out0 = v$G6_484_out0;
assign v$COUTD_7053_out0 = v$G6_575_out0;
assign v$COUTD_7058_out0 = v$G6_580_out0;
assign v$COUTD_7064_out0 = v$G6_586_out0;
assign v$COUTD_7067_out0 = v$G6_589_out0;
assign v$COUTD_7072_out0 = v$G6_594_out0;
assign v$COUTD_7085_out0 = v$G6_607_out0;
assign v$G4_11616_out0 = v$G5_4695_out0 || v$G$CD_1023_out0;
assign v$G4_11620_out0 = v$G5_4699_out0 || v$G$CD_1027_out0;
assign v$G4_11639_out0 = v$G5_4718_out0 || v$G$CD_1046_out0;
assign v$G4_11647_out0 = v$G5_4726_out0 || v$G$CD_1054_out0;
assign v$G4_11649_out0 = v$G5_4728_out0 || v$G$CD_1056_out0;
assign v$G4_11739_out0 = v$G5_4818_out0 || v$G$CD_1146_out0;
assign v$G4_11743_out0 = v$G5_4822_out0 || v$G$CD_1150_out0;
assign v$G4_11762_out0 = v$G5_4841_out0 || v$G$CD_1169_out0;
assign v$G4_11770_out0 = v$G5_4849_out0 || v$G$CD_1177_out0;
assign v$G4_11772_out0 = v$G5_4851_out0 || v$G$CD_1179_out0;
assign v$C4_1413_out0 = v$COUTD_6935_out0;
assign v$C4_1416_out0 = v$COUTD_7058_out0;
assign v$P$AB_2180_out0 = v$P$AD_753_out0;
assign v$P$AB_2187_out0 = v$P$AD_753_out0;
assign v$P$AB_2191_out0 = v$P$AD_774_out0;
assign v$P$AB_2194_out0 = v$P$AD_774_out0;
assign v$P$AB_2202_out0 = v$P$AD_753_out0;
assign v$P$AB_2303_out0 = v$P$AD_876_out0;
assign v$P$AB_2310_out0 = v$P$AD_876_out0;
assign v$P$AB_2314_out0 = v$P$AD_897_out0;
assign v$P$AB_2317_out0 = v$P$AD_897_out0;
assign v$P$AB_2325_out0 = v$P$AD_876_out0;
assign v$END27_2414_out0 = v$P$AD_783_out0;
assign v$END27_2417_out0 = v$P$AD_906_out0;
assign v$END21_4504_out0 = v$P$AD_763_out0;
assign v$END21_4507_out0 = v$P$AD_886_out0;
assign v$END40_6062_out0 = v$COUTD_6949_out0;
assign v$END40_6065_out0 = v$COUTD_7072_out0;
assign v$END29_6161_out0 = v$P$AD_774_out0;
assign v$END29_6164_out0 = v$P$AD_897_out0;
assign v$CINA_8776_out0 = v$COUTD_6962_out0;
assign v$CINA_8780_out0 = v$COUTD_6962_out0;
assign v$CINA_8799_out0 = v$COUTD_6962_out0;
assign v$CINA_8807_out0 = v$COUTD_6949_out0;
assign v$CINA_8809_out0 = v$COUTD_6962_out0;
assign v$CINA_8899_out0 = v$COUTD_7085_out0;
assign v$CINA_8903_out0 = v$COUTD_7085_out0;
assign v$CINA_8922_out0 = v$COUTD_7085_out0;
assign v$CINA_8930_out0 = v$COUTD_7072_out0;
assign v$CINA_8932_out0 = v$COUTD_7085_out0;
assign v$END4_9737_out0 = v$COUTD_6930_out0;
assign v$END4_9740_out0 = v$COUTD_7053_out0;
assign v$END52_12549_out0 = v$P$AD_776_out0;
assign v$END52_12552_out0 = v$P$AD_899_out0;
assign v$END60_15741_out0 = v$COUTD_6944_out0;
assign v$END60_15744_out0 = v$COUTD_7067_out0;
assign v$MUX2_15820_out0 = v$EN_4966_out0 ? v$MUX1_2560_out0 : v$IN_16199_out0;
assign v$MUX2_15822_out0 = v$EN_4968_out0 ? v$MUX1_2570_out0 : v$IN_16201_out0;
assign v$MUX2_15826_out0 = v$EN_4972_out0 ? v$MUX1_2591_out0 : v$IN_16205_out0;
assign v$MUX2_15828_out0 = v$EN_4974_out0 ? v$MUX1_2601_out0 : v$IN_16207_out0;
assign v$C3_16323_out0 = v$COUTD_6941_out0;
assign v$C3_16326_out0 = v$COUTD_7064_out0;
assign v$C5_16519_out0 = v$COUTD_6962_out0;
assign v$C5_16522_out0 = v$COUTD_7085_out0;
assign v$END23_17336_out0 = v$P$AD_784_out0;
assign v$END23_17339_out0 = v$P$AD_907_out0;
assign v$END25_17666_out0 = v$P$AD_762_out0;
assign v$END25_17669_out0 = v$P$AD_885_out0;
assign v$G$AD_17690_out0 = v$G4_11616_out0;
assign v$G$AD_17694_out0 = v$G4_11620_out0;
assign v$G$AD_17713_out0 = v$G4_11639_out0;
assign v$G$AD_17721_out0 = v$G4_11647_out0;
assign v$G$AD_17723_out0 = v$G4_11649_out0;
assign v$G$AD_17813_out0 = v$G4_11739_out0;
assign v$G$AD_17817_out0 = v$G4_11743_out0;
assign v$G$AD_17836_out0 = v$G4_11762_out0;
assign v$G$AD_17844_out0 = v$G4_11770_out0;
assign v$G$AD_17846_out0 = v$G4_11772_out0;
assign v$END16_222_out0 = v$G$AD_17723_out0;
assign v$END16_225_out0 = v$G$AD_17846_out0;
assign v$END14_284_out0 = v$G$AD_17694_out0;
assign v$END14_287_out0 = v$G$AD_17817_out0;
assign v$G$CD_1043_out0 = v$G$AD_17721_out0;
assign v$G$CD_1166_out0 = v$G$AD_17844_out0;
assign {v$A7A_1815_out1,v$A7A_1815_out0 } = v$A5_6901_out0 + v$B5_18978_out0 + v$C4_1413_out0;
assign {v$A7A_1818_out1,v$A7A_1818_out0 } = v$A5_6904_out0 + v$B5_18981_out0 + v$C4_1416_out0;
assign v$C4_2038_out0 = v$C4_1413_out0;
assign v$C4_2041_out0 = v$C4_1416_out0;
assign {v$A6A_3334_out1,v$A6A_3334_out0 } = v$A6_320_out0 + v$B6_13883_out0 + v$C5_16519_out0;
assign {v$A6A_3337_out1,v$A6A_3337_out0 } = v$A6_323_out0 + v$B6_13886_out0 + v$C5_16522_out0;
assign v$G1_5779_out0 = v$P$AB_2180_out0 && v$P$CD_10922_out0;
assign v$G1_5786_out0 = v$P$AB_2187_out0 && v$P$CD_10929_out0;
assign v$G1_5790_out0 = v$P$AB_2191_out0 && v$P$CD_10933_out0;
assign v$G1_5793_out0 = v$P$AB_2194_out0 && v$P$CD_10936_out0;
assign v$G1_5801_out0 = v$P$AB_2202_out0 && v$P$CD_10944_out0;
assign v$G1_5902_out0 = v$P$AB_2303_out0 && v$P$CD_11045_out0;
assign v$G1_5909_out0 = v$P$AB_2310_out0 && v$P$CD_11052_out0;
assign v$G1_5913_out0 = v$P$AB_2314_out0 && v$P$CD_11056_out0;
assign v$G1_5916_out0 = v$P$AB_2317_out0 && v$P$CD_11059_out0;
assign v$G1_5924_out0 = v$P$AB_2325_out0 && v$P$CD_11067_out0;
assign v$G$AB_9467_out0 = v$G$AD_17713_out0;
assign v$G$AB_9476_out0 = v$G$AD_17713_out0;
assign v$G$AB_9477_out0 = v$G$AD_17690_out0;
assign v$G$AB_9488_out0 = v$G$AD_17713_out0;
assign v$G$AB_9490_out0 = v$G$AD_17713_out0;
assign v$G$AB_9497_out0 = v$G$AD_17713_out0;
assign v$G$AB_9498_out0 = v$G$AD_17690_out0;
assign v$G$AB_9590_out0 = v$G$AD_17836_out0;
assign v$G$AB_9599_out0 = v$G$AD_17836_out0;
assign v$G$AB_9600_out0 = v$G$AD_17813_out0;
assign v$G$AB_9611_out0 = v$G$AD_17836_out0;
assign v$G$AB_9613_out0 = v$G$AD_17836_out0;
assign v$G$AB_9620_out0 = v$G$AD_17836_out0;
assign v$G$AB_9621_out0 = v$G$AD_17813_out0;
assign v$G8_11931_out0 = v$CINA_8776_out0 && v$P$AB_2170_out0;
assign v$G8_11935_out0 = v$CINA_8780_out0 && v$P$AB_2174_out0;
assign v$G8_11954_out0 = v$CINA_8799_out0 && v$P$AB_2193_out0;
assign v$G8_11962_out0 = v$CINA_8807_out0 && v$P$AB_2201_out0;
assign v$G8_11964_out0 = v$CINA_8809_out0 && v$P$AB_2203_out0;
assign v$G8_12054_out0 = v$CINA_8899_out0 && v$P$AB_2293_out0;
assign v$G8_12058_out0 = v$CINA_8903_out0 && v$P$AB_2297_out0;
assign v$G8_12077_out0 = v$CINA_8922_out0 && v$P$AB_2316_out0;
assign v$G8_12085_out0 = v$CINA_8930_out0 && v$P$AB_2324_out0;
assign v$G8_12087_out0 = v$CINA_8932_out0 && v$P$AB_2326_out0;
assign v$C5_12253_out0 = v$C5_16519_out0;
assign v$C5_12256_out0 = v$C5_16522_out0;
assign v$END18_12519_out0 = v$G$AD_17690_out0;
assign v$END18_12522_out0 = v$G$AD_17813_out0;
assign v$OUT_15532_out0 = v$MUX2_15820_out0;
assign v$OUT_15542_out0 = v$MUX2_15822_out0;
assign v$OUT_15563_out0 = v$MUX2_15826_out0;
assign v$OUT_15573_out0 = v$MUX2_15828_out0;
assign v$C3_16420_out0 = v$C3_16323_out0;
assign v$C3_16423_out0 = v$C3_16326_out0;
assign {v$A5A_16709_out1,v$A5A_16709_out0 } = v$A4_18138_out0 + v$B4_15266_out0 + v$C3_16323_out0;
assign {v$A5A_16712_out1,v$A5A_16712_out0 } = v$A4_18141_out0 + v$B4_15269_out0 + v$C3_16326_out0;
assign v$_82_out0 = { v$A5A_16709_out0,v$A7A_1815_out0 };
assign v$_85_out0 = { v$A5A_16712_out0,v$A7A_1818_out0 };
assign v$P$AD_766_out0 = v$G1_5779_out0;
assign v$P$AD_773_out0 = v$G1_5786_out0;
assign v$P$AD_777_out0 = v$G1_5790_out0;
assign v$P$AD_780_out0 = v$G1_5793_out0;
assign v$P$AD_788_out0 = v$G1_5801_out0;
assign v$P$AD_889_out0 = v$G1_5902_out0;
assign v$P$AD_896_out0 = v$G1_5909_out0;
assign v$P$AD_900_out0 = v$G1_5913_out0;
assign v$P$AD_903_out0 = v$G1_5916_out0;
assign v$P$AD_911_out0 = v$G1_5924_out0;
assign v$_2646_out0 = { v$C4_2038_out0,v$C5_12253_out0 };
assign v$_2649_out0 = { v$C4_2041_out0,v$C5_12256_out0 };
assign v$END5_4301_out0 = v$A7A_1815_out1;
assign v$END5_4304_out0 = v$A7A_1818_out1;
assign v$G5_4692_out0 = v$G$AB_9467_out0 && v$P$CD_10909_out0;
assign v$G5_4701_out0 = v$G$AB_9476_out0 && v$P$CD_10918_out0;
assign v$G5_4702_out0 = v$G$AB_9477_out0 && v$P$CD_10919_out0;
assign v$G5_4713_out0 = v$G$AB_9488_out0 && v$P$CD_10930_out0;
assign v$G5_4715_out0 = v$G$AB_9490_out0 && v$P$CD_10932_out0;
assign v$G5_4722_out0 = v$G$AB_9497_out0 && v$P$CD_10939_out0;
assign v$G5_4723_out0 = v$G$AB_9498_out0 && v$P$CD_10940_out0;
assign v$G5_4815_out0 = v$G$AB_9590_out0 && v$P$CD_11032_out0;
assign v$G5_4824_out0 = v$G$AB_9599_out0 && v$P$CD_11041_out0;
assign v$G5_4825_out0 = v$G$AB_9600_out0 && v$P$CD_11042_out0;
assign v$G5_4836_out0 = v$G$AB_9611_out0 && v$P$CD_11053_out0;
assign v$G5_4838_out0 = v$G$AB_9613_out0 && v$P$CD_11055_out0;
assign v$G5_4845_out0 = v$G$AB_9620_out0 && v$P$CD_11062_out0;
assign v$G5_4846_out0 = v$G$AB_9621_out0 && v$P$CD_11063_out0;
assign v$IN_5381_out0 = v$OUT_15532_out0;
assign v$IN_5391_out0 = v$OUT_15542_out0;
assign v$IN_5412_out0 = v$OUT_15563_out0;
assign v$IN_5422_out0 = v$OUT_15573_out0;
assign v$END4_5463_out0 = v$A5A_16709_out1;
assign v$END4_5466_out0 = v$A5A_16712_out1;
assign v$G7_10023_out0 = v$G8_11931_out0 && v$P$CD_10912_out0;
assign v$G7_10027_out0 = v$G8_11935_out0 && v$P$CD_10916_out0;
assign v$G7_10046_out0 = v$G8_11954_out0 && v$P$CD_10935_out0;
assign v$G7_10054_out0 = v$G8_11962_out0 && v$P$CD_10943_out0;
assign v$G7_10056_out0 = v$G8_11964_out0 && v$P$CD_10945_out0;
assign v$G7_10146_out0 = v$G8_12054_out0 && v$P$CD_11035_out0;
assign v$G7_10150_out0 = v$G8_12058_out0 && v$P$CD_11039_out0;
assign v$G7_10169_out0 = v$G8_12077_out0 && v$P$CD_11058_out0;
assign v$G7_10177_out0 = v$G8_12085_out0 && v$P$CD_11066_out0;
assign v$G7_10179_out0 = v$G8_12087_out0 && v$P$CD_11068_out0;
assign v$_15614_out0 = { v$C2_18777_out0,v$C3_16420_out0 };
assign v$_15617_out0 = { v$C2_18780_out0,v$C3_16423_out0 };
assign v$END6_15831_out0 = v$A6A_3334_out1;
assign v$END6_15834_out0 = v$A6A_3337_out1;
assign v$END33_273_out0 = v$P$AD_780_out0;
assign v$END33_276_out0 = v$P$AD_903_out0;
assign v$G6_458_out0 = v$G4_11616_out0 || v$G7_10023_out0;
assign v$G6_462_out0 = v$G4_11620_out0 || v$G7_10027_out0;
assign v$G6_481_out0 = v$G4_11639_out0 || v$G7_10046_out0;
assign v$G6_489_out0 = v$G4_11647_out0 || v$G7_10054_out0;
assign v$G6_491_out0 = v$G4_11649_out0 || v$G7_10056_out0;
assign v$G6_581_out0 = v$G4_11739_out0 || v$G7_10146_out0;
assign v$G6_585_out0 = v$G4_11743_out0 || v$G7_10150_out0;
assign v$G6_604_out0 = v$G4_11762_out0 || v$G7_10169_out0;
assign v$G6_612_out0 = v$G4_11770_out0 || v$G7_10177_out0;
assign v$G6_614_out0 = v$G4_11772_out0 || v$G7_10179_out0;
assign v$P$AB_2173_out0 = v$P$AD_773_out0;
assign v$P$AB_2192_out0 = v$P$AD_773_out0;
assign v$P$AB_2296_out0 = v$P$AD_896_out0;
assign v$P$AB_2315_out0 = v$P$AD_896_out0;
assign v$END47_2876_out0 = v$P$AD_773_out0;
assign v$END47_2879_out0 = v$P$AD_896_out0;
assign v$IN_5239_out0 = v$IN_5381_out0;
assign v$IN_5242_out0 = v$IN_5391_out0;
assign v$IN_5249_out0 = v$IN_5412_out0;
assign v$IN_5252_out0 = v$IN_5422_out0;
assign v$_7568_out0 = { v$_9235_out0,v$_15614_out0 };
assign v$_7571_out0 = { v$_9238_out0,v$_15617_out0 };
assign v$G4_11613_out0 = v$G5_4692_out0 || v$G$CD_1020_out0;
assign v$G4_11622_out0 = v$G5_4701_out0 || v$G$CD_1029_out0;
assign v$G4_11623_out0 = v$G5_4702_out0 || v$G$CD_1030_out0;
assign v$G4_11634_out0 = v$G5_4713_out0 || v$G$CD_1041_out0;
assign v$G4_11636_out0 = v$G5_4715_out0 || v$G$CD_1043_out0;
assign v$G4_11643_out0 = v$G5_4722_out0 || v$G$CD_1050_out0;
assign v$G4_11644_out0 = v$G5_4723_out0 || v$G$CD_1051_out0;
assign v$G4_11736_out0 = v$G5_4815_out0 || v$G$CD_1143_out0;
assign v$G4_11745_out0 = v$G5_4824_out0 || v$G$CD_1152_out0;
assign v$G4_11746_out0 = v$G5_4825_out0 || v$G$CD_1153_out0;
assign v$G4_11757_out0 = v$G5_4836_out0 || v$G$CD_1164_out0;
assign v$G4_11759_out0 = v$G5_4838_out0 || v$G$CD_1166_out0;
assign v$G4_11766_out0 = v$G5_4845_out0 || v$G$CD_1173_out0;
assign v$G4_11767_out0 = v$G5_4846_out0 || v$G$CD_1174_out0;
assign v$END44_16258_out0 = v$P$AD_788_out0;
assign v$END44_16261_out0 = v$P$AD_911_out0;
assign v$END42_18916_out0 = v$P$AD_766_out0;
assign v$END42_18919_out0 = v$P$AD_889_out0;
assign v$END31_19131_out0 = v$P$AD_777_out0;
assign v$END31_19134_out0 = v$P$AD_900_out0;
assign v$G1_5772_out0 = v$P$AB_2173_out0 && v$P$CD_10915_out0;
assign v$G1_5791_out0 = v$P$AB_2192_out0 && v$P$CD_10934_out0;
assign v$G1_5895_out0 = v$P$AB_2296_out0 && v$P$CD_11038_out0;
assign v$G1_5914_out0 = v$P$AB_2315_out0 && v$P$CD_11057_out0;
assign v$COUTD_6936_out0 = v$G6_458_out0;
assign v$COUTD_6940_out0 = v$G6_462_out0;
assign v$COUTD_6959_out0 = v$G6_481_out0;
assign v$COUTD_6967_out0 = v$G6_489_out0;
assign v$COUTD_6969_out0 = v$G6_491_out0;
assign v$COUTD_7059_out0 = v$G6_581_out0;
assign v$COUTD_7063_out0 = v$G6_585_out0;
assign v$COUTD_7082_out0 = v$G6_604_out0;
assign v$COUTD_7090_out0 = v$G6_612_out0;
assign v$COUTD_7092_out0 = v$G6_614_out0;
assign v$SEL1_9062_out0 = v$IN_5239_out0[23:8];
assign v$SEL1_9072_out0 = v$IN_5242_out0[23:8];
assign v$SEL1_9093_out0 = v$IN_5249_out0[23:8];
assign v$SEL1_9103_out0 = v$IN_5252_out0[23:8];
assign v$SEL1_15990_out0 = v$IN_5239_out0[15:0];
assign v$SEL1_16000_out0 = v$IN_5242_out0[15:0];
assign v$SEL1_16021_out0 = v$IN_5249_out0[15:0];
assign v$SEL1_16031_out0 = v$IN_5252_out0[15:0];
assign v$G$AD_17687_out0 = v$G4_11613_out0;
assign v$G$AD_17696_out0 = v$G4_11622_out0;
assign v$G$AD_17697_out0 = v$G4_11623_out0;
assign v$G$AD_17708_out0 = v$G4_11634_out0;
assign v$G$AD_17710_out0 = v$G4_11636_out0;
assign v$G$AD_17717_out0 = v$G4_11643_out0;
assign v$G$AD_17718_out0 = v$G4_11644_out0;
assign v$G$AD_17810_out0 = v$G4_11736_out0;
assign v$G$AD_17819_out0 = v$G4_11745_out0;
assign v$G$AD_17820_out0 = v$G4_11746_out0;
assign v$G$AD_17831_out0 = v$G4_11757_out0;
assign v$G$AD_17833_out0 = v$G4_11759_out0;
assign v$G$AD_17840_out0 = v$G4_11766_out0;
assign v$G$AD_17841_out0 = v$G4_11767_out0;
assign v$END53_330_out0 = v$G$AD_17710_out0;
assign v$END53_333_out0 = v$G$AD_17833_out0;
assign v$P$AD_759_out0 = v$G1_5772_out0;
assign v$P$AD_778_out0 = v$G1_5791_out0;
assign v$P$AD_882_out0 = v$G1_5895_out0;
assign v$P$AD_901_out0 = v$G1_5914_out0;
assign v$_4422_out0 = { v$C2_120_out0,v$SEL1_15990_out0 };
assign v$_4432_out0 = { v$C2_130_out0,v$SEL1_16000_out0 };
assign v$_4453_out0 = { v$C2_151_out0,v$SEL1_16021_out0 };
assign v$_4463_out0 = { v$C2_161_out0,v$SEL1_16031_out0 };
assign v$END26_6678_out0 = v$G$AD_17717_out0;
assign v$END26_6681_out0 = v$G$AD_17840_out0;
assign v$C8_7748_out0 = v$COUTD_6936_out0;
assign v$C8_7751_out0 = v$COUTD_7059_out0;
assign v$CINA_8773_out0 = v$COUTD_6959_out0;
assign v$CINA_8782_out0 = v$COUTD_6959_out0;
assign v$CINA_8783_out0 = v$COUTD_6936_out0;
assign v$CINA_8794_out0 = v$COUTD_6959_out0;
assign v$CINA_8796_out0 = v$COUTD_6959_out0;
assign v$CINA_8803_out0 = v$COUTD_6959_out0;
assign v$CINA_8804_out0 = v$COUTD_6936_out0;
assign v$CINA_8896_out0 = v$COUTD_7082_out0;
assign v$CINA_8905_out0 = v$COUTD_7082_out0;
assign v$CINA_8906_out0 = v$COUTD_7059_out0;
assign v$CINA_8917_out0 = v$COUTD_7082_out0;
assign v$CINA_8919_out0 = v$COUTD_7082_out0;
assign v$CINA_8926_out0 = v$COUTD_7082_out0;
assign v$CINA_8927_out0 = v$COUTD_7059_out0;
assign v$_9323_out0 = { v$SEL1_9062_out0,v$C1_6258_out0 };
assign v$_9333_out0 = { v$SEL1_9072_out0,v$C1_6268_out0 };
assign v$_9354_out0 = { v$SEL1_9093_out0,v$C1_6289_out0 };
assign v$_9364_out0 = { v$SEL1_9103_out0,v$C1_6299_out0 };
assign v$G$AB_9480_out0 = v$G$AD_17687_out0;
assign v$G$AB_9487_out0 = v$G$AD_17687_out0;
assign v$G$AB_9491_out0 = v$G$AD_17708_out0;
assign v$G$AB_9494_out0 = v$G$AD_17708_out0;
assign v$G$AB_9502_out0 = v$G$AD_17687_out0;
assign v$G$AB_9603_out0 = v$G$AD_17810_out0;
assign v$G$AB_9610_out0 = v$G$AD_17810_out0;
assign v$G$AB_9614_out0 = v$G$AD_17831_out0;
assign v$G$AB_9617_out0 = v$G$AD_17831_out0;
assign v$G$AB_9625_out0 = v$G$AD_17810_out0;
assign v$C6_9966_out0 = v$COUTD_6940_out0;
assign v$C6_9969_out0 = v$COUTD_7063_out0;
assign v$C7_11475_out0 = v$COUTD_6969_out0;
assign v$C7_11478_out0 = v$COUTD_7092_out0;
assign v$END20_13847_out0 = v$G$AD_17697_out0;
assign v$END20_13850_out0 = v$G$AD_17820_out0;
assign v$END28_14248_out0 = v$G$AD_17708_out0;
assign v$END28_14251_out0 = v$G$AD_17831_out0;
assign v$C11_15404_out0 = v$COUTD_6959_out0;
assign v$C11_15407_out0 = v$COUTD_7082_out0;
assign v$END22_16073_out0 = v$G$AD_17718_out0;
assign v$END22_16076_out0 = v$G$AD_17841_out0;
assign v$END24_17022_out0 = v$G$AD_17696_out0;
assign v$END24_17025_out0 = v$G$AD_17819_out0;
assign v$END61_18570_out0 = v$COUTD_6967_out0;
assign v$END61_18573_out0 = v$COUTD_7090_out0;
assign {v$A8A_1659_out1,v$A8A_1659_out0 } = v$A7_15891_out0 + v$B7_17634_out0 + v$C6_9966_out0;
assign {v$A8A_1662_out1,v$A8A_1662_out0 } = v$A7_15894_out0 + v$B7_17637_out0 + v$C6_9969_out0;
assign v$MUX1_2559_out0 = v$LEFT$SHIT_3271_out0 ? v$_4422_out0 : v$_9323_out0;
assign v$MUX1_2569_out0 = v$LEFT$SHIT_3281_out0 ? v$_4432_out0 : v$_9333_out0;
assign v$MUX1_2590_out0 = v$LEFT$SHIT_3302_out0 ? v$_4453_out0 : v$_9354_out0;
assign v$MUX1_2600_out0 = v$LEFT$SHIT_3312_out0 ? v$_4463_out0 : v$_9364_out0;
assign {v$A17A_2682_out1,v$A17A_2682_out0 } = v$A12_3355_out0 + v$B12_2114_out0 + v$C11_15404_out0;
assign {v$A17A_2685_out1,v$A17A_2685_out0 } = v$A12_3358_out0 + v$B12_2117_out0 + v$C11_15407_out0;
assign v$G5_4705_out0 = v$G$AB_9480_out0 && v$P$CD_10922_out0;
assign v$G5_4712_out0 = v$G$AB_9487_out0 && v$P$CD_10929_out0;
assign v$G5_4716_out0 = v$G$AB_9491_out0 && v$P$CD_10933_out0;
assign v$G5_4719_out0 = v$G$AB_9494_out0 && v$P$CD_10936_out0;
assign v$G5_4727_out0 = v$G$AB_9502_out0 && v$P$CD_10944_out0;
assign v$G5_4828_out0 = v$G$AB_9603_out0 && v$P$CD_11045_out0;
assign v$G5_4835_out0 = v$G$AB_9610_out0 && v$P$CD_11052_out0;
assign v$G5_4839_out0 = v$G$AB_9614_out0 && v$P$CD_11056_out0;
assign v$G5_4842_out0 = v$G$AB_9617_out0 && v$P$CD_11059_out0;
assign v$G5_4850_out0 = v$G$AB_9625_out0 && v$P$CD_11067_out0;
assign v$C6_7341_out0 = v$C6_9966_out0;
assign v$C6_7344_out0 = v$C6_9969_out0;
assign v$C11_9887_out0 = v$C11_15404_out0;
assign v$C11_9890_out0 = v$C11_15407_out0;
assign {v$A9A_10862_out1,v$A9A_10862_out0 } = v$A8_18697_out0 + v$B8_13715_out0 + v$C7_11475_out0;
assign {v$A9A_10865_out1,v$A9A_10865_out0 } = v$A8_18700_out0 + v$B8_13718_out0 + v$C7_11478_out0;
assign v$G8_11928_out0 = v$CINA_8773_out0 && v$P$AB_2167_out0;
assign v$G8_11937_out0 = v$CINA_8782_out0 && v$P$AB_2176_out0;
assign v$G8_11938_out0 = v$CINA_8783_out0 && v$P$AB_2177_out0;
assign v$G8_11949_out0 = v$CINA_8794_out0 && v$P$AB_2188_out0;
assign v$G8_11951_out0 = v$CINA_8796_out0 && v$P$AB_2190_out0;
assign v$G8_11958_out0 = v$CINA_8803_out0 && v$P$AB_2197_out0;
assign v$G8_11959_out0 = v$CINA_8804_out0 && v$P$AB_2198_out0;
assign v$G8_12051_out0 = v$CINA_8896_out0 && v$P$AB_2290_out0;
assign v$G8_12060_out0 = v$CINA_8905_out0 && v$P$AB_2299_out0;
assign v$G8_12061_out0 = v$CINA_8906_out0 && v$P$AB_2300_out0;
assign v$G8_12072_out0 = v$CINA_8917_out0 && v$P$AB_2311_out0;
assign v$G8_12074_out0 = v$CINA_8919_out0 && v$P$AB_2313_out0;
assign v$G8_12081_out0 = v$CINA_8926_out0 && v$P$AB_2320_out0;
assign v$G8_12082_out0 = v$CINA_8927_out0 && v$P$AB_2321_out0;
assign v$END51_12242_out0 = v$P$AD_759_out0;
assign v$END51_12245_out0 = v$P$AD_882_out0;
assign {v$A10A_16612_out1,v$A10A_16612_out0 } = v$A9_3643_out0 + v$B9_4220_out0 + v$C8_7748_out0;
assign {v$A10A_16615_out1,v$A10A_16615_out0 } = v$A9_3646_out0 + v$B9_4223_out0 + v$C8_7751_out0;
assign v$C7_17051_out0 = v$C7_11475_out0;
assign v$C7_17054_out0 = v$C7_11478_out0;
assign v$END49_19059_out0 = v$P$AD_778_out0;
assign v$END49_19062_out0 = v$P$AD_901_out0;
assign v$C8_19107_out0 = v$C8_7748_out0;
assign v$C8_19110_out0 = v$C8_7751_out0;
assign v$MUX2_2694_out0 = v$EN_1499_out0 ? v$MUX1_2559_out0 : v$IN_5239_out0;
assign v$MUX2_2697_out0 = v$EN_1502_out0 ? v$MUX1_2569_out0 : v$IN_5242_out0;
assign v$MUX2_2704_out0 = v$EN_1509_out0 ? v$MUX1_2590_out0 : v$IN_5249_out0;
assign v$MUX2_2707_out0 = v$EN_1512_out0 ? v$MUX1_2600_out0 : v$IN_5252_out0;
assign v$END7_3582_out0 = v$A8A_1659_out1;
assign v$END7_3585_out0 = v$A8A_1662_out1;
assign v$_3826_out0 = { v$A6A_3334_out0,v$A8A_1659_out0 };
assign v$_3829_out0 = { v$A6A_3337_out0,v$A8A_1662_out0 };
assign v$END8_4070_out0 = v$A9A_10862_out1;
assign v$END8_4073_out0 = v$A9A_10865_out1;
assign v$END9_4392_out0 = v$A10A_16612_out1;
assign v$END9_4395_out0 = v$A10A_16615_out1;
assign v$ENDw_9930_out0 = v$A17A_2682_out1;
assign v$ENDw_9933_out0 = v$A17A_2685_out1;
assign v$G7_10020_out0 = v$G8_11928_out0 && v$P$CD_10909_out0;
assign v$G7_10029_out0 = v$G8_11937_out0 && v$P$CD_10918_out0;
assign v$G7_10030_out0 = v$G8_11938_out0 && v$P$CD_10919_out0;
assign v$G7_10041_out0 = v$G8_11949_out0 && v$P$CD_10930_out0;
assign v$G7_10043_out0 = v$G8_11951_out0 && v$P$CD_10932_out0;
assign v$G7_10050_out0 = v$G8_11958_out0 && v$P$CD_10939_out0;
assign v$G7_10051_out0 = v$G8_11959_out0 && v$P$CD_10940_out0;
assign v$G7_10143_out0 = v$G8_12051_out0 && v$P$CD_11032_out0;
assign v$G7_10152_out0 = v$G8_12060_out0 && v$P$CD_11041_out0;
assign v$G7_10153_out0 = v$G8_12061_out0 && v$P$CD_11042_out0;
assign v$G7_10164_out0 = v$G8_12072_out0 && v$P$CD_11053_out0;
assign v$G7_10166_out0 = v$G8_12074_out0 && v$P$CD_11055_out0;
assign v$G7_10173_out0 = v$G8_12081_out0 && v$P$CD_11062_out0;
assign v$G7_10174_out0 = v$G8_12082_out0 && v$P$CD_11063_out0;
assign v$G4_11626_out0 = v$G5_4705_out0 || v$G$CD_1033_out0;
assign v$G4_11633_out0 = v$G5_4712_out0 || v$G$CD_1040_out0;
assign v$G4_11637_out0 = v$G5_4716_out0 || v$G$CD_1044_out0;
assign v$G4_11640_out0 = v$G5_4719_out0 || v$G$CD_1047_out0;
assign v$G4_11648_out0 = v$G5_4727_out0 || v$G$CD_1055_out0;
assign v$G4_11749_out0 = v$G5_4828_out0 || v$G$CD_1156_out0;
assign v$G4_11756_out0 = v$G5_4835_out0 || v$G$CD_1163_out0;
assign v$G4_11760_out0 = v$G5_4839_out0 || v$G$CD_1167_out0;
assign v$G4_11763_out0 = v$G5_4842_out0 || v$G$CD_1170_out0;
assign v$G4_11771_out0 = v$G5_4850_out0 || v$G$CD_1178_out0;
assign v$_15630_out0 = { v$A9A_10862_out0,v$A10A_16612_out0 };
assign v$_15633_out0 = { v$A9A_10865_out0,v$A10A_16615_out0 };
assign v$_16924_out0 = { v$C6_7341_out0,v$C7_17051_out0 };
assign v$_16927_out0 = { v$C6_7344_out0,v$C7_17054_out0 };
assign v$G6_455_out0 = v$G4_11613_out0 || v$G7_10020_out0;
assign v$G6_464_out0 = v$G4_11622_out0 || v$G7_10029_out0;
assign v$G6_465_out0 = v$G4_11623_out0 || v$G7_10030_out0;
assign v$G6_476_out0 = v$G4_11634_out0 || v$G7_10041_out0;
assign v$G6_478_out0 = v$G4_11636_out0 || v$G7_10043_out0;
assign v$G6_485_out0 = v$G4_11643_out0 || v$G7_10050_out0;
assign v$G6_486_out0 = v$G4_11644_out0 || v$G7_10051_out0;
assign v$G6_578_out0 = v$G4_11736_out0 || v$G7_10143_out0;
assign v$G6_587_out0 = v$G4_11745_out0 || v$G7_10152_out0;
assign v$G6_588_out0 = v$G4_11746_out0 || v$G7_10153_out0;
assign v$G6_599_out0 = v$G4_11757_out0 || v$G7_10164_out0;
assign v$G6_601_out0 = v$G4_11759_out0 || v$G7_10166_out0;
assign v$G6_608_out0 = v$G4_11766_out0 || v$G7_10173_out0;
assign v$G6_609_out0 = v$G4_11767_out0 || v$G7_10174_out0;
assign v$_7719_out0 = { v$_2646_out0,v$_16924_out0 };
assign v$_7722_out0 = { v$_2649_out0,v$_16927_out0 };
assign v$OUT_15531_out0 = v$MUX2_2694_out0;
assign v$OUT_15541_out0 = v$MUX2_2697_out0;
assign v$OUT_15562_out0 = v$MUX2_2704_out0;
assign v$OUT_15572_out0 = v$MUX2_2707_out0;
assign v$G$AD_17700_out0 = v$G4_11626_out0;
assign v$G$AD_17707_out0 = v$G4_11633_out0;
assign v$G$AD_17711_out0 = v$G4_11637_out0;
assign v$G$AD_17714_out0 = v$G4_11640_out0;
assign v$G$AD_17722_out0 = v$G4_11648_out0;
assign v$G$AD_17823_out0 = v$G4_11749_out0;
assign v$G$AD_17830_out0 = v$G4_11756_out0;
assign v$G$AD_17834_out0 = v$G4_11760_out0;
assign v$G$AD_17837_out0 = v$G4_11763_out0;
assign v$G$AD_17845_out0 = v$G4_11771_out0;
assign v$_18579_out0 = { v$_82_out0,v$_3826_out0 };
assign v$_18582_out0 = { v$_85_out0,v$_3829_out0 };
assign v$END32_2664_out0 = v$G$AD_17714_out0;
assign v$END32_2667_out0 = v$G$AD_17837_out0;
assign v$IN_5383_out0 = v$OUT_15531_out0;
assign v$IN_5393_out0 = v$OUT_15541_out0;
assign v$IN_5414_out0 = v$OUT_15562_out0;
assign v$IN_5424_out0 = v$OUT_15572_out0;
assign v$COUTD_6933_out0 = v$G6_455_out0;
assign v$COUTD_6942_out0 = v$G6_464_out0;
assign v$COUTD_6943_out0 = v$G6_465_out0;
assign v$COUTD_6954_out0 = v$G6_476_out0;
assign v$COUTD_6956_out0 = v$G6_478_out0;
assign v$COUTD_6963_out0 = v$G6_485_out0;
assign v$COUTD_6964_out0 = v$G6_486_out0;
assign v$COUTD_7056_out0 = v$G6_578_out0;
assign v$COUTD_7065_out0 = v$G6_587_out0;
assign v$COUTD_7066_out0 = v$G6_588_out0;
assign v$COUTD_7077_out0 = v$G6_599_out0;
assign v$COUTD_7079_out0 = v$G6_601_out0;
assign v$COUTD_7086_out0 = v$G6_608_out0;
assign v$COUTD_7087_out0 = v$G6_609_out0;
assign v$_8112_out0 = { v$_7568_out0,v$_7719_out0 };
assign v$_8115_out0 = { v$_7571_out0,v$_7722_out0 };
assign v$G$AB_9473_out0 = v$G$AD_17707_out0;
assign v$G$AB_9492_out0 = v$G$AD_17707_out0;
assign v$G$AB_9596_out0 = v$G$AD_17830_out0;
assign v$G$AB_9615_out0 = v$G$AD_17830_out0;
assign v$END43_13771_out0 = v$G$AD_17722_out0;
assign v$END43_13774_out0 = v$G$AD_17845_out0;
assign v$END46_15663_out0 = v$G$AD_17707_out0;
assign v$END46_15666_out0 = v$G$AD_17830_out0;
assign v$END30_16309_out0 = v$G$AD_17711_out0;
assign v$END30_16312_out0 = v$G$AD_17834_out0;
assign v$END41_17286_out0 = v$G$AD_17700_out0;
assign v$END41_17289_out0 = v$G$AD_17823_out0;
assign v$_18358_out0 = { v$_10817_out0,v$_18579_out0 };
assign v$_18361_out0 = { v$_10820_out0,v$_18582_out0 };
assign v$C14_290_out0 = v$COUTD_6954_out0;
assign v$C14_293_out0 = v$COUTD_7077_out0;
assign v$C17_2716_out0 = v$COUTD_6933_out0;
assign v$C17_2719_out0 = v$COUTD_7056_out0;
assign v$IN_4040_out0 = v$IN_5383_out0;
assign v$IN_4043_out0 = v$IN_5393_out0;
assign v$IN_4049_out0 = v$IN_5414_out0;
assign v$IN_4052_out0 = v$IN_5424_out0;
assign v$G5_4698_out0 = v$G$AB_9473_out0 && v$P$CD_10915_out0;
assign v$G5_4717_out0 = v$G$AB_9492_out0 && v$P$CD_10934_out0;
assign v$G5_4821_out0 = v$G$AB_9596_out0 && v$P$CD_11038_out0;
assign v$G5_4840_out0 = v$G$AB_9615_out0 && v$P$CD_11057_out0;
assign v$C23_5056_out0 = v$COUTD_6956_out0;
assign v$C23_5059_out0 = v$COUTD_7079_out0;
assign v$C9_6216_out0 = v$COUTD_6943_out0;
assign v$C9_6219_out0 = v$COUTD_7066_out0;
assign v$CINA_8786_out0 = v$COUTD_6933_out0;
assign v$CINA_8793_out0 = v$COUTD_6933_out0;
assign v$CINA_8797_out0 = v$COUTD_6954_out0;
assign v$CINA_8800_out0 = v$COUTD_6954_out0;
assign v$CINA_8808_out0 = v$COUTD_6933_out0;
assign v$CINA_8909_out0 = v$COUTD_7056_out0;
assign v$CINA_8916_out0 = v$COUTD_7056_out0;
assign v$CINA_8920_out0 = v$COUTD_7077_out0;
assign v$CINA_8923_out0 = v$COUTD_7077_out0;
assign v$CINA_8931_out0 = v$COUTD_7056_out0;
assign v$C13_12346_out0 = v$COUTD_6963_out0;
assign v$C13_12349_out0 = v$COUTD_7086_out0;
assign v$C10_13301_out0 = v$COUTD_6964_out0;
assign v$C10_13304_out0 = v$COUTD_7087_out0;
assign v$C12_14094_out0 = v$COUTD_6942_out0;
assign v$C12_14097_out0 = v$COUTD_7065_out0;
assign v$C14_340_out0 = v$C14_290_out0;
assign v$C14_343_out0 = v$C14_293_out0;
assign v$C10_2103_out0 = v$C10_13301_out0;
assign v$C10_2106_out0 = v$C10_13304_out0;
assign {v$A12A_4613_out1,v$A12A_4613_out0 } = v$A11_10386_out0 + v$B11_9443_out0 + v$C10_13301_out0;
assign {v$A12A_4616_out1,v$A12A_4616_out0 } = v$A11_10389_out0 + v$B11_9446_out0 + v$C10_13304_out0;
assign v$C17_6342_out0 = v$C17_2716_out0;
assign v$C17_6345_out0 = v$C17_2719_out0;
assign {v$A13_7554_out1,v$A13_7554_out0 } = v$A15_17957_out0 + v$B15_10446_out0 + v$C14_290_out0;
assign {v$A13_7557_out1,v$A13_7557_out0 } = v$A15_17960_out0 + v$B15_10449_out0 + v$C14_293_out0;
assign v$SEL1_9064_out0 = v$IN_4040_out0[23:16];
assign v$SEL1_9074_out0 = v$IN_4043_out0[23:16];
assign v$SEL1_9095_out0 = v$IN_4049_out0[23:16];
assign v$SEL1_9105_out0 = v$IN_4052_out0[23:16];
assign v$C12_9767_out0 = v$C12_14094_out0;
assign v$C12_9770_out0 = v$C12_14097_out0;
assign {v$A18_10458_out1,v$A18_10458_out0 } = v$A13_14445_out0 + v$B13_9022_out0 + v$C12_14094_out0;
assign {v$A18_10461_out1,v$A18_10461_out0 } = v$A13_14448_out0 + v$B13_9025_out0 + v$C12_14097_out0;
assign v$G4_11619_out0 = v$G5_4698_out0 || v$G$CD_1026_out0;
assign v$G4_11638_out0 = v$G5_4717_out0 || v$G$CD_1045_out0;
assign v$G4_11742_out0 = v$G5_4821_out0 || v$G$CD_1149_out0;
assign v$G4_11761_out0 = v$G5_4840_out0 || v$G$CD_1168_out0;
assign v$G8_11941_out0 = v$CINA_8786_out0 && v$P$AB_2180_out0;
assign v$G8_11948_out0 = v$CINA_8793_out0 && v$P$AB_2187_out0;
assign v$G8_11952_out0 = v$CINA_8797_out0 && v$P$AB_2191_out0;
assign v$G8_11955_out0 = v$CINA_8800_out0 && v$P$AB_2194_out0;
assign v$G8_11963_out0 = v$CINA_8808_out0 && v$P$AB_2202_out0;
assign v$G8_12064_out0 = v$CINA_8909_out0 && v$P$AB_2303_out0;
assign v$G8_12071_out0 = v$CINA_8916_out0 && v$P$AB_2310_out0;
assign v$G8_12075_out0 = v$CINA_8920_out0 && v$P$AB_2314_out0;
assign v$G8_12078_out0 = v$CINA_8923_out0 && v$P$AB_2317_out0;
assign v$G8_12086_out0 = v$CINA_8931_out0 && v$P$AB_2325_out0;
assign v$C9_12716_out0 = v$C9_6216_out0;
assign v$C9_12719_out0 = v$C9_6219_out0;
assign {v$A15_13797_out1,v$A15_13797_out0 } = v$A18_18300_out0 + v$B18_11368_out0 + v$C17_2716_out0;
assign {v$A15_13800_out1,v$A15_13800_out0 } = v$A18_18303_out0 + v$B18_11371_out0 + v$C17_2719_out0;
assign {v$A16A_15158_out1,v$A16A_15158_out0 } = v$A10_1703_out0 + v$B10_10297_out0 + v$C9_6216_out0;
assign {v$A16A_15161_out1,v$A16A_15161_out0 } = v$A10_1706_out0 + v$B10_10300_out0 + v$C9_6219_out0;
assign v$SEL1_15992_out0 = v$IN_4040_out0[7:0];
assign v$SEL1_16002_out0 = v$IN_4043_out0[7:0];
assign v$SEL1_16023_out0 = v$IN_4049_out0[7:0];
assign v$SEL1_16033_out0 = v$IN_4052_out0[7:0];
assign v$C23_16758_out0 = v$C23_5056_out0;
assign v$C23_16761_out0 = v$C23_5059_out0;
assign {v$A20_16992_out1,v$A20_16992_out0 } = v$A14_738_out0 + v$B14_4158_out0 + v$C13_12346_out0;
assign {v$A20_16995_out1,v$A20_16995_out0 } = v$A14_741_out0 + v$B14_4161_out0 + v$C13_12349_out0;
assign v$C13_19197_out0 = v$C13_12346_out0;
assign v$C13_19200_out0 = v$C13_12349_out0;
assign v$ENDq_1609_out0 = v$A12A_4613_out1;
assign v$ENDq_1612_out0 = v$A12A_4616_out1;
assign v$_4424_out0 = { v$C2_122_out0,v$SEL1_15992_out0 };
assign v$_4434_out0 = { v$C2_132_out0,v$SEL1_16002_out0 };
assign v$_4455_out0 = { v$C2_153_out0,v$SEL1_16023_out0 };
assign v$_4465_out0 = { v$C2_163_out0,v$SEL1_16033_out0 };
assign v$_6173_out0 = { v$A17A_2682_out0,v$A18_10458_out0 };
assign v$_6176_out0 = { v$A17A_2685_out0,v$A18_10461_out0 };
assign v$CARRY_6582_out0 = v$C23_16758_out0;
assign v$CARRY_6585_out0 = v$C23_16761_out0;
assign v$ENDr_7842_out0 = v$A20_16992_out1;
assign v$ENDr_7845_out0 = v$A20_16995_out1;
assign v$_7874_out0 = { v$C8_19107_out0,v$C9_12716_out0 };
assign v$_7877_out0 = { v$C8_19110_out0,v$C9_12719_out0 };
assign v$ENDi_9030_out0 = v$A15_13797_out1;
assign v$ENDi_9033_out0 = v$A15_13800_out1;
assign v$_9325_out0 = { v$SEL1_9064_out0,v$C1_6260_out0 };
assign v$_9335_out0 = { v$SEL1_9074_out0,v$C1_6270_out0 };
assign v$_9356_out0 = { v$SEL1_9095_out0,v$C1_6291_out0 };
assign v$_9366_out0 = { v$SEL1_9105_out0,v$C1_6301_out0 };
assign v$END0_9721_out0 = v$A16A_15158_out1;
assign v$END0_9724_out0 = v$A16A_15161_out1;
assign v$G7_10033_out0 = v$G8_11941_out0 && v$P$CD_10922_out0;
assign v$G7_10040_out0 = v$G8_11948_out0 && v$P$CD_10929_out0;
assign v$G7_10044_out0 = v$G8_11952_out0 && v$P$CD_10933_out0;
assign v$G7_10047_out0 = v$G8_11955_out0 && v$P$CD_10936_out0;
assign v$G7_10055_out0 = v$G8_11963_out0 && v$P$CD_10944_out0;
assign v$G7_10156_out0 = v$G8_12064_out0 && v$P$CD_11045_out0;
assign v$G7_10163_out0 = v$G8_12071_out0 && v$P$CD_11052_out0;
assign v$G7_10167_out0 = v$G8_12075_out0 && v$P$CD_11056_out0;
assign v$G7_10170_out0 = v$G8_12078_out0 && v$P$CD_11059_out0;
assign v$G7_10178_out0 = v$G8_12086_out0 && v$P$CD_11067_out0;
assign v$_10689_out0 = { v$C12_9767_out0,v$C13_19197_out0 };
assign v$_10692_out0 = { v$C12_9770_out0,v$C13_19200_out0 };
assign v$ENDt_10711_out0 = v$A13_7554_out1;
assign v$ENDt_10714_out0 = v$A13_7557_out1;
assign v$_11463_out0 = { v$A16A_15158_out0,v$A12A_4613_out0 };
assign v$_11466_out0 = { v$A16A_15161_out0,v$A12A_4616_out0 };
assign v$_15446_out0 = { v$C10_2103_out0,v$C11_9887_out0 };
assign v$_15449_out0 = { v$C10_2106_out0,v$C11_9890_out0 };
assign v$G$AD_17693_out0 = v$G4_11619_out0;
assign v$G$AD_17712_out0 = v$G4_11638_out0;
assign v$G$AD_17816_out0 = v$G4_11742_out0;
assign v$G$AD_17835_out0 = v$G4_11761_out0;
assign v$_18098_out0 = { v$A20_16992_out0,v$A13_7554_out0 };
assign v$_18101_out0 = { v$A20_16995_out0,v$A13_7557_out0 };
assign v$ENDe_18504_out0 = v$A18_10458_out1;
assign v$ENDe_18507_out0 = v$A18_10461_out1;
assign v$G6_468_out0 = v$G4_11626_out0 || v$G7_10033_out0;
assign v$G6_475_out0 = v$G4_11633_out0 || v$G7_10040_out0;
assign v$G6_479_out0 = v$G4_11637_out0 || v$G7_10044_out0;
assign v$G6_482_out0 = v$G4_11640_out0 || v$G7_10047_out0;
assign v$G6_490_out0 = v$G4_11648_out0 || v$G7_10055_out0;
assign v$G6_591_out0 = v$G4_11749_out0 || v$G7_10156_out0;
assign v$G6_598_out0 = v$G4_11756_out0 || v$G7_10163_out0;
assign v$G6_602_out0 = v$G4_11760_out0 || v$G7_10167_out0;
assign v$G6_605_out0 = v$G4_11763_out0 || v$G7_10170_out0;
assign v$G6_613_out0 = v$G4_11771_out0 || v$G7_10178_out0;
assign v$_1713_out0 = { v$_15630_out0,v$_11463_out0 };
assign v$_1716_out0 = { v$_15633_out0,v$_11466_out0 };
assign v$MUX1_2561_out0 = v$LEFT$SHIT_3273_out0 ? v$_4424_out0 : v$_9325_out0;
assign v$MUX1_2571_out0 = v$LEFT$SHIT_3283_out0 ? v$_4434_out0 : v$_9335_out0;
assign v$MUX1_2592_out0 = v$LEFT$SHIT_3304_out0 ? v$_4455_out0 : v$_9356_out0;
assign v$MUX1_2602_out0 = v$LEFT$SHIT_3314_out0 ? v$_4465_out0 : v$_9366_out0;
assign v$TWOS$COMPLEMENT$ADDER$COUT_3639_out0 = v$CARRY_6582_out0;
assign v$TWOS$COMPLEMENT$ADDER$COUT_3640_out0 = v$CARRY_6585_out0;
assign v$END50_7729_out0 = v$G$AD_17693_out0;
assign v$END50_7732_out0 = v$G$AD_17816_out0;
assign v$END48_10827_out0 = v$G$AD_17712_out0;
assign v$END48_10830_out0 = v$G$AD_17835_out0;
assign v$_14896_out0 = { v$_6173_out0,v$_18098_out0 };
assign v$_14899_out0 = { v$_6176_out0,v$_18101_out0 };
assign v$_18907_out0 = { v$_7874_out0,v$_15446_out0 };
assign v$_18910_out0 = { v$_7877_out0,v$_15449_out0 };
assign v$_1319_out0 = { v$_1713_out0,v$_14896_out0 };
assign v$_1322_out0 = { v$_1716_out0,v$_14899_out0 };
assign v$COUTD_6946_out0 = v$G6_468_out0;
assign v$COUTD_6953_out0 = v$G6_475_out0;
assign v$COUTD_6957_out0 = v$G6_479_out0;
assign v$COUTD_6960_out0 = v$G6_482_out0;
assign v$COUTD_6968_out0 = v$G6_490_out0;
assign v$COUTD_7069_out0 = v$G6_591_out0;
assign v$COUTD_7076_out0 = v$G6_598_out0;
assign v$COUTD_7080_out0 = v$G6_602_out0;
assign v$COUTD_7083_out0 = v$G6_605_out0;
assign v$COUTD_7091_out0 = v$G6_613_out0;
assign v$MUX2_19188_out0 = v$EN_5430_out0 ? v$MUX1_2561_out0 : v$IN_4040_out0;
assign v$MUX2_19190_out0 = v$EN_5432_out0 ? v$MUX1_2571_out0 : v$IN_4043_out0;
assign v$MUX2_19194_out0 = v$EN_5436_out0 ? v$MUX1_2592_out0 : v$IN_4049_out0;
assign v$MUX2_19196_out0 = v$EN_5438_out0 ? v$MUX1_2602_out0 : v$IN_4052_out0;
assign v$C16_1423_out0 = v$COUTD_6960_out0;
assign v$C16_1426_out0 = v$COUTD_7083_out0;
assign v$C15_8447_out0 = v$COUTD_6957_out0;
assign v$C15_8450_out0 = v$COUTD_7080_out0;
assign v$C19_8467_out0 = v$COUTD_6968_out0;
assign v$C19_8470_out0 = v$COUTD_7091_out0;
assign v$CINA_8779_out0 = v$COUTD_6953_out0;
assign v$CINA_8798_out0 = v$COUTD_6953_out0;
assign v$CINA_8902_out0 = v$COUTD_7076_out0;
assign v$CINA_8921_out0 = v$COUTD_7076_out0;
assign v$OUT_15533_out0 = v$MUX2_19188_out0;
assign v$OUT_15543_out0 = v$MUX2_19190_out0;
assign v$OUT_15564_out0 = v$MUX2_19194_out0;
assign v$OUT_15574_out0 = v$MUX2_19196_out0;
assign v$C20_16079_out0 = v$COUTD_6953_out0;
assign v$C20_16082_out0 = v$COUTD_7076_out0;
assign v$C18_16902_out0 = v$COUTD_6946_out0;
assign v$C18_16905_out0 = v$COUTD_7069_out0;
assign v$_18834_out0 = { v$_18358_out0,v$_1319_out0 };
assign v$_18837_out0 = { v$_18361_out0,v$_1322_out0 };
assign v$OUT_5128_out0 = v$OUT_15533_out0;
assign v$OUT_5129_out0 = v$OUT_15543_out0;
assign v$OUT_5130_out0 = v$OUT_15564_out0;
assign v$OUT_5131_out0 = v$OUT_15574_out0;
assign v$G8_11934_out0 = v$CINA_8779_out0 && v$P$AB_2173_out0;
assign v$G8_11953_out0 = v$CINA_8798_out0 && v$P$AB_2192_out0;
assign v$G8_12057_out0 = v$CINA_8902_out0 && v$P$AB_2296_out0;
assign v$G8_12076_out0 = v$CINA_8921_out0 && v$P$AB_2315_out0;
assign v$C15_13707_out0 = v$C15_8447_out0;
assign v$C15_13710_out0 = v$C15_8450_out0;
assign v$C19_14421_out0 = v$C19_8467_out0;
assign v$C19_14424_out0 = v$C19_8470_out0;
assign v$C20_15592_out0 = v$C20_16079_out0;
assign v$C20_15595_out0 = v$C20_16082_out0;
assign v$C16_15768_out0 = v$C16_1423_out0;
assign v$C16_15771_out0 = v$C16_1426_out0;
assign {v$A14_15941_out1,v$A14_15941_out0 } = v$A16_14191_out0 + v$B16_17034_out0 + v$C15_8447_out0;
assign {v$A14_15944_out1,v$A14_15944_out0 } = v$A16_14194_out0 + v$B16_17037_out0 + v$C15_8450_out0;
assign {v$A19_16511_out1,v$A19_16511_out0 } = v$A19_1363_out0 + v$B19_17410_out0 + v$C18_16902_out0;
assign {v$A19_16514_out1,v$A19_16514_out0 } = v$A19_1366_out0 + v$B19_17413_out0 + v$C18_16905_out0;
assign {v$A24_17569_out1,v$A24_17569_out0 } = v$A21_2792_out0 + v$B21_18689_out0 + v$C20_16079_out0;
assign {v$A24_17572_out1,v$A24_17572_out0 } = v$A21_2795_out0 + v$B21_18692_out0 + v$C20_16082_out0;
assign {v$A22_18127_out1,v$A22_18127_out0 } = v$A20_4603_out0 + v$B20_4112_out0 + v$C19_8467_out0;
assign {v$A22_18130_out1,v$A22_18130_out0 } = v$A20_4606_out0 + v$B20_4115_out0 + v$C19_8470_out0;
assign {v$A11_18484_out1,v$A11_18484_out0 } = v$A17_17342_out0 + v$B17_16125_out0 + v$C16_1423_out0;
assign {v$A11_18487_out1,v$A11_18487_out0 } = v$A17_17345_out0 + v$B17_16128_out0 + v$C16_1426_out0;
assign v$C18_18609_out0 = v$C18_16902_out0;
assign v$C18_18612_out0 = v$C18_16905_out0;
assign v$_1347_out0 = { v$A15_13797_out0,v$A19_16511_out0 };
assign v$_1350_out0 = { v$A15_13800_out0,v$A19_16514_out0 };
assign v$_1954_out0 = { v$A22_18127_out0,v$A24_17569_out0 };
assign v$_1957_out0 = { v$A22_18130_out0,v$A24_17572_out0 };
assign v$_3064_out0 = { v$C14_340_out0,v$C15_13707_out0 };
assign v$_3067_out0 = { v$C14_343_out0,v$C15_13710_out0 };
assign v$ENDp_3409_out0 = v$A22_18127_out1;
assign v$ENDp_3412_out0 = v$A22_18130_out1;
assign v$ENDy_4271_out0 = v$A14_15941_out1;
assign v$ENDy_4274_out0 = v$A14_15944_out1;
assign v$SEL1_6308_out0 = v$OUT_5129_out0[22:0];
assign v$SEL1_6309_out0 = v$OUT_5131_out0[22:0];
assign v$ENDu_7313_out0 = v$A11_18484_out1;
assign v$ENDu_7316_out0 = v$A11_18487_out1;
assign v$_8193_out0 = { v$C16_15768_out0,v$C17_6342_out0 };
assign v$_8196_out0 = { v$C16_15771_out0,v$C17_6345_out0 };
assign v$SEL2_8412_out0 = v$OUT_5128_out0[22:13];
assign v$SEL2_8413_out0 = v$OUT_5130_out0[22:13];
assign v$_8641_out0 = { v$C18_18609_out0,v$C19_14421_out0 };
assign v$_8644_out0 = { v$C18_18612_out0,v$C19_14424_out0 };
assign v$G7_10026_out0 = v$G8_11934_out0 && v$P$CD_10915_out0;
assign v$G7_10045_out0 = v$G8_11953_out0 && v$P$CD_10934_out0;
assign v$G7_10149_out0 = v$G8_12057_out0 && v$P$CD_11038_out0;
assign v$G7_10168_out0 = v$G8_12076_out0 && v$P$CD_11057_out0;
assign v$_13877_out0 = { v$A14_15941_out0,v$A11_18484_out0 };
assign v$_13880_out0 = { v$A14_15944_out0,v$A11_18487_out0 };
assign v$ENDa_17183_out0 = v$A24_17569_out1;
assign v$ENDa_17186_out0 = v$A24_17572_out1;
assign v$ENDo_19304_out0 = v$A19_16511_out1;
assign v$ENDo_19307_out0 = v$A19_16514_out1;
assign v$G6_461_out0 = v$G4_11619_out0 || v$G7_10026_out0;
assign v$G6_480_out0 = v$G4_11638_out0 || v$G7_10045_out0;
assign v$G6_584_out0 = v$G4_11742_out0 || v$G7_10149_out0;
assign v$G6_603_out0 = v$G4_11761_out0 || v$G7_10168_out0;
assign v$_1395_out0 = { v$_10689_out0,v$_3064_out0 };
assign v$_1398_out0 = { v$_10692_out0,v$_3067_out0 };
assign v$_10811_out0 = { v$_8193_out0,v$_8641_out0 };
assign v$_10814_out0 = { v$_8196_out0,v$_8644_out0 };
assign v$_16450_out0 = { v$SEL2_8412_out0,v$A2_10470_out0 };
assign v$_16451_out0 = { v$SEL1_6308_out0,v$A2_10471_out0 };
assign v$_16452_out0 = { v$SEL2_8413_out0,v$A2_10472_out0 };
assign v$_16453_out0 = { v$SEL1_6309_out0,v$A2_10473_out0 };
assign v$_16866_out0 = { v$_13877_out0,v$_1347_out0 };
assign v$_16869_out0 = { v$_13880_out0,v$_1350_out0 };
assign v$COUTD_6939_out0 = v$G6_461_out0;
assign v$COUTD_6958_out0 = v$G6_480_out0;
assign v$COUTD_7062_out0 = v$G6_584_out0;
assign v$COUTD_7081_out0 = v$G6_603_out0;
assign v$MUX2_14208_out0 = v$Z_16411_out0 ? v$C4_8566_out0 : v$_16450_out0;
assign v$MUX2_14209_out0 = v$Z_16412_out0 ? v$C4_8567_out0 : v$_16451_out0;
assign v$MUX2_14210_out0 = v$Z_16413_out0 ? v$C4_8568_out0 : v$_16452_out0;
assign v$MUX2_14211_out0 = v$Z_16414_out0 ? v$C4_8569_out0 : v$_16453_out0;
assign v$_17995_out0 = { v$_18907_out0,v$_1395_out0 };
assign v$_17998_out0 = { v$_18910_out0,v$_1398_out0 };
assign v$_5082_out0 = { v$_8112_out0,v$_17995_out0 };
assign v$_5085_out0 = { v$_8115_out0,v$_17998_out0 };
assign v$C21_11258_out0 = v$COUTD_6958_out0;
assign v$C21_11261_out0 = v$COUTD_7081_out0;
assign v$C22_11488_out0 = v$COUTD_6939_out0;
assign v$C22_11491_out0 = v$COUTD_7062_out0;
assign v$_19023_out0 = { v$MUX2_14208_out0,v$SIGN_1529_out0 };
assign v$_19024_out0 = { v$MUX2_14209_out0,v$SIGN_1530_out0 };
assign v$_19025_out0 = { v$MUX2_14210_out0,v$SIGN_1531_out0 };
assign v$_19026_out0 = { v$MUX2_14211_out0,v$SIGN_1532_out0 };
assign v$C21_6608_out0 = v$C21_11258_out0;
assign v$C21_6611_out0 = v$C21_11261_out0;
assign v$C22_8714_out0 = v$C22_11488_out0;
assign v$C22_8717_out0 = v$C22_11491_out0;
assign {v$A23_9924_out1,v$A23_9924_out0 } = v$A23_5281_out0 + v$B23_1441_out0 + v$C22_11488_out0;
assign {v$A23_9927_out1,v$A23_9927_out0 } = v$A23_5284_out0 + v$B23_1444_out0 + v$C22_11491_out0;
assign v$OUT_13072_out0 = v$_19023_out0;
assign v$OUT_13073_out0 = v$_19024_out0;
assign v$OUT_13074_out0 = v$_19025_out0;
assign v$OUT_13075_out0 = v$_19026_out0;
assign {v$A21_19179_out1,v$A21_19179_out0 } = v$A22_4590_out0 + v$B22_11300_out0 + v$C21_11258_out0;
assign {v$A21_19182_out1,v$A21_19182_out0 } = v$A22_4593_out0 + v$B22_11303_out0 + v$C21_11261_out0;
assign v$_710_out0 = { v$C20_15592_out0,v$C21_6608_out0 };
assign v$_713_out0 = { v$C20_15595_out0,v$C21_6611_out0 };
assign v$_1733_out0 = { v$A21_19179_out0,v$A23_9924_out0 };
assign v$_1736_out0 = { v$A21_19182_out0,v$A23_9927_out0 };
assign v$ENDs_3435_out0 = v$A21_19179_out1;
assign v$ENDs_3438_out0 = v$A21_19182_out1;
assign v$MUX11_9016_out0 = v$G5_6460_out0 ? v$C9_19371_out0 : v$OUT_13072_out0;
assign v$MUX11_9017_out0 = v$G5_6461_out0 ? v$C9_19372_out0 : v$OUT_13074_out0;
assign v$MUX3_9291_out0 = v$G3_16620_out0 ? v$C1_15809_out0 : v$OUT_13073_out0;
assign v$MUX3_9292_out0 = v$G3_16621_out0 ? v$C1_15810_out0 : v$OUT_13075_out0;
assign v$ENDd_11330_out0 = v$A23_9924_out1;
assign v$ENDd_11333_out0 = v$A23_9927_out1;
assign v$_16303_out0 = { v$C22_8714_out0,v$C23_16758_out0 };
assign v$_16306_out0 = { v$C22_8717_out0,v$C23_16761_out0 };
assign v$SINGLE$PRECISION_8227_out0 = v$MUX3_9291_out0;
assign v$SINGLE$PRECISION_8228_out0 = v$MUX3_9292_out0;
assign v$_9865_out0 = { v$_1954_out0,v$_1733_out0 };
assign v$_9868_out0 = { v$_1957_out0,v$_1736_out0 };
assign v$_14314_out0 = { v$_710_out0,v$_16303_out0 };
assign v$_14317_out0 = { v$_713_out0,v$_16306_out0 };
assign v$_17630_out0 = { v$C10_6624_out0,v$MUX11_9016_out0 };
assign v$_17631_out0 = { v$C10_6625_out0,v$MUX11_9017_out0 };
assign v$_4248_out0 = { v$_10811_out0,v$_14314_out0 };
assign v$_4251_out0 = { v$_10814_out0,v$_14317_out0 };
assign v$_6893_out0 = { v$_16866_out0,v$_9865_out0 };
assign v$_6896_out0 = { v$_16869_out0,v$_9868_out0 };
assign v$HALF$PRECISION_10767_out0 = v$_17630_out0;
assign v$HALF$PRECISION_10768_out0 = v$_17631_out0;
assign v$_3939_out0 = { v$_5082_out0,v$_4248_out0 };
assign v$_3942_out0 = { v$_5085_out0,v$_4251_out0 };
assign v$_10327_out0 = { v$_18834_out0,v$_6893_out0 };
assign v$_10330_out0 = { v$_18837_out0,v$_6896_out0 };
assign v$MUX12_17418_out0 = v$IS$32$BITS_3203_out0 ? v$SINGLE$PRECISION_8227_out0 : v$HALF$PRECISION_10767_out0;
assign v$MUX12_17419_out0 = v$IS$32$BITS_3204_out0 ? v$SINGLE$PRECISION_8228_out0 : v$HALF$PRECISION_10768_out0;
assign v$OUT_3588_out0 = v$MUX12_17418_out0;
assign v$OUT_3589_out0 = v$MUX12_17419_out0;
assign v$SUM_9731_out0 = v$_10327_out0;
assign v$SUM_9734_out0 = v$_10330_out0;
assign v$SUM1_13397_out0 = v$_3939_out0;
assign v$SUM1_13400_out0 = v$_3942_out0;
assign v$END_2032_out0 = v$SUM1_13397_out0;
assign v$END_2033_out0 = v$SUM1_13400_out0;
assign v$MUX5_6486_out0 = v$IS$A$LARGER_10896_out0 ? v$SUM_2068_out0 : v$SUM_9731_out0;
assign v$MUX5_6487_out0 = v$IS$A$LARGER_10897_out0 ? v$SUM_2069_out0 : v$SUM_9734_out0;
assign v$LZD$INPUT_9184_out0 = v$MUX5_6486_out0;
assign v$LZD$INPUT_9185_out0 = v$MUX5_6487_out0;
assign v$IN_13745_out0 = v$LZD$INPUT_9184_out0;
assign v$IN_13749_out0 = v$LZD$INPUT_9185_out0;
assign v$IN_18605_out0 = v$LZD$INPUT_9184_out0;
assign v$IN_18606_out0 = v$LZD$INPUT_9185_out0;
assign v$SEL1_368_out0 = v$IN_18605_out0[23:16];
assign v$SEL1_369_out0 = v$IN_18606_out0[23:16];
assign v$IN_5377_out0 = v$IN_13745_out0;
assign v$IN_5408_out0 = v$IN_13749_out0;
assign v$SEL2_18013_out0 = v$IN_18605_out0[15:8];
assign v$SEL2_18014_out0 = v$IN_18606_out0[15:8];
assign v$SEL1_18066_out0 = v$IN_18605_out0[7:0];
assign v$SEL1_18067_out0 = v$IN_18606_out0[7:0];
assign v$IN_4038_out0 = v$IN_5377_out0;
assign v$IN_4047_out0 = v$IN_5408_out0;
assign v$IN_15465_out0 = v$SEL1_368_out0;
assign v$IN_15466_out0 = v$SEL2_18013_out0;
assign v$IN_15467_out0 = v$SEL1_18066_out0;
assign v$IN_15470_out0 = v$SEL1_369_out0;
assign v$IN_15471_out0 = v$SEL2_18014_out0;
assign v$IN_15472_out0 = v$SEL1_18067_out0;
assign v$SEL2_3235_out0 = v$IN_15465_out0[7:4];
assign v$SEL2_3236_out0 = v$IN_15466_out0[7:4];
assign v$SEL2_3237_out0 = v$IN_15467_out0[7:4];
assign v$SEL2_3240_out0 = v$IN_15470_out0[7:4];
assign v$SEL2_3241_out0 = v$IN_15471_out0[7:4];
assign v$SEL2_3242_out0 = v$IN_15472_out0[7:4];
assign v$SEL1_9058_out0 = v$IN_4038_out0[23:1];
assign v$SEL1_9089_out0 = v$IN_4047_out0[23:1];
assign v$SEL1_15986_out0 = v$IN_4038_out0[22:0];
assign v$SEL1_16017_out0 = v$IN_4047_out0[22:0];
assign v$SEL1_17079_out0 = v$IN_15465_out0[3:0];
assign v$SEL1_17080_out0 = v$IN_15466_out0[3:0];
assign v$SEL1_17081_out0 = v$IN_15467_out0[3:0];
assign v$SEL1_17084_out0 = v$IN_15470_out0[3:0];
assign v$SEL1_17085_out0 = v$IN_15471_out0[3:0];
assign v$SEL1_17086_out0 = v$IN_15472_out0[3:0];
assign v$_4418_out0 = { v$C2_116_out0,v$SEL1_15986_out0 };
assign v$_4449_out0 = { v$C2_147_out0,v$SEL1_16017_out0 };
assign v$_9319_out0 = { v$SEL1_9058_out0,v$C1_6254_out0 };
assign v$_9350_out0 = { v$SEL1_9089_out0,v$C1_6285_out0 };
assign v$IN_15677_out0 = v$SEL1_17079_out0;
assign v$IN_15678_out0 = v$SEL2_3235_out0;
assign v$IN_15679_out0 = v$SEL1_17080_out0;
assign v$IN_15680_out0 = v$SEL2_3236_out0;
assign v$IN_15681_out0 = v$SEL1_17081_out0;
assign v$IN_15682_out0 = v$SEL2_3237_out0;
assign v$IN_15695_out0 = v$SEL1_17084_out0;
assign v$IN_15696_out0 = v$SEL2_3240_out0;
assign v$IN_15697_out0 = v$SEL1_17085_out0;
assign v$IN_15698_out0 = v$SEL2_3241_out0;
assign v$IN_15699_out0 = v$SEL1_17086_out0;
assign v$IN_15700_out0 = v$SEL2_3242_out0;
assign v$SEL3_2499_out0 = v$IN_15677_out0[2:2];
assign v$SEL3_2500_out0 = v$IN_15678_out0[2:2];
assign v$SEL3_2501_out0 = v$IN_15679_out0[2:2];
assign v$SEL3_2502_out0 = v$IN_15680_out0[2:2];
assign v$SEL3_2503_out0 = v$IN_15681_out0[2:2];
assign v$SEL3_2504_out0 = v$IN_15682_out0[2:2];
assign v$SEL3_2517_out0 = v$IN_15695_out0[2:2];
assign v$SEL3_2518_out0 = v$IN_15696_out0[2:2];
assign v$SEL3_2519_out0 = v$IN_15697_out0[2:2];
assign v$SEL3_2520_out0 = v$IN_15698_out0[2:2];
assign v$SEL3_2521_out0 = v$IN_15699_out0[2:2];
assign v$SEL3_2522_out0 = v$IN_15700_out0[2:2];
assign v$MUX1_2555_out0 = v$LEFT$SHIT_3267_out0 ? v$_4418_out0 : v$_9319_out0;
assign v$MUX1_2586_out0 = v$LEFT$SHIT_3298_out0 ? v$_4449_out0 : v$_9350_out0;
assign v$SEL4_6356_out0 = v$IN_15677_out0[3:3];
assign v$SEL4_6357_out0 = v$IN_15678_out0[3:3];
assign v$SEL4_6358_out0 = v$IN_15679_out0[3:3];
assign v$SEL4_6359_out0 = v$IN_15680_out0[3:3];
assign v$SEL4_6360_out0 = v$IN_15681_out0[3:3];
assign v$SEL4_6361_out0 = v$IN_15682_out0[3:3];
assign v$SEL4_6374_out0 = v$IN_15695_out0[3:3];
assign v$SEL4_6375_out0 = v$IN_15696_out0[3:3];
assign v$SEL4_6376_out0 = v$IN_15697_out0[3:3];
assign v$SEL4_6377_out0 = v$IN_15698_out0[3:3];
assign v$SEL4_6378_out0 = v$IN_15699_out0[3:3];
assign v$SEL4_6379_out0 = v$IN_15700_out0[3:3];
assign v$SEL2_7999_out0 = v$IN_15677_out0[1:1];
assign v$SEL2_8000_out0 = v$IN_15678_out0[1:1];
assign v$SEL2_8001_out0 = v$IN_15679_out0[1:1];
assign v$SEL2_8002_out0 = v$IN_15680_out0[1:1];
assign v$SEL2_8003_out0 = v$IN_15681_out0[1:1];
assign v$SEL2_8004_out0 = v$IN_15682_out0[1:1];
assign v$SEL2_8017_out0 = v$IN_15695_out0[1:1];
assign v$SEL2_8018_out0 = v$IN_15696_out0[1:1];
assign v$SEL2_8019_out0 = v$IN_15697_out0[1:1];
assign v$SEL2_8020_out0 = v$IN_15698_out0[1:1];
assign v$SEL2_8021_out0 = v$IN_15699_out0[1:1];
assign v$SEL2_8022_out0 = v$IN_15700_out0[1:1];
assign v$SEL1_14044_out0 = v$IN_15677_out0[0:0];
assign v$SEL1_14045_out0 = v$IN_15678_out0[0:0];
assign v$SEL1_14046_out0 = v$IN_15679_out0[0:0];
assign v$SEL1_14047_out0 = v$IN_15680_out0[0:0];
assign v$SEL1_14048_out0 = v$IN_15681_out0[0:0];
assign v$SEL1_14049_out0 = v$IN_15682_out0[0:0];
assign v$SEL1_14062_out0 = v$IN_15695_out0[0:0];
assign v$SEL1_14063_out0 = v$IN_15696_out0[0:0];
assign v$SEL1_14064_out0 = v$IN_15697_out0[0:0];
assign v$SEL1_14065_out0 = v$IN_15698_out0[0:0];
assign v$SEL1_14066_out0 = v$IN_15699_out0[0:0];
assign v$SEL1_14067_out0 = v$IN_15700_out0[0:0];
assign v$G10_1543_out0 = !(v$SEL1_14044_out0 || v$SEL2_7999_out0);
assign v$G10_1544_out0 = !(v$SEL1_14045_out0 || v$SEL2_8000_out0);
assign v$G10_1545_out0 = !(v$SEL1_14046_out0 || v$SEL2_8001_out0);
assign v$G10_1546_out0 = !(v$SEL1_14047_out0 || v$SEL2_8002_out0);
assign v$G10_1547_out0 = !(v$SEL1_14048_out0 || v$SEL2_8003_out0);
assign v$G10_1548_out0 = !(v$SEL1_14049_out0 || v$SEL2_8004_out0);
assign v$G10_1561_out0 = !(v$SEL1_14062_out0 || v$SEL2_8017_out0);
assign v$G10_1562_out0 = !(v$SEL1_14063_out0 || v$SEL2_8018_out0);
assign v$G10_1563_out0 = !(v$SEL1_14064_out0 || v$SEL2_8019_out0);
assign v$G10_1564_out0 = !(v$SEL1_14065_out0 || v$SEL2_8020_out0);
assign v$G10_1565_out0 = !(v$SEL1_14066_out0 || v$SEL2_8021_out0);
assign v$G10_1566_out0 = !(v$SEL1_14067_out0 || v$SEL2_8022_out0);
assign v$G6_3756_out0 = ! v$SEL2_7999_out0;
assign v$G6_3757_out0 = ! v$SEL2_8000_out0;
assign v$G6_3758_out0 = ! v$SEL2_8001_out0;
assign v$G6_3759_out0 = ! v$SEL2_8002_out0;
assign v$G6_3760_out0 = ! v$SEL2_8003_out0;
assign v$G6_3761_out0 = ! v$SEL2_8004_out0;
assign v$G6_3774_out0 = ! v$SEL2_8017_out0;
assign v$G6_3775_out0 = ! v$SEL2_8018_out0;
assign v$G6_3776_out0 = ! v$SEL2_8019_out0;
assign v$G6_3777_out0 = ! v$SEL2_8020_out0;
assign v$G6_3778_out0 = ! v$SEL2_8021_out0;
assign v$G6_3779_out0 = ! v$SEL2_8022_out0;
assign v$G5_6119_out0 = ! v$SEL4_6356_out0;
assign v$G5_6120_out0 = ! v$SEL4_6357_out0;
assign v$G5_6121_out0 = ! v$SEL4_6358_out0;
assign v$G5_6122_out0 = ! v$SEL4_6359_out0;
assign v$G5_6123_out0 = ! v$SEL4_6360_out0;
assign v$G5_6124_out0 = ! v$SEL4_6361_out0;
assign v$G5_6137_out0 = ! v$SEL4_6374_out0;
assign v$G5_6138_out0 = ! v$SEL4_6375_out0;
assign v$G5_6139_out0 = ! v$SEL4_6376_out0;
assign v$G5_6140_out0 = ! v$SEL4_6377_out0;
assign v$G5_6141_out0 = ! v$SEL4_6378_out0;
assign v$G5_6142_out0 = ! v$SEL4_6379_out0;
assign v$G11_9189_out0 = !(v$SEL3_2499_out0 || v$SEL4_6356_out0);
assign v$G11_9190_out0 = !(v$SEL3_2500_out0 || v$SEL4_6357_out0);
assign v$G11_9191_out0 = !(v$SEL3_2501_out0 || v$SEL4_6358_out0);
assign v$G11_9192_out0 = !(v$SEL3_2502_out0 || v$SEL4_6359_out0);
assign v$G11_9193_out0 = !(v$SEL3_2503_out0 || v$SEL4_6360_out0);
assign v$G11_9194_out0 = !(v$SEL3_2504_out0 || v$SEL4_6361_out0);
assign v$G11_9207_out0 = !(v$SEL3_2517_out0 || v$SEL4_6374_out0);
assign v$G11_9208_out0 = !(v$SEL3_2518_out0 || v$SEL4_6375_out0);
assign v$G11_9209_out0 = !(v$SEL3_2519_out0 || v$SEL4_6376_out0);
assign v$G11_9210_out0 = !(v$SEL3_2520_out0 || v$SEL4_6377_out0);
assign v$G11_9211_out0 = !(v$SEL3_2521_out0 || v$SEL4_6378_out0);
assign v$G11_9212_out0 = !(v$SEL3_2522_out0 || v$SEL4_6379_out0);
assign v$G8_12567_out0 = ! v$SEL3_2499_out0;
assign v$G8_12568_out0 = ! v$SEL3_2500_out0;
assign v$G8_12569_out0 = ! v$SEL3_2501_out0;
assign v$G8_12570_out0 = ! v$SEL3_2502_out0;
assign v$G8_12571_out0 = ! v$SEL3_2503_out0;
assign v$G8_12572_out0 = ! v$SEL3_2504_out0;
assign v$G8_12585_out0 = ! v$SEL3_2517_out0;
assign v$G8_12586_out0 = ! v$SEL3_2518_out0;
assign v$G8_12587_out0 = ! v$SEL3_2519_out0;
assign v$G8_12588_out0 = ! v$SEL3_2520_out0;
assign v$G8_12589_out0 = ! v$SEL3_2521_out0;
assign v$G8_12590_out0 = ! v$SEL3_2522_out0;
assign v$G3_13244_out0 = v$G10_1543_out0 && v$G11_9189_out0;
assign v$G3_13245_out0 = v$G10_1544_out0 && v$G11_9190_out0;
assign v$G3_13246_out0 = v$G10_1545_out0 && v$G11_9191_out0;
assign v$G3_13247_out0 = v$G10_1546_out0 && v$G11_9192_out0;
assign v$G3_13248_out0 = v$G10_1547_out0 && v$G11_9193_out0;
assign v$G3_13249_out0 = v$G10_1548_out0 && v$G11_9194_out0;
assign v$G3_13262_out0 = v$G10_1561_out0 && v$G11_9207_out0;
assign v$G3_13263_out0 = v$G10_1562_out0 && v$G11_9208_out0;
assign v$G3_13264_out0 = v$G10_1563_out0 && v$G11_9209_out0;
assign v$G3_13265_out0 = v$G10_1564_out0 && v$G11_9210_out0;
assign v$G3_13266_out0 = v$G10_1565_out0 && v$G11_9211_out0;
assign v$G3_13267_out0 = v$G10_1566_out0 && v$G11_9212_out0;
assign v$G9_18211_out0 = v$G8_12567_out0 && v$G5_6119_out0;
assign v$G9_18212_out0 = v$G8_12568_out0 && v$G5_6120_out0;
assign v$G9_18213_out0 = v$G8_12569_out0 && v$G5_6121_out0;
assign v$G9_18214_out0 = v$G8_12570_out0 && v$G5_6122_out0;
assign v$G9_18215_out0 = v$G8_12571_out0 && v$G5_6123_out0;
assign v$G9_18216_out0 = v$G8_12572_out0 && v$G5_6124_out0;
assign v$G9_18229_out0 = v$G8_12585_out0 && v$G5_6137_out0;
assign v$G9_18230_out0 = v$G8_12586_out0 && v$G5_6138_out0;
assign v$G9_18231_out0 = v$G8_12587_out0 && v$G5_6139_out0;
assign v$G9_18232_out0 = v$G8_12588_out0 && v$G5_6140_out0;
assign v$G9_18233_out0 = v$G8_12589_out0 && v$G5_6141_out0;
assign v$G9_18234_out0 = v$G8_12590_out0 && v$G5_6142_out0;
assign v$G7_18741_out0 = v$G6_3756_out0 || v$SEL3_2499_out0;
assign v$G7_18742_out0 = v$G6_3757_out0 || v$SEL3_2500_out0;
assign v$G7_18743_out0 = v$G6_3758_out0 || v$SEL3_2501_out0;
assign v$G7_18744_out0 = v$G6_3759_out0 || v$SEL3_2502_out0;
assign v$G7_18745_out0 = v$G6_3760_out0 || v$SEL3_2503_out0;
assign v$G7_18746_out0 = v$G6_3761_out0 || v$SEL3_2504_out0;
assign v$G7_18759_out0 = v$G6_3774_out0 || v$SEL3_2517_out0;
assign v$G7_18760_out0 = v$G6_3775_out0 || v$SEL3_2518_out0;
assign v$G7_18761_out0 = v$G6_3776_out0 || v$SEL3_2519_out0;
assign v$G7_18762_out0 = v$G6_3777_out0 || v$SEL3_2520_out0;
assign v$G7_18763_out0 = v$G6_3778_out0 || v$SEL3_2521_out0;
assign v$G7_18764_out0 = v$G6_3779_out0 || v$SEL3_2522_out0;
assign v$Z_13147_out0 = v$G3_13244_out0;
assign v$Z_13148_out0 = v$G3_13245_out0;
assign v$Z_13149_out0 = v$G3_13246_out0;
assign v$Z_13150_out0 = v$G3_13247_out0;
assign v$Z_13151_out0 = v$G3_13248_out0;
assign v$Z_13152_out0 = v$G3_13249_out0;
assign v$Z_13165_out0 = v$G3_13262_out0;
assign v$Z_13166_out0 = v$G3_13263_out0;
assign v$Z_13167_out0 = v$G3_13264_out0;
assign v$Z_13168_out0 = v$G3_13265_out0;
assign v$Z_13169_out0 = v$G3_13266_out0;
assign v$Z_13170_out0 = v$G3_13267_out0;
assign v$G4_18158_out0 = v$G7_18741_out0 && v$G5_6119_out0;
assign v$G4_18159_out0 = v$G7_18742_out0 && v$G5_6120_out0;
assign v$G4_18160_out0 = v$G7_18743_out0 && v$G5_6121_out0;
assign v$G4_18161_out0 = v$G7_18744_out0 && v$G5_6122_out0;
assign v$G4_18162_out0 = v$G7_18745_out0 && v$G5_6123_out0;
assign v$G4_18163_out0 = v$G7_18746_out0 && v$G5_6124_out0;
assign v$G4_18176_out0 = v$G7_18759_out0 && v$G5_6137_out0;
assign v$G4_18177_out0 = v$G7_18760_out0 && v$G5_6138_out0;
assign v$G4_18178_out0 = v$G7_18761_out0 && v$G5_6139_out0;
assign v$G4_18179_out0 = v$G7_18762_out0 && v$G5_6140_out0;
assign v$G4_18180_out0 = v$G7_18763_out0 && v$G5_6141_out0;
assign v$G4_18181_out0 = v$G7_18764_out0 && v$G5_6142_out0;
assign v$Z2_180_out0 = v$Z_13147_out0;
assign v$Z2_181_out0 = v$Z_13149_out0;
assign v$Z2_182_out0 = v$Z_13151_out0;
assign v$Z2_185_out0 = v$Z_13165_out0;
assign v$Z2_186_out0 = v$Z_13167_out0;
assign v$Z2_187_out0 = v$Z_13169_out0;
assign v$Z1_6049_out0 = v$Z_13148_out0;
assign v$Z1_6050_out0 = v$Z_13150_out0;
assign v$Z1_6051_out0 = v$Z_13152_out0;
assign v$Z1_6054_out0 = v$Z_13166_out0;
assign v$Z1_6055_out0 = v$Z_13168_out0;
assign v$Z1_6056_out0 = v$Z_13170_out0;
assign v$_6532_out0 = { v$G4_18158_out0,v$G9_18211_out0 };
assign v$_6533_out0 = { v$G4_18159_out0,v$G9_18212_out0 };
assign v$_6534_out0 = { v$G4_18160_out0,v$G9_18213_out0 };
assign v$_6535_out0 = { v$G4_18161_out0,v$G9_18214_out0 };
assign v$_6536_out0 = { v$G4_18162_out0,v$G9_18215_out0 };
assign v$_6537_out0 = { v$G4_18163_out0,v$G9_18216_out0 };
assign v$_6550_out0 = { v$G4_18176_out0,v$G9_18229_out0 };
assign v$_6551_out0 = { v$G4_18177_out0,v$G9_18230_out0 };
assign v$_6552_out0 = { v$G4_18178_out0,v$G9_18231_out0 };
assign v$_6553_out0 = { v$G4_18179_out0,v$G9_18232_out0 };
assign v$_6554_out0 = { v$G4_18180_out0,v$G9_18233_out0 };
assign v$_6555_out0 = { v$G4_18181_out0,v$G9_18234_out0 };
assign v$Y_6731_out0 = v$_6532_out0;
assign v$Y_6732_out0 = v$_6533_out0;
assign v$Y_6733_out0 = v$_6534_out0;
assign v$Y_6734_out0 = v$_6535_out0;
assign v$Y_6735_out0 = v$_6536_out0;
assign v$Y_6736_out0 = v$_6537_out0;
assign v$Y_6749_out0 = v$_6550_out0;
assign v$Y_6750_out0 = v$_6551_out0;
assign v$Y_6751_out0 = v$_6552_out0;
assign v$Y_6752_out0 = v$_6553_out0;
assign v$Y_6753_out0 = v$_6554_out0;
assign v$Y_6754_out0 = v$_6555_out0;
assign v$G1_15191_out0 = v$Z1_6049_out0 && v$Z2_180_out0;
assign v$G1_15192_out0 = v$Z1_6050_out0 && v$Z2_181_out0;
assign v$G1_15193_out0 = v$Z1_6051_out0 && v$Z2_182_out0;
assign v$G1_15196_out0 = v$Z1_6054_out0 && v$Z2_185_out0;
assign v$G1_15197_out0 = v$Z1_6055_out0 && v$Z2_186_out0;
assign v$G1_15198_out0 = v$Z1_6056_out0 && v$Z2_187_out0;
assign v$_5705_out0 = { v$Y_6732_out0,v$C1_18266_out0 };
assign v$_5706_out0 = { v$Y_6734_out0,v$C1_18267_out0 };
assign v$_5707_out0 = { v$Y_6736_out0,v$C1_18268_out0 };
assign v$_5710_out0 = { v$Y_6750_out0,v$C1_18271_out0 };
assign v$_5711_out0 = { v$Y_6752_out0,v$C1_18272_out0 };
assign v$_5712_out0 = { v$Y_6754_out0,v$C1_18273_out0 };
assign v$_8453_out0 = { v$Y_6731_out0,v$C2_7951_out0 };
assign v$_8454_out0 = { v$Y_6733_out0,v$C2_7952_out0 };
assign v$_8455_out0 = { v$Y_6735_out0,v$C2_7953_out0 };
assign v$_8458_out0 = { v$Y_6749_out0,v$C2_7956_out0 };
assign v$_8459_out0 = { v$Y_6751_out0,v$C2_7957_out0 };
assign v$_8460_out0 = { v$Y_6753_out0,v$C2_7958_out0 };
assign v$Z_10787_out0 = v$G1_15191_out0;
assign v$Z_10788_out0 = v$G1_15192_out0;
assign v$Z_10789_out0 = v$G1_15193_out0;
assign v$Z_10792_out0 = v$G1_15196_out0;
assign v$Z_10793_out0 = v$G1_15197_out0;
assign v$Z_10794_out0 = v$G1_15198_out0;
assign v$Z2_2463_out0 = v$Z_10788_out0;
assign v$Z2_2464_out0 = v$Z_10793_out0;
assign v$Z3_12563_out0 = v$Z_10787_out0;
assign v$Z3_12564_out0 = v$Z_10792_out0;
assign v$MUX1_15297_out0 = v$Z1_6049_out0 ? v$_8453_out0 : v$_5705_out0;
assign v$MUX1_15298_out0 = v$Z1_6050_out0 ? v$_8454_out0 : v$_5706_out0;
assign v$MUX1_15299_out0 = v$Z1_6051_out0 ? v$_8455_out0 : v$_5707_out0;
assign v$MUX1_15302_out0 = v$Z1_6054_out0 ? v$_8458_out0 : v$_5710_out0;
assign v$MUX1_15303_out0 = v$Z1_6055_out0 ? v$_8459_out0 : v$_5711_out0;
assign v$MUX1_15304_out0 = v$Z1_6056_out0 ? v$_8460_out0 : v$_5712_out0;
assign v$Z1_18330_out0 = v$Z_10789_out0;
assign v$Z1_18331_out0 = v$Z_10794_out0;
assign v$Y_8074_out0 = v$MUX1_15297_out0;
assign v$Y_8075_out0 = v$MUX1_15298_out0;
assign v$Y_8076_out0 = v$MUX1_15299_out0;
assign v$Y_8079_out0 = v$MUX1_15302_out0;
assign v$Y_8080_out0 = v$MUX1_15303_out0;
assign v$Y_8081_out0 = v$MUX1_15304_out0;
assign v$G2_16466_out0 = v$Z2_2463_out0 && v$Z3_12563_out0;
assign v$G2_16467_out0 = v$Z2_2464_out0 && v$Z3_12564_out0;
assign v$_1487_out0 = { v$Y_8076_out0,v$C1_8041_out0 };
assign v$_1488_out0 = { v$Y_8081_out0,v$C1_8042_out0 };
assign v$_2872_out0 = { v$Y_8075_out0,v$C2_13971_out0 };
assign v$_2873_out0 = { v$Y_8080_out0,v$C2_13972_out0 };
assign v$_3551_out0 = { v$Y_8074_out0,v$C4_16916_out0 };
assign v$_3552_out0 = { v$Y_8079_out0,v$C4_16917_out0 };
assign v$G1_17610_out0 = v$Z1_18330_out0 && v$G2_16466_out0;
assign v$G1_17611_out0 = v$Z1_18331_out0 && v$G2_16467_out0;
assign v$Z_14128_out0 = v$G1_17610_out0;
assign v$Z_14129_out0 = v$G1_17611_out0;
assign v$MUX1_15871_out0 = v$Z2_2463_out0 ? v$_1487_out0 : v$_2872_out0;
assign v$MUX1_15872_out0 = v$Z2_2464_out0 ? v$_1488_out0 : v$_2873_out0;
assign v$MUX2_14121_out0 = v$Z3_12563_out0 ? v$MUX1_15871_out0 : v$_3551_out0;
assign v$MUX2_14122_out0 = v$Z3_12564_out0 ? v$MUX1_15872_out0 : v$_3552_out0;
assign v$IS$SUM$0_16216_out0 = v$Z_14128_out0;
assign v$IS$SUM$0_16217_out0 = v$Z_14129_out0;
assign v$OUT_9253_out0 = v$MUX2_14121_out0;
assign v$OUT_9254_out0 = v$MUX2_14122_out0;
assign v$IS$SUM$0_16276_out0 = v$IS$SUM$0_16216_out0;
assign v$IS$SUM$0_16277_out0 = v$IS$SUM$0_16217_out0;
assign v$IS$SUM$0_1000_out0 = v$IS$SUM$0_16276_out0;
assign v$IS$SUM$0_1001_out0 = v$IS$SUM$0_16277_out0;
assign v$_10833_out0 = { v$OUT_9253_out0,v$C10_14117_out0 };
assign v$_10834_out0 = { v$OUT_9254_out0,v$C10_14118_out0 };
assign v$NORMALIZATION$SHIFT_3477_out0 = v$_10833_out0;
assign v$NORMALIZATION$SHIFT_3478_out0 = v$_10834_out0;
assign v$NORMALIZATION$SHIFT_1311_out0 = v$NORMALIZATION$SHIFT_3477_out0;
assign v$NORMALIZATION$SHIFT_1312_out0 = v$NORMALIZATION$SHIFT_3478_out0;
assign v$SHIFT$AMOUNT_7704_out0 = v$NORMALIZATION$SHIFT_3477_out0;
assign v$SHIFT$AMOUNT_7708_out0 = v$NORMALIZATION$SHIFT_3478_out0;
assign v$SEL3_1283_out0 = v$SHIFT$AMOUNT_7704_out0[2:2];
assign v$SEL3_1287_out0 = v$SHIFT$AMOUNT_7708_out0[2:2];
assign v$SEL1_2477_out0 = v$SHIFT$AMOUNT_7704_out0[0:0];
assign v$SEL1_2481_out0 = v$SHIFT$AMOUNT_7708_out0[0:0];
assign v$SEL4_5154_out0 = v$SHIFT$AMOUNT_7704_out0[3:3];
assign v$SEL4_5158_out0 = v$SHIFT$AMOUNT_7708_out0[3:3];
assign v$SEL7_6598_out0 = v$SHIFT$AMOUNT_7704_out0[5:5];
assign v$SEL7_6602_out0 = v$SHIFT$AMOUNT_7708_out0[5:5];
assign v$SEL5_12783_out0 = v$SHIFT$AMOUNT_7704_out0[4:4];
assign v$SEL5_12787_out0 = v$SHIFT$AMOUNT_7708_out0[4:4];
assign v$SEL6_14367_out0 = v$SHIFT$AMOUNT_7704_out0[6:6];
assign v$SEL6_14371_out0 = v$SHIFT$AMOUNT_7708_out0[6:6];
assign v$SEL8_17192_out0 = v$SHIFT$AMOUNT_7704_out0[7:7];
assign v$SEL8_17196_out0 = v$SHIFT$AMOUNT_7708_out0[7:7];
assign v$SEL2_18962_out0 = v$SHIFT$AMOUNT_7704_out0[1:1];
assign v$SEL2_18966_out0 = v$SHIFT$AMOUNT_7708_out0[1:1];
assign v$NORMALIZATION$SHIFT_19233_out0 = v$NORMALIZATION$SHIFT_1311_out0;
assign v$NORMALIZATION$SHIFT_19234_out0 = v$NORMALIZATION$SHIFT_1312_out0;
assign v$EN_1497_out0 = v$SEL5_12783_out0;
assign v$EN_1498_out0 = v$SEL4_5154_out0;
assign v$EN_1507_out0 = v$SEL5_12787_out0;
assign v$EN_1508_out0 = v$SEL4_5158_out0;
assign v$EN_4965_out0 = v$SEL3_1283_out0;
assign v$EN_4971_out0 = v$SEL3_1287_out0;
assign v$EN_5429_out0 = v$SEL1_2477_out0;
assign v$EN_5435_out0 = v$SEL1_2481_out0;
assign v$EN_8201_out0 = v$SEL2_18962_out0;
assign v$EN_8207_out0 = v$SEL2_18966_out0;
assign v$SEL14_9427_out0 = v$NORMALIZATION$SHIFT_19233_out0[4:0];
assign v$SEL14_9428_out0 = v$NORMALIZATION$SHIFT_19234_out0[4:0];
assign v$NORMALIZATION$SHIFT_11230_out0 = v$NORMALIZATION$SHIFT_19233_out0;
assign v$NORMALIZATION$SHIFT_11231_out0 = v$NORMALIZATION$SHIFT_19234_out0;
assign v$G1_16645_out0 = v$SEL7_6598_out0 || v$SEL6_14367_out0;
assign v$G1_16649_out0 = v$SEL7_6602_out0 || v$SEL6_14371_out0;
assign v$NORMALIZATION$SHIFT_4562_out0 = v$SEL14_9427_out0;
assign v$NORMALIZATION$SHIFT_4563_out0 = v$SEL14_9428_out0;
assign v$XOR1_15146_out0 = v$NORMALIZATION$SHIFT_11230_out0 ^ v$C1_1711_out0;
assign v$XOR1_15147_out0 = v$NORMALIZATION$SHIFT_11231_out0 ^ v$C1_1712_out0;
assign v$G2_18056_out0 = v$G1_16645_out0 || v$SEL8_17192_out0;
assign v$G2_18060_out0 = v$G1_16649_out0 || v$SEL8_17196_out0;
assign v$MUX2_19187_out0 = v$EN_5429_out0 ? v$MUX1_2555_out0 : v$IN_4038_out0;
assign v$MUX2_19193_out0 = v$EN_5435_out0 ? v$MUX1_2586_out0 : v$IN_4047_out0;
assign {v$A1_698_out1,v$A1_698_out0 } = v$EXPONENT_1521_out0 + v$XOR1_15146_out0 + v$C2_3185_out0;
assign {v$A1_699_out1,v$A1_699_out0 } = v$EXPONENT_1522_out0 + v$XOR1_15147_out0 + v$C2_3186_out0;
assign v$XOR1_11435_out0 = v$NORMALIZATION$SHIFT_4562_out0 ^ v$C1_16332_out0;
assign v$XOR1_11436_out0 = v$NORMALIZATION$SHIFT_4563_out0 ^ v$C1_16333_out0;
assign v$OUT_15527_out0 = v$MUX2_19187_out0;
assign v$OUT_15558_out0 = v$MUX2_19193_out0;
assign v$IN_5379_out0 = v$OUT_15527_out0;
assign v$IN_5410_out0 = v$OUT_15558_out0;
assign {v$A1_8047_out1,v$A1_8047_out0 } = v$EXPONENT_17014_out0 + v$XOR1_11435_out0 + v$C2_1607_out0;
assign {v$A1_8048_out1,v$A1_8048_out0 } = v$EXPONENT_17015_out0 + v$XOR1_11436_out0 + v$C2_1608_out0;
assign v$IGNORE_12272_out0 = v$A1_698_out1;
assign v$IGNORE_12273_out0 = v$A1_699_out1;
assign v$OUT_16707_out0 = v$A1_698_out0;
assign v$OUT_16708_out0 = v$A1_699_out0;
assign v$OUT_6454_out0 = v$A1_8047_out0;
assign v$OUT_6455_out0 = v$A1_8048_out0;
assign v$IN_12354_out0 = v$IN_5379_out0;
assign v$IN_12360_out0 = v$IN_5410_out0;
assign v$IGNORE_17180_out0 = v$A1_8047_out1;
assign v$IGNORE_17181_out0 = v$A1_8048_out1;
assign v$SEL1_9060_out0 = v$IN_12354_out0[23:2];
assign v$SEL1_9091_out0 = v$IN_12360_out0[23:2];
assign v$SEL1_15988_out0 = v$IN_12354_out0[21:0];
assign v$SEL1_16019_out0 = v$IN_12360_out0[21:0];
assign v$_4420_out0 = { v$C2_118_out0,v$SEL1_15988_out0 };
assign v$_4451_out0 = { v$C2_149_out0,v$SEL1_16019_out0 };
assign v$_9321_out0 = { v$SEL1_9060_out0,v$C1_6256_out0 };
assign v$_9352_out0 = { v$SEL1_9091_out0,v$C1_6287_out0 };
assign v$MUX1_2557_out0 = v$LEFT$SHIT_3269_out0 ? v$_4420_out0 : v$_9321_out0;
assign v$MUX1_2588_out0 = v$LEFT$SHIT_3300_out0 ? v$_4451_out0 : v$_9352_out0;
assign v$MUX2_2672_out0 = v$EN_8201_out0 ? v$MUX1_2557_out0 : v$IN_12354_out0;
assign v$MUX2_2678_out0 = v$EN_8207_out0 ? v$MUX1_2588_out0 : v$IN_12360_out0;
assign v$OUT_15529_out0 = v$MUX2_2672_out0;
assign v$OUT_15560_out0 = v$MUX2_2678_out0;
assign v$IN_5378_out0 = v$OUT_15529_out0;
assign v$IN_5409_out0 = v$OUT_15560_out0;
assign v$IN_16198_out0 = v$IN_5378_out0;
assign v$IN_16204_out0 = v$IN_5409_out0;
assign v$SEL1_9059_out0 = v$IN_16198_out0[23:4];
assign v$SEL1_9090_out0 = v$IN_16204_out0[23:4];
assign v$SEL1_15987_out0 = v$IN_16198_out0[19:0];
assign v$SEL1_16018_out0 = v$IN_16204_out0[19:0];
assign v$_4419_out0 = { v$C2_117_out0,v$SEL1_15987_out0 };
assign v$_4450_out0 = { v$C2_148_out0,v$SEL1_16018_out0 };
assign v$_9320_out0 = { v$SEL1_9059_out0,v$C1_6255_out0 };
assign v$_9351_out0 = { v$SEL1_9090_out0,v$C1_6286_out0 };
assign v$MUX1_2556_out0 = v$LEFT$SHIT_3268_out0 ? v$_4419_out0 : v$_9320_out0;
assign v$MUX1_2587_out0 = v$LEFT$SHIT_3299_out0 ? v$_4450_out0 : v$_9351_out0;
assign v$MUX2_15819_out0 = v$EN_4965_out0 ? v$MUX1_2556_out0 : v$IN_16198_out0;
assign v$MUX2_15825_out0 = v$EN_4971_out0 ? v$MUX1_2587_out0 : v$IN_16204_out0;
assign v$OUT_15528_out0 = v$MUX2_15819_out0;
assign v$OUT_15559_out0 = v$MUX2_15825_out0;
assign v$IN_5376_out0 = v$OUT_15528_out0;
assign v$IN_5407_out0 = v$OUT_15559_out0;
assign v$IN_5238_out0 = v$IN_5376_out0;
assign v$IN_5248_out0 = v$IN_5407_out0;
assign v$SEL1_9057_out0 = v$IN_5238_out0[23:8];
assign v$SEL1_9088_out0 = v$IN_5248_out0[23:8];
assign v$SEL1_15985_out0 = v$IN_5238_out0[15:0];
assign v$SEL1_16016_out0 = v$IN_5248_out0[15:0];
assign v$_4417_out0 = { v$C2_115_out0,v$SEL1_15985_out0 };
assign v$_4448_out0 = { v$C2_146_out0,v$SEL1_16016_out0 };
assign v$_9318_out0 = { v$SEL1_9057_out0,v$C1_6253_out0 };
assign v$_9349_out0 = { v$SEL1_9088_out0,v$C1_6284_out0 };
assign v$MUX1_2554_out0 = v$LEFT$SHIT_3266_out0 ? v$_4417_out0 : v$_9318_out0;
assign v$MUX1_2585_out0 = v$LEFT$SHIT_3297_out0 ? v$_4448_out0 : v$_9349_out0;
assign v$MUX2_2693_out0 = v$EN_1498_out0 ? v$MUX1_2554_out0 : v$IN_5238_out0;
assign v$MUX2_2703_out0 = v$EN_1508_out0 ? v$MUX1_2585_out0 : v$IN_5248_out0;
assign v$OUT_15526_out0 = v$MUX2_2693_out0;
assign v$OUT_15557_out0 = v$MUX2_2703_out0;
assign v$IN_5375_out0 = v$OUT_15526_out0;
assign v$IN_5406_out0 = v$OUT_15557_out0;
assign v$IN_5237_out0 = v$IN_5375_out0;
assign v$IN_5247_out0 = v$IN_5406_out0;
assign v$SEL1_9056_out0 = v$IN_5237_out0[23:16];
assign v$SEL1_9087_out0 = v$IN_5247_out0[23:16];
assign v$SEL1_15984_out0 = v$IN_5237_out0[7:0];
assign v$SEL1_16015_out0 = v$IN_5247_out0[7:0];
assign v$_4416_out0 = { v$C2_114_out0,v$SEL1_15984_out0 };
assign v$_4447_out0 = { v$C2_145_out0,v$SEL1_16015_out0 };
assign v$_9317_out0 = { v$SEL1_9056_out0,v$C1_6252_out0 };
assign v$_9348_out0 = { v$SEL1_9087_out0,v$C1_6283_out0 };
assign v$MUX1_2553_out0 = v$LEFT$SHIT_3265_out0 ? v$_4416_out0 : v$_9317_out0;
assign v$MUX1_2584_out0 = v$LEFT$SHIT_3296_out0 ? v$_4447_out0 : v$_9348_out0;
assign v$MUX2_2692_out0 = v$EN_1497_out0 ? v$MUX1_2553_out0 : v$IN_5237_out0;
assign v$MUX2_2702_out0 = v$EN_1507_out0 ? v$MUX1_2584_out0 : v$IN_5247_out0;
assign v$OUT_15525_out0 = v$MUX2_2692_out0;
assign v$OUT_15556_out0 = v$MUX2_2702_out0;
assign v$MUX1_12193_out0 = v$G2_18056_out0 ? v$C1_4625_out0 : v$OUT_15525_out0;
assign v$MUX1_12197_out0 = v$G2_18060_out0 ? v$C1_4629_out0 : v$OUT_15556_out0;
assign v$OUT_10438_out0 = v$MUX1_12193_out0;
assign v$OUT_10442_out0 = v$MUX1_12197_out0;
assign v$SEL2_6314_out0 = v$OUT_10438_out0[22:0];
assign v$SEL2_6315_out0 = v$OUT_10442_out0[22:0];
assign v$MUX2_3183_out0 = v$IS$SUM$0_16216_out0 ? v$C5_16212_out0 : v$SEL2_6314_out0;
assign v$MUX2_3184_out0 = v$IS$SUM$0_16217_out0 ? v$C5_16213_out0 : v$SEL2_6315_out0;
assign v$MUX6_13339_out0 = v$IS$SUB_13643_out0 ? v$MUX2_3183_out0 : v$SEL3_14851_out0;
assign v$MUX6_13340_out0 = v$IS$SUB_13644_out0 ? v$MUX2_3184_out0 : v$SEL3_14852_out0;
assign v$OUT1_10858_out0 = v$MUX6_13339_out0;
assign v$OUT1_10859_out0 = v$MUX6_13340_out0;
assign v$MANTISA$RESULT_6779_out0 = v$OUT1_10858_out0;
assign v$MANTISA$RESULT_6780_out0 = v$OUT1_10859_out0;
assign v$SEL10_3429_out0 = v$MANTISA$RESULT_6779_out0[22:13];
assign v$SEL10_3430_out0 = v$MANTISA$RESULT_6780_out0[22:13];
assign v$SEL7_3499_out0 = v$MANTISA$RESULT_6779_out0[22:13];
assign v$SEL7_3500_out0 = v$MANTISA$RESULT_6780_out0[22:13];
assign v$_7305_out0 = { v$MANTISA$RESULT_6779_out0,v$OUT_15386_out0 };
assign v$_7306_out0 = { v$MANTISA$RESULT_6780_out0,v$OUT_15387_out0 };
assign v$_15939_out0 = { v$MANTISA$RESULT_6779_out0,v$OUT_16707_out0 };
assign v$_15940_out0 = { v$MANTISA$RESULT_6780_out0,v$OUT_16708_out0 };
assign v$_11912_out0 = { v$SEL10_3429_out0,v$OUT_6454_out0 };
assign v$_11913_out0 = { v$SEL10_3430_out0,v$OUT_6455_out0 };
assign v$_15764_out0 = { v$SEL7_3499_out0,v$OUT_170_out0 };
assign v$_15765_out0 = { v$SEL7_3500_out0,v$OUT_171_out0 };
assign v$_58_out0 = { v$C9_3525_out0,v$_11912_out0 };
assign v$_59_out0 = { v$C9_3526_out0,v$_11913_out0 };
assign v$_12403_out0 = { v$C7_1867_out0,v$_15764_out0 };
assign v$_12404_out0 = { v$C7_1868_out0,v$_15765_out0 };
assign v$MUX12_15750_out0 = v$IS$32$BIT_11362_out0 ? v$_7305_out0 : v$_12403_out0;
assign v$MUX12_15751_out0 = v$IS$32$BIT_11363_out0 ? v$_7306_out0 : v$_12404_out0;
assign v$MUX6_18078_out0 = v$IS$32$BIT_11362_out0 ? v$_15939_out0 : v$_58_out0;
assign v$MUX6_18079_out0 = v$IS$32$BIT_11363_out0 ? v$_15940_out0 : v$_59_out0;
assign v$_17132_out0 = { v$MUX12_15750_out0,v$SEL13_18204_out0 };
assign v$_17133_out0 = { v$MUX12_15751_out0,v$SEL13_18205_out0 };
assign v$_17422_out0 = { v$MUX6_18078_out0,v$SUBTRACTION$SIGN_12445_out0 };
assign v$_17423_out0 = { v$MUX6_18079_out0,v$SUBTRACTION$SIGN_12446_out0 };
assign v$MUX1_14132_out0 = v$IS$SUB_4611_out0 ? v$_17422_out0 : v$_17132_out0;
assign v$MUX1_14133_out0 = v$IS$SUB_4612_out0 ? v$_17423_out0 : v$_17133_out0;
assign v$MUX7_5078_out0 = v$IS$SUM$0_1000_out0 ? v$C5_4269_out0 : v$MUX1_14132_out0;
assign v$MUX7_5079_out0 = v$IS$SUM$0_1001_out0 ? v$C5_4270_out0 : v$MUX1_14133_out0;
assign v$OUT1_18415_out0 = v$MUX7_5078_out0;
assign v$OUT1_18416_out0 = v$MUX7_5079_out0;
assign v$MUX2_16839_out0 = v$G2_3905_out0 ? v$OUT1_18415_out0 : v$C4_14636_out0;
assign v$MUX2_16840_out0 = v$G2_3906_out0 ? v$OUT1_18416_out0 : v$C4_14637_out0;
assign v$MUX4_1411_out0 = v$FINISHED_8327_out0 ? v$OUT_3588_out0 : v$MUX2_16839_out0;
assign v$MUX4_1412_out0 = v$FINISHED_8328_out0 ? v$OUT_3589_out0 : v$MUX2_16840_out0;
assign v$SEL4_9936_out0 = v$MUX4_1411_out0[15:0];
assign v$SEL4_9937_out0 = v$MUX4_1412_out0[15:0];
assign v$SEL5_14164_out0 = v$MUX4_1411_out0[31:16];
assign v$SEL5_14165_out0 = v$MUX4_1412_out0[31:16];
assign v$MUX3_18992_out0 = v$G12_12555_out0 ? v$REG3_12336_out0 : v$SEL5_14164_out0;
assign v$MUX3_18993_out0 = v$G12_12556_out0 ? v$REG3_12337_out0 : v$SEL5_14165_out0;
assign v$OUT_1483_out0 = v$MUX3_18992_out0;
assign v$OUT_1484_out0 = v$MUX3_18993_out0;
assign v$FPU$OUT_17605_out0 = v$OUT_1483_out0;
assign v$FPU$OUT_17606_out0 = v$OUT_1484_out0;
assign v$MUX6_7758_out0 = v$G21_19292_out0 ? v$FPU$OUT_17605_out0 : v$MUX4_46_out0;
assign v$MUX6_7759_out0 = v$G21_19293_out0 ? v$FPU$OUT_17606_out0 : v$MUX4_47_out0;
assign v$MUX14_19331_out0 = v$FINISHED_14451_out0 ? v$FPU$OUT_17605_out0 : v$MUX6_7758_out0;
assign v$MUX14_19332_out0 = v$FINISHED_14452_out0 ? v$FPU$OUT_17606_out0 : v$MUX6_7759_out0;
assign v$DIN3_15022_out0 = v$MUX14_19331_out0;
assign v$DIN3_15023_out0 = v$MUX14_19332_out0;


endmodule

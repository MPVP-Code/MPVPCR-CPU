

    module v$RAM1_8558(q, a, d, we, clk);
    output reg [15:0] q;
    input [15:0] d;
    input [11:0] a;
    input we, clk;
    reg [15:0] ram [4095:0];
     always @(posedge clk) begin
         if (we)
             ram[a] <= d;
         q <= ram[a];
     end

    integer i;
    initial
    begin
        for (i=0; i < 4096; i=i+1)
        begin
            ram[i] = 0;
        end

        ram[0] = 16;
ram[1] = 32;
ram[2] = 48;
ram[3] = 64;
ram[4] = 80;
    end
    endmodule

    

    module v$AROM1_11322(q, a);
    output[43:0] q;
    input [5:0] a;
    reg [43:0] rom [63:0];

    assign q = rom[a];
    integer i;
    initial
    begin
        for (i=0; i < 64; i=i+1)
        begin
            rom[i] = 0;
        end
    
        rom[0] = 1030792151295;
rom[1] = 64424509695;
rom[2] = 1095216660735;
rom[3] = 4026532095;
rom[4] = 1034818683135;
rom[5] = 68451041535;
rom[6] = 1099243192575;
rom[7] = 251658495;
rom[8] = 1031043809535;
rom[9] = 64676167935;
rom[10] = 0;
    end
    endmodule
     

    module v$AROM1_11323(q, a);
    output[43:0] q;
    input [5:0] a;
    reg [43:0] rom [63:0];

    assign q = rom[a];
    integer i;
    initial
    begin
        for (i=0; i < 64; i=i+1)
        begin
            rom[i] = 0;
        end
    
        rom[0] = 1030792151295;
rom[1] = 64424509695;
rom[2] = 1095216660735;
rom[3] = 4026532095;
rom[4] = 1034818683135;
rom[5] = 68451041535;
rom[6] = 1099243192575;
rom[7] = 251658495;
rom[8] = 1031043809535;
rom[9] = 64676167935;
rom[10] = 0;
    end
    endmodule
     

    module v$ROM1_12254(q, a, clk);
    output reg [15:0] q;
    input clk;
    input [11:0] a;
    reg [15:0] rom [4095:0];
    always @(posedge clk) q <= rom[a];
    integer i;
    initial
    begin
        for (i=0; i < 4096; i=i+1)
        begin
            rom[i] = 0;
        end
    
        rom[0] = 52740;
rom[1] = 1860;
rom[2] = 34817;
rom[3] = 53251;
rom[4] = 20481;
rom[5] = 51238;
rom[6] = 52752;
rom[7] = 2115;
rom[8] = 28672;
rom[9] = 7713;
rom[10] = 6912;
rom[11] = 7104;
rom[12] = 7713;
rom[13] = 6912;
rom[14] = 7040;
rom[15] = 5411;
rom[16] = 4864;
rom[17] = 52740;
rom[18] = 327;
rom[19] = 1027;
rom[20] = 52736;
rom[21] = 839;
rom[22] = 4992;
rom[23] = 1863;
rom[24] = 52742;
rom[25] = 2887;
rom[26] = 7104;
rom[27] = 3587;
rom[28] = 7713;
rom[29] = 6912;
rom[30] = 7104;
rom[31] = 7713;
rom[32] = 6912;
rom[33] = 7104;
rom[34] = 7713;
rom[35] = 6912;
rom[36] = 7104;
rom[37] = 7713;
rom[38] = 6912;
rom[39] = 7104;
rom[40] = 7713;
rom[41] = 6912;
rom[42] = 50692;
rom[43] = 837;
rom[44] = 1537;
rom[45] = 5056;
rom[46] = 7040;
rom[47] = 5155;
rom[48] = 4864;
rom[49] = 52744;
rom[50] = 327;
rom[51] = 1027;
rom[52] = 52736;
rom[53] = 839;
rom[54] = 4992;
rom[55] = 1863;
rom[56] = 52746;
rom[57] = 2887;
rom[58] = 7104;
rom[59] = 3587;
rom[60] = 7713;
rom[61] = 6912;
rom[62] = 7104;
rom[63] = 7713;
rom[64] = 6912;
rom[65] = 7104;
rom[66] = 7713;
rom[67] = 6912;
rom[68] = 7104;
rom[69] = 7713;
rom[70] = 6912;
rom[71] = 7104;
rom[72] = 7713;
rom[73] = 6912;
rom[74] = 7104;
rom[75] = 7713;
rom[76] = 6912;
rom[77] = 7104;
rom[78] = 7713;
rom[79] = 6912;
rom[80] = 50696;
rom[81] = 837;
rom[82] = 1537;
rom[83] = 5056;
rom[84] = 7040;
rom[85] = 5411;
rom[86] = 4864;
rom[87] = 52748;
rom[88] = 327;
rom[89] = 1027;
rom[90] = 28672;
    end
    endmodule
     

    module v$ROM1_12255(q, a, clk);
    output reg [15:0] q;
    input clk;
    input [11:0] a;
    reg [15:0] rom [4095:0];
    always @(posedge clk) q <= rom[a];
    integer i;
    initial
    begin
        for (i=0; i < 4096; i=i+1)
        begin
            rom[i] = 0;
        end
    
        rom[0] = 52744;
rom[1] = 516;
rom[2] = 1860;
rom[3] = 34817;
rom[4] = 53251;
rom[5] = 20482;
rom[6] = 51238;
rom[7] = 52752;
rom[8] = 1603;
rom[9] = 35073;
rom[10] = 51222;
rom[11] = 2115;
rom[12] = 28672;
    end
    endmodule
     
module main (
	clk);
input clk;
reg  [11:0] v$INT0_11100_out0 = 12'h0;
reg  [11:0] v$INT0_11101_out0 = 12'h0;
reg  [11:0] v$INT1_13185_out0 = 12'h0;
reg  [11:0] v$INT1_13186_out0 = 12'h0;
reg  [11:0] v$INT2_221_out0 = 12'h0;
reg  [11:0] v$INT2_222_out0 = 12'h0;
reg  [11:0] v$INT3_233_out0 = 12'h0;
reg  [11:0] v$INT3_234_out0 = 12'h0;
reg  [11:0] v$PCINTERRUPT_12603_out0 = 12'h0;
reg  [11:0] v$PCINTERRUPT_12604_out0 = 12'h0;
reg  [11:0] v$PCNORMAL_8422_out0 = 12'h0;
reg  [11:0] v$PCNORMAL_8423_out0 = 12'h0;
reg  [11:0] v$REG12_2023_out0 = 12'h0;
reg  [11:0] v$REG9_11269_out0 = 12'h0;
reg  [15:0] v$REG0_11406_out0 = 16'h0;
reg  [15:0] v$REG0_11407_out0 = 16'h0;
reg  [15:0] v$REG10_11541_out0 = 16'h0;
reg  [15:0] v$REG11_6578_out0 = 16'h0;
reg  [15:0] v$REG1_3286_out0 = 16'h0;
reg  [15:0] v$REG1_3287_out0 = 16'h0;
reg  [15:0] v$REG1_457_out0 = 16'h0;
reg  [15:0] v$REG1_458_out0 = 16'h0;
reg  [15:0] v$REG1_9161_out0 = 16'h0;
reg  [15:0] v$REG1_9162_out0 = 16'h0;
reg  [15:0] v$REG1_9488_out0 = 16'h0;
reg  [15:0] v$REG1_9489_out0 = 16'h0;
reg  [15:0] v$REG2_10321_out0 = 16'h0;
reg  [15:0] v$REG2_10322_out0 = 16'h0;
reg  [15:0] v$REG2_10886_out0 = 16'h0;
reg  [15:0] v$REG2_10887_out0 = 16'h0;
reg  [15:0] v$REG2_11460_out0 = 16'h0;
reg  [15:0] v$REG2_11461_out0 = 16'h0;
reg  [15:0] v$REG2_12278_out0 = 16'h0;
reg  [15:0] v$REG2_12279_out0 = 16'h0;
reg  [15:0] v$REG3_1589_out0 = 16'h0;
reg  [15:0] v$REG3_1590_out0 = 16'h0;
reg  [15:0] v$REG3_7255_out0 = 16'h0;
reg  [15:0] v$REG3_7256_out0 = 16'h0;
reg  [15:0] v$REG3_7578_out0 = 16'h0;
reg  [15:0] v$REG3_7579_out0 = 16'h0;
reg  [15:0] v$REG4_4650_out0 = 16'h0;
reg  [15:0] v$REG4_4651_out0 = 16'h0;
reg  [1:0] v$REG1_7183_out0 = 2'h0;
reg  [1:0] v$REG1_7184_out0 = 2'h0;
reg  [35:0] v$REG3_4759_out0 = 36'h0;
reg  [35:0] v$REG3_4760_out0 = 36'h0;
reg  [3:0] v$REG1_13298_out0 = 4'h0;
reg  [3:0] v$REG1_13299_out0 = 4'h0;
reg  [3:0] v$REG1_6141_out0 = 4'h0;
reg  [3:0] v$REG1_6142_out0 = 4'h0;
reg  [5:0] v$REG1_10179_out0 = 6'h0;
reg  [5:0] v$REG1_10180_out0 = 6'h0;
reg  [5:0] v$REG2_376_out0 = 6'h0;
reg  [5:0] v$REG2_377_out0 = 6'h0;
reg  [7:0] v$REG1_2760_out0 = 8'h0;
reg  [7:0] v$REG1_2761_out0 = 8'h0;
reg  [7:0] v$REG1_6863_out0 = 8'h0;
reg  [7:0] v$REG1_6864_out0 = 8'h0;
reg v$FF0_2992_out0 = 1'b0;
reg v$FF0_2993_out0 = 1'b0;
reg v$FF0_3399_out0 = 1'b0;
reg v$FF0_3400_out0 = 1'b0;
reg v$FF0_374_out0 = 1'b0;
reg v$FF0_375_out0 = 1'b0;
reg v$FF0_6397_out0 = 1'b0;
reg v$FF0_6398_out0 = 1'b0;
reg v$FF10_5406_out0 = 1'b0;
reg v$FF10_5407_out0 = 1'b0;
reg v$FF10_9601_out0 = 1'b0;
reg v$FF10_9602_out0 = 1'b0;
reg v$FF11_1377_out0 = 1'b0;
reg v$FF11_1378_out0 = 1'b0;
reg v$FF12_11522_out0 = 1'b0;
reg v$FF12_11523_out0 = 1'b0;
reg v$FF13_13193_out0 = 1'b0;
reg v$FF13_13194_out0 = 1'b0;
reg v$FF14_7185_out0 = 1'b0;
reg v$FF14_7186_out0 = 1'b0;
reg v$FF15_8373_out0 = 1'b0;
reg v$FF15_8374_out0 = 1'b0;
reg v$FF1_11255_out0 = 1'b0;
reg v$FF1_11256_out0 = 1'b0;
reg v$FF1_11257_out0 = 1'b0;
reg v$FF1_11258_out0 = 1'b0;
reg v$FF1_11259_out0 = 1'b0;
reg v$FF1_11260_out0 = 1'b0;
reg v$FF1_11261_out0 = 1'b0;
reg v$FF1_11262_out0 = 1'b0;
reg v$FF1_11263_out0 = 1'b0;
reg v$FF1_11264_out0 = 1'b0;
reg v$FF1_11265_out0 = 1'b0;
reg v$FF1_11266_out0 = 1'b0;
reg v$FF1_11343_out0 = 1'b0;
reg v$FF1_11344_out0 = 1'b0;
reg v$FF1_11440_out0 = 1'b0;
reg v$FF1_11441_out0 = 1'b0;
reg v$FF1_1433_out0 = 1'b0;
reg v$FF1_1434_out0 = 1'b0;
reg v$FF1_178_out0 = 1'b0;
reg v$FF1_179_out0 = 1'b0;
reg v$FF1_2_out0 = 1'b0;
reg v$FF1_3605_out0 = 1'b0;
reg v$FF1_3606_out0 = 1'b0;
reg v$FF1_3695_out0 = 1'b0;
reg v$FF1_3_out0 = 1'b0;
reg v$FF1_4029_out0 = 1'b0;
reg v$FF1_4030_out0 = 1'b0;
reg v$FF1_4163_out0 = 1'b0;
reg v$FF1_4164_out0 = 1'b0;
reg v$FF1_467_out0 = 1'b0;
reg v$FF1_468_out0 = 1'b0;
reg v$FF1_5716_out0 = 1'b0;
reg v$FF1_5717_out0 = 1'b0;
reg v$FF1_601_out0 = 1'b0;
reg v$FF1_602_out0 = 1'b0;
reg v$FF1_6417_out0 = 1'b0;
reg v$FF1_6418_out0 = 1'b0;
reg v$FF1_6568_out0 = 1'b0;
reg v$FF1_6569_out0 = 1'b0;
reg v$FF1_6586_out0 = 1'b0;
reg v$FF1_6587_out0 = 1'b0;
reg v$FF1_6867_out0 = 1'b0;
reg v$FF1_6868_out0 = 1'b0;
reg v$FF1_7292_out0 = 1'b0;
reg v$FF1_7293_out0 = 1'b0;
reg v$FF1_8718_out0 = 1'b0;
reg v$FF1_8719_out0 = 1'b0;
reg v$FF1_9226_out0 = 1'b0;
reg v$FF1_9227_out0 = 1'b0;
reg v$FF2_10133_out0 = 1'b0;
reg v$FF2_10134_out0 = 1'b0;
reg v$FF2_10135_out0 = 1'b0;
reg v$FF2_10136_out0 = 1'b0;
reg v$FF2_10137_out0 = 1'b0;
reg v$FF2_10138_out0 = 1'b0;
reg v$FF2_10139_out0 = 1'b0;
reg v$FF2_10140_out0 = 1'b0;
reg v$FF2_10141_out0 = 1'b0;
reg v$FF2_10142_out0 = 1'b0;
reg v$FF2_10143_out0 = 1'b0;
reg v$FF2_10144_out0 = 1'b0;
reg v$FF2_10772_out0 = 1'b0;
reg v$FF2_10773_out0 = 1'b0;
reg v$FF2_11450_out0 = 1'b0;
reg v$FF2_11451_out0 = 1'b0;
reg v$FF2_11724_out0 = 1'b0;
reg v$FF2_11725_out0 = 1'b0;
reg v$FF2_1717_out0 = 1'b0;
reg v$FF2_1718_out0 = 1'b0;
reg v$FF2_3000_out0 = 1'b0;
reg v$FF2_3001_out0 = 1'b0;
reg v$FF2_469_out0 = 1'b0;
reg v$FF2_470_out0 = 1'b0;
reg v$FF2_6413_out0 = 1'b0;
reg v$FF2_6414_out0 = 1'b0;
reg v$FF2_779_out0 = 1'b0;
reg v$FF2_780_out0 = 1'b0;
reg v$FF2_8662_out0 = 1'b0;
reg v$FF2_8663_out0 = 1'b0;
reg v$FF2_8664_out0 = 1'b0;
reg v$FF2_8665_out0 = 1'b0;
reg v$FF2_8666_out0 = 1'b0;
reg v$FF2_8667_out0 = 1'b0;
reg v$FF2_8668_out0 = 1'b0;
reg v$FF2_8669_out0 = 1'b0;
reg v$FF2_8670_out0 = 1'b0;
reg v$FF2_8671_out0 = 1'b0;
reg v$FF2_8672_out0 = 1'b0;
reg v$FF2_8673_out0 = 1'b0;
reg v$FF2_8674_out0 = 1'b0;
reg v$FF2_8675_out0 = 1'b0;
reg v$FF2_8676_out0 = 1'b0;
reg v$FF2_8677_out0 = 1'b0;
reg v$FF2_8678_out0 = 1'b0;
reg v$FF2_8679_out0 = 1'b0;
reg v$FF2_8680_out0 = 1'b0;
reg v$FF2_8681_out0 = 1'b0;
reg v$FF2_8682_out0 = 1'b0;
reg v$FF2_8683_out0 = 1'b0;
reg v$FF2_9024_out0 = 1'b0;
reg v$FF2_9998_out0 = 1'b0;
reg v$FF2_9999_out0 = 1'b0;
reg v$FF3_10341_out0 = 1'b0;
reg v$FF3_10342_out0 = 1'b0;
reg v$FF3_11154_out0 = 1'b0;
reg v$FF3_11155_out0 = 1'b0;
reg v$FF3_12851_out0 = 1'b0;
reg v$FF3_12852_out0 = 1'b0;
reg v$FF3_2072_out0 = 1'b0;
reg v$FF3_227_out0 = 1'b0;
reg v$FF3_228_out0 = 1'b0;
reg v$FF3_4929_out0 = 1'b0;
reg v$FF3_4930_out0 = 1'b0;
reg v$FF3_5109_out0 = 1'b0;
reg v$FF3_5110_out0 = 1'b0;
reg v$FF3_532_out0 = 1'b0;
reg v$FF3_533_out0 = 1'b0;
reg v$FF3_6686_out0 = 1'b0;
reg v$FF3_6687_out0 = 1'b0;
reg v$FF3_6688_out0 = 1'b0;
reg v$FF3_6689_out0 = 1'b0;
reg v$FF3_6690_out0 = 1'b0;
reg v$FF3_6691_out0 = 1'b0;
reg v$FF3_6692_out0 = 1'b0;
reg v$FF3_6693_out0 = 1'b0;
reg v$FF3_6694_out0 = 1'b0;
reg v$FF3_6695_out0 = 1'b0;
reg v$FF3_6696_out0 = 1'b0;
reg v$FF3_6697_out0 = 1'b0;
reg v$FF3_7189_out0 = 1'b0;
reg v$FF3_7190_out0 = 1'b0;
reg v$FF4_11162_out0 = 1'b0;
reg v$FF4_11163_out0 = 1'b0;
reg v$FF4_11164_out0 = 1'b0;
reg v$FF4_11165_out0 = 1'b0;
reg v$FF4_11166_out0 = 1'b0;
reg v$FF4_11167_out0 = 1'b0;
reg v$FF4_11168_out0 = 1'b0;
reg v$FF4_11169_out0 = 1'b0;
reg v$FF4_11170_out0 = 1'b0;
reg v$FF4_11171_out0 = 1'b0;
reg v$FF4_11172_out0 = 1'b0;
reg v$FF4_11173_out0 = 1'b0;
reg v$FF4_12634_out0 = 1'b0;
reg v$FF4_12635_out0 = 1'b0;
reg v$FF4_1281_out0 = 1'b0;
reg v$FF4_1282_out0 = 1'b0;
reg v$FF4_13119_out0 = 1'b0;
reg v$FF4_13120_out0 = 1'b0;
reg v$FF4_2489_out0 = 1'b0;
reg v$FF4_2490_out0 = 1'b0;
reg v$FF4_4776_out0 = 1'b0;
reg v$FF4_4777_out0 = 1'b0;
reg v$FF4_5562_out0 = 1'b0;
reg v$FF4_5563_out0 = 1'b0;
reg v$FF4_5735_out0 = 1'b0;
reg v$FF4_5736_out0 = 1'b0;
reg v$FF4_9118_out0 = 1'b0;
reg v$FF5_11452_out0 = 1'b0;
reg v$FF5_11453_out0 = 1'b0;
reg v$FF5_11521_out0 = 1'b0;
reg v$FF5_13141_out0 = 1'b0;
reg v$FF5_13142_out0 = 1'b0;
reg v$FF5_3159_out0 = 1'b0;
reg v$FF5_3160_out0 = 1'b0;
reg v$FF5_933_out0 = 1'b0;
reg v$FF5_934_out0 = 1'b0;
reg v$FF5_935_out0 = 1'b0;
reg v$FF5_936_out0 = 1'b0;
reg v$FF5_937_out0 = 1'b0;
reg v$FF5_938_out0 = 1'b0;
reg v$FF5_939_out0 = 1'b0;
reg v$FF5_940_out0 = 1'b0;
reg v$FF5_941_out0 = 1'b0;
reg v$FF5_942_out0 = 1'b0;
reg v$FF5_943_out0 = 1'b0;
reg v$FF5_944_out0 = 1'b0;
reg v$FF6_10631_out0 = 1'b0;
reg v$FF6_10632_out0 = 1'b0;
reg v$FF6_11336_out0 = 1'b0;
reg v$FF6_1523_out0 = 1'b0;
reg v$FF6_1524_out0 = 1'b0;
reg v$FF6_1525_out0 = 1'b0;
reg v$FF6_1526_out0 = 1'b0;
reg v$FF6_1527_out0 = 1'b0;
reg v$FF6_1528_out0 = 1'b0;
reg v$FF6_1529_out0 = 1'b0;
reg v$FF6_1530_out0 = 1'b0;
reg v$FF6_1531_out0 = 1'b0;
reg v$FF6_1532_out0 = 1'b0;
reg v$FF6_1533_out0 = 1'b0;
reg v$FF6_1534_out0 = 1'b0;
reg v$FF6_6215_out0 = 1'b0;
reg v$FF6_6216_out0 = 1'b0;
reg v$FF7_12855_out0 = 1'b0;
reg v$FF7_12856_out0 = 1'b0;
reg v$FF7_5594_out0 = 1'b0;
reg v$FF7_5595_out0 = 1'b0;
reg v$FF7_5772_out0 = 1'b0;
reg v$FF7_5773_out0 = 1'b0;
reg v$FF7_5774_out0 = 1'b0;
reg v$FF7_5775_out0 = 1'b0;
reg v$FF7_5776_out0 = 1'b0;
reg v$FF7_5777_out0 = 1'b0;
reg v$FF7_5778_out0 = 1'b0;
reg v$FF7_5779_out0 = 1'b0;
reg v$FF7_5780_out0 = 1'b0;
reg v$FF7_5781_out0 = 1'b0;
reg v$FF7_5782_out0 = 1'b0;
reg v$FF7_5783_out0 = 1'b0;
reg v$FF7_8410_out0 = 1'b0;
reg v$FF7_8411_out0 = 1'b0;
reg v$FF7_9941_out0 = 1'b0;
reg v$FF7_9942_out0 = 1'b0;
reg v$FF8_11778_out0 = 1'b0;
reg v$FF8_11779_out0 = 1'b0;
reg v$FF8_5529_out0 = 1'b0;
reg v$FF8_5530_out0 = 1'b0;
reg v$FF8_6889_out0 = 1'b0;
reg v$FF8_6890_out0 = 1'b0;
reg v$FF8_9843_out0 = 1'b0;
reg v$FF8_9844_out0 = 1'b0;
reg v$FF8_9845_out0 = 1'b0;
reg v$FF8_9846_out0 = 1'b0;
reg v$FF8_9847_out0 = 1'b0;
reg v$FF8_9848_out0 = 1'b0;
reg v$FF8_9849_out0 = 1'b0;
reg v$FF8_9850_out0 = 1'b0;
reg v$FF8_9851_out0 = 1'b0;
reg v$FF8_9852_out0 = 1'b0;
reg v$FF8_9853_out0 = 1'b0;
reg v$FF8_9854_out0 = 1'b0;
reg v$FF9_11201_out0 = 1'b0;
reg v$FF9_11202_out0 = 1'b0;
reg v$FF9_6996_out0 = 1'b0;
reg v$FF9_6997_out0 = 1'b0;
reg v$LSB$FF_13171_out0 = 1'b0;
reg v$LSB$FF_13172_out0 = 1'b0;
reg v$REG13_248_out0 = 1'b0;
reg v$REG14_3705_out0 = 1'b0;
reg v$REG1_4808_out0 = 1'b0;
reg v$REG1_6069_out0 = 1'b0;
reg v$REG2_13074_out0 = 1'b0;
reg v$REG2_13075_out0 = 1'b0;
reg v$REG2_3503_out0 = 1'b0;
reg v$REG2_7598_out0 = 1'b0;
reg v$REG2_7599_out0 = 1'b0;
reg v$REG3_12548_out0 = 1'b0;
reg v$REG3_12549_out0 = 1'b0;
reg v$REG4_7248_out0 = 1'b0;
reg v$REG7_4199_out0 = 1'b0;
reg v$REG8_2804_out0 = 1'b0;
reg v$S$FF_7118_out0 = 1'b0;
reg v$S$FF_7119_out0 = 1'b0;
wire  [10:0] v$C1_11027_out0;
wire  [10:0] v$C1_11028_out0;
wire  [10:0] v$SEL5_11341_out0;
wire  [10:0] v$SEL5_11342_out0;
wire  [10:0] v$SEL6_6954_out0;
wire  [10:0] v$SEL6_6955_out0;
wire  [11:0] v$A1_10168_out0;
wire  [11:0] v$A1_10169_out0;
wire  [11:0] v$ADDRESS_10499_out0;
wire  [11:0] v$ADDRESS_10500_out0;
wire  [11:0] v$ADDRESS_11116_out0;
wire  [11:0] v$ADDRESS_11117_out0;
wire  [11:0] v$ADDRESS_3831_out0;
wire  [11:0] v$ADDRESS_3832_out0;
wire  [11:0] v$ADD_1721_out0;
wire  [11:0] v$ADD_1722_out0;
wire  [11:0] v$A_1452_out0;
wire  [11:0] v$A_1453_out0;
wire  [11:0] v$A_1454_out0;
wire  [11:0] v$A_1455_out0;
wire  [11:0] v$B_7905_out0;
wire  [11:0] v$B_7906_out0;
wire  [11:0] v$B_7907_out0;
wire  [11:0] v$B_7908_out0;
wire  [11:0] v$C1_11144_out0;
wire  [11:0] v$C1_11145_out0;
wire  [11:0] v$C4_11121_out0;
wire  [11:0] v$C4_11122_out0;
wire  [11:0] v$END_11670_out0;
wire  [11:0] v$END_11671_out0;
wire  [11:0] v$MUX1_1023_out0;
wire  [11:0] v$MUX2_2435_out0;
wire  [11:0] v$MUX2_2436_out0;
wire  [11:0] v$MUX3_6357_out0;
wire  [11:0] v$MUX4_781_out0;
wire  [11:0] v$MUX4_782_out0;
wire  [11:0] v$MUX5_12042_out0;
wire  [11:0] v$MUX5_12043_out0;
wire  [11:0] v$MUX6_4683_out0;
wire  [11:0] v$MUX6_9803_out0;
wire  [11:0] v$MUX6_9804_out0;
wire  [11:0] v$MUX7_435_out0;
wire  [11:0] v$MUX7_436_out0;
wire  [11:0] v$MUX8_8058_out0;
wire  [11:0] v$MUX8_8059_out0;
wire  [11:0] v$N$VIEWER_819_out0;
wire  [11:0] v$N$VIEWER_820_out0;
wire  [11:0] v$NEXTINSTRUCTIONADDRESS_13095_out0;
wire  [11:0] v$NEXTINSTRUCTIONADDRESS_13096_out0;
wire  [11:0] v$N_10183_out0;
wire  [11:0] v$N_10184_out0;
wire  [11:0] v$N_12713_out0;
wire  [11:0] v$N_12714_out0;
wire  [11:0] v$N_13005_out0;
wire  [11:0] v$N_13006_out0;
wire  [11:0] v$N_5753_out0;
wire  [11:0] v$N_5754_out0;
wire  [11:0] v$N_7568_out0;
wire  [11:0] v$N_7569_out0;
wire  [11:0] v$N_7740_out0;
wire  [11:0] v$N_7741_out0;
wire  [11:0] v$N_825_out0;
wire  [11:0] v$N_826_out0;
wire  [11:0] v$N_9895_out0;
wire  [11:0] v$N_9896_out0;
wire  [11:0] v$PC$NEXT0_1086_out0;
wire  [11:0] v$PC$NEXT1_2199_out0;
wire  [11:0] v$PCNEXT$VIEWER_11005_out0;
wire  [11:0] v$PCNEXT$VIEWER_11006_out0;
wire  [11:0] v$PCNEXT_4654_out0;
wire  [11:0] v$PCNEXT_4655_out0;
wire  [11:0] v$PC_1881_out0;
wire  [11:0] v$PC_1882_out0;
wire  [11:0] v$RAM$ADDR$VIEWER_11138_out0;
wire  [11:0] v$RAM$ADDR$VIEWER_11139_out0;
wire  [11:0] v$RAM$ADDR0_8161_out0;
wire  [11:0] v$RAM$ADDR1_4451_out0;
wire  [11:0] v$RAM$ADDR_10549_out0;
wire  [11:0] v$RAM$ADDR_10550_out0;
wire  [11:0] v$RAM$ADDR_4425_out0;
wire  [11:0] v$RAM$ADDR_4426_out0;
wire  [11:0] v$RAMADDR0_12041_out0;
wire  [11:0] v$RAMADDR1_8300_out0;
wire  [11:0] v$RAMADDRESS_4749_out0;
wire  [11:0] v$RAMADDRESS_4750_out0;
wire  [11:0] v$RAMADDRESS_8378_out0;
wire  [11:0] v$RAMADDRESS_8379_out0;
wire  [11:0] v$RAMADDRMUX_3221_out0;
wire  [11:0] v$RAMADDRMUX_3222_out0;
wire  [11:0] v$RAMADDRMUX_347_out0;
wire  [11:0] v$RAMADDRMUX_348_out0;
wire  [11:0] v$RAMADDRMUX_9758_out0;
wire  [11:0] v$RAMADDRMUX_9759_out0;
wire  [11:0] v$RAMADDR_13293_out0;
wire  [11:0] v$RAMADDR_6006_out0;
wire  [11:0] v$RAMADDR_9169_out0;
wire  [11:0] v$RAMAddress_1183_out0;
wire  [11:0] v$RAMAddress_1184_out0;
wire  [11:0] v$SEL1_1953_out0;
wire  [11:0] v$SEL1_1954_out0;
wire  [11:0] v$SEL1_7748_out0;
wire  [11:0] v$SEL1_7749_out0;
wire  [11:0] v$SEL2_9281_out0;
wire  [11:0] v$SEL2_9282_out0;
wire  [11:0] v$SEL3_513_out0;
wire  [11:0] v$SEL3_514_out0;
wire  [11:0] v$SEL4_589_out0;
wire  [11:0] v$SEL4_590_out0;
wire  [11:0] v$SEL8_8402_out0;
wire  [11:0] v$SEL8_8403_out0;
wire  [11:0] v$SUM_9219_out0;
wire  [11:0] v$SUM_9220_out0;
wire  [11:0] v$_10004_out0;
wire  [11:0] v$_10008_out0;
wire  [11:0] v$_11477_out0;
wire  [11:0] v$_11478_out0;
wire  [11:0] v$_11796_out0;
wire  [11:0] v$_11800_out0;
wire  [11:0] v$_3211_out0;
wire  [11:0] v$_3215_out0;
wire  [11:0] v$_5263_out0;
wire  [11:0] v$_5264_out0;
wire  [11:0] v$_9417_out0;
wire  [11:0] v$_9418_out0;
wire  [11:0] v$_9978_out0;
wire  [11:0] v$_9982_out0;
wire  [12:0] v$C10_6197_out0;
wire  [12:0] v$C10_6198_out0;
wire  [12:0] v$C4_1379_out0;
wire  [12:0] v$C4_1380_out0;
wire  [12:0] v$C5_6_out0;
wire  [12:0] v$C5_7_out0;
wire  [12:0] v$C6_757_out0;
wire  [12:0] v$C6_758_out0;
wire  [12:0] v$C7_4039_out0;
wire  [12:0] v$C7_4040_out0;
wire  [12:0] v$C8_5698_out0;
wire  [12:0] v$C8_5699_out0;
wire  [13:0] v$_10003_out0;
wire  [13:0] v$_10007_out0;
wire  [13:0] v$_11795_out0;
wire  [13:0] v$_11799_out0;
wire  [13:0] v$_3210_out0;
wire  [13:0] v$_3214_out0;
wire  [13:0] v$_9977_out0;
wire  [13:0] v$_9981_out0;
wire  [14:0] v$C2_12781_out0;
wire  [14:0] v$C2_12782_out0;
wire  [14:0] v$C4_5739_out0;
wire  [14:0] v$C4_5741_out0;
wire  [14:0] v$MUX2_9187_out0;
wire  [14:0] v$MUX2_9189_out0;
wire  [14:0] v$SEL2_4179_out0;
wire  [14:0] v$SEL2_4180_out0;
wire  [14:0] v$_10002_out0;
wire  [14:0] v$_10006_out0;
wire  [14:0] v$_10451_out0;
wire  [14:0] v$_10452_out0;
wire  [14:0] v$_11064_out0;
wire  [14:0] v$_11066_out0;
wire  [14:0] v$_11794_out0;
wire  [14:0] v$_11798_out0;
wire  [14:0] v$_3209_out0;
wire  [14:0] v$_3213_out0;
wire  [14:0] v$_7424_out0;
wire  [14:0] v$_7425_out0;
wire  [14:0] v$_9976_out0;
wire  [14:0] v$_9980_out0;
wire  [15:0] v$A$COMPARATOR$IN_699_out0;
wire  [15:0] v$A$COMPARATOR$IN_700_out0;
wire  [15:0] v$A$IN$MULTIPLIER_2784_out0;
wire  [15:0] v$A$IN$MULTIPLIER_2785_out0;
wire  [15:0] v$A$SAVED_10000_out0;
wire  [15:0] v$A$SAVED_10001_out0;
wire  [15:0] v$A$SAVED_11604_out0;
wire  [15:0] v$A$SAVED_11605_out0;
wire  [15:0] v$A$SAVED_2413_out0;
wire  [15:0] v$A$SAVED_2414_out0;
wire  [15:0] v$A$SAVED_6682_out0;
wire  [15:0] v$A$SAVED_6683_out0;
wire  [15:0] v$A$VIEW_11438_out0;
wire  [15:0] v$A$VIEW_11439_out0;
wire  [15:0] v$A1_4421_out0;
wire  [15:0] v$A1_4422_out0;
wire  [15:0] v$A1_6425_out0;
wire  [15:0] v$A1_6426_out0;
wire  [15:0] v$A1_9247_out0;
wire  [15:0] v$A1_9248_out0;
wire  [15:0] v$ADDEROUT_2206_out0;
wire  [15:0] v$ADDEROUT_2207_out0;
wire  [15:0] v$ALUOUT$LOADSTORE_13269_out0;
wire  [15:0] v$ALUOUT$LOADSTORE_13270_out0;
wire  [15:0] v$ALUOUT_11622_out0;
wire  [15:0] v$ALUOUT_11623_out0;
wire  [15:0] v$ALUOUT_12827_out0;
wire  [15:0] v$ALUOUT_12828_out0;
wire  [15:0] v$ALUOUT_3788_out0;
wire  [15:0] v$ALUOUT_3789_out0;
wire  [15:0] v$ALUOUT_4692_out0;
wire  [15:0] v$ALUOUT_4693_out0;
wire  [15:0] v$ALUOUT_6795_out0;
wire  [15:0] v$ALUOUT_6796_out0;
wire  [15:0] v$ANDOUT_4975_out0;
wire  [15:0] v$ANDOUT_4976_out0;
wire  [15:0] v$A_11271_out0;
wire  [15:0] v$A_11272_out0;
wire  [15:0] v$A_11516_out0;
wire  [15:0] v$A_11517_out0;
wire  [15:0] v$A_12094_out0;
wire  [15:0] v$A_12095_out0;
wire  [15:0] v$A_13003_out0;
wire  [15:0] v$A_13004_out0;
wire  [15:0] v$A_1456_out0;
wire  [15:0] v$A_1457_out0;
wire  [15:0] v$A_1951_out0;
wire  [15:0] v$A_1952_out0;
wire  [15:0] v$A_2886_out0;
wire  [15:0] v$A_2887_out0;
wire  [15:0] v$A_5932_out0;
wire  [15:0] v$A_5933_out0;
wire  [15:0] v$A_6399_out0;
wire  [15:0] v$A_6400_out0;
wire  [15:0] v$A_7280_out0;
wire  [15:0] v$A_7281_out0;
wire  [15:0] v$A_9334_out0;
wire  [15:0] v$A_9336_out0;
wire  [15:0] v$A_9338_out0;
wire  [15:0] v$A_9340_out0;
wire  [15:0] v$B$COMPARATOR$IN_12733_out0;
wire  [15:0] v$B$COMPARATOR$IN_12734_out0;
wire  [15:0] v$B$IN$MULTIPLIER_10764_out0;
wire  [15:0] v$B$IN$MULTIPLIER_10765_out0;
wire  [15:0] v$B$IN_7490_out0;
wire  [15:0] v$B$IN_7491_out0;
wire  [15:0] v$B$MERGE_11664_out0;
wire  [15:0] v$B$MERGE_11665_out0;
wire  [15:0] v$B$SAVED_12540_out0;
wire  [15:0] v$B$SAVED_12541_out0;
wire  [15:0] v$B$SAVED_2592_out0;
wire  [15:0] v$B$SAVED_2593_out0;
wire  [15:0] v$B$SAVED_3014_out0;
wire  [15:0] v$B$SAVED_3015_out0;
wire  [15:0] v$B$SAVED_3161_out0;
wire  [15:0] v$B$SAVED_3162_out0;
wire  [15:0] v$B_12100_out0;
wire  [15:0] v$B_12101_out0;
wire  [15:0] v$B_12546_out0;
wire  [15:0] v$B_12547_out0;
wire  [15:0] v$B_12739_out0;
wire  [15:0] v$B_12740_out0;
wire  [15:0] v$B_12845_out0;
wire  [15:0] v$B_12846_out0;
wire  [15:0] v$B_2056_out0;
wire  [15:0] v$B_2057_out0;
wire  [15:0] v$B_3230_out0;
wire  [15:0] v$B_3232_out0;
wire  [15:0] v$B_3234_out0;
wire  [15:0] v$B_3236_out0;
wire  [15:0] v$B_6722_out0;
wire  [15:0] v$B_6723_out0;
wire  [15:0] v$B_7540_out0;
wire  [15:0] v$B_7541_out0;
wire  [15:0] v$B_7913_out0;
wire  [15:0] v$B_7914_out0;
wire  [15:0] v$B_9458_out0;
wire  [15:0] v$B_9459_out0;
wire  [15:0] v$C10_4403_out0;
wire  [15:0] v$C10_4404_out0;
wire  [15:0] v$C1_11442_out0;
wire  [15:0] v$C1_11443_out0;
wire  [15:0] v$C1_12939_out0;
wire  [15:0] v$C1_12940_out0;
wire  [15:0] v$C1_3963_out0;
wire  [15:0] v$C1_3971_out0;
wire  [15:0] v$C1_3977_out0;
wire  [15:0] v$C1_3980_out0;
wire  [15:0] v$C1_3985_out0;
wire  [15:0] v$C1_3990_out0;
wire  [15:0] v$C1_3995_out0;
wire  [15:0] v$C1_4003_out0;
wire  [15:0] v$C1_4009_out0;
wire  [15:0] v$C1_4012_out0;
wire  [15:0] v$C1_4017_out0;
wire  [15:0] v$C1_4022_out0;
wire  [15:0] v$C2_104_out0;
wire  [15:0] v$C2_110_out0;
wire  [15:0] v$C2_113_out0;
wire  [15:0] v$C2_118_out0;
wire  [15:0] v$C2_123_out0;
wire  [15:0] v$C2_128_out0;
wire  [15:0] v$C2_136_out0;
wire  [15:0] v$C2_142_out0;
wire  [15:0] v$C2_145_out0;
wire  [15:0] v$C2_150_out0;
wire  [15:0] v$C2_155_out0;
wire  [15:0] v$C2_6724_out0;
wire  [15:0] v$C2_6725_out0;
wire  [15:0] v$C2_7980_out0;
wire  [15:0] v$C2_7981_out0;
wire  [15:0] v$C2_96_out0;
wire  [15:0] v$C3_7978_out0;
wire  [15:0] v$C3_7979_out0;
wire  [15:0] v$C7_893_out0;
wire  [15:0] v$C7_894_out0;
wire  [15:0] v$C9_13387_out0;
wire  [15:0] v$C9_13388_out0;
wire  [15:0] v$C9_1999_out0;
wire  [15:0] v$C9_2000_out0;
wire  [15:0] v$COUNTERTHRESHOLD_12725_out0;
wire  [15:0] v$COUNTERTHRESHOLD_12726_out0;
wire  [15:0] v$COUNTERVALUE_1747_out0;
wire  [15:0] v$COUNTERVALUE_1748_out0;
wire  [15:0] v$C_12847_out0;
wire  [15:0] v$C_12848_out0;
wire  [15:0] v$DATA$IN0_6953_out0;
wire  [15:0] v$DATA$IN1_10600_out0;
wire  [15:0] v$DATA$IN_4809_out0;
wire  [15:0] v$DATA$IN_4810_out0;
wire  [15:0] v$DATA$IN_811_out0;
wire  [15:0] v$DATA$IN_812_out0;
wire  [15:0] v$DATA$OUT0_8072_out0;
wire  [15:0] v$DATA$OUT1_10871_out0;
wire  [15:0] v$DATA$OUT_5146_out0;
wire  [15:0] v$DATA$OUT_5147_out0;
wire  [15:0] v$DATA$OUT_538_out0;
wire  [15:0] v$DATA$OUT_539_out0;
wire  [15:0] v$DATAIN0_7296_out0;
wire  [15:0] v$DATAIN1_6590_out0;
wire  [15:0] v$DATAINCP_7244_out0;
wire  [15:0] v$DATAINCP_7245_out0;
wire  [15:0] v$DATA_3010_out0;
wire  [15:0] v$DATA_3011_out0;
wire  [15:0] v$DATA_9478_out0;
wire  [15:0] v$DATA_9479_out0;
wire  [15:0] v$DIN$FIRST$MUX_5070_out0;
wire  [15:0] v$DIN$FIRST$MUX_5071_out0;
wire  [15:0] v$DIN3$VIEWER_1146_out0;
wire  [15:0] v$DIN3$VIEWER_1147_out0;
wire  [15:0] v$DIN3_9801_out0;
wire  [15:0] v$DIN3_9802_out0;
wire  [15:0] v$DIN_903_out0;
wire  [15:0] v$DIN_904_out0;
wire  [15:0] v$DIN_977_out0;
wire  [15:0] v$DIN_978_out0;
wire  [15:0] v$DM1_5380_out0;
wire  [15:0] v$DM1_5380_out1;
wire  [15:0] v$DOUT1_1887_out0;
wire  [15:0] v$DOUT1_1888_out0;
wire  [15:0] v$DOUT2_2214_out0;
wire  [15:0] v$DOUT2_2215_out0;
wire  [15:0] v$FPU$A_11096_out0;
wire  [15:0] v$FPU$A_11097_out0;
wire  [15:0] v$FPU$B_4772_out0;
wire  [15:0] v$FPU$B_4773_out0;
wire  [15:0] v$FPU$OUT_12069_out0;
wire  [15:0] v$FPU$OUT_12070_out0;
wire  [15:0] v$HAZ$DECTECTOR$A_12727_out0;
wire  [15:0] v$HAZ$DECTECTOR$A_12728_out0;
wire  [15:0] v$HAZ$DETECTOR$B_3447_out0;
wire  [15:0] v$HAZ$DETECTOR$B_3448_out0;
wire  [15:0] v$INSTR$READ0_9560_out0;
wire  [15:0] v$INSTR$READ1_7747_out0;
wire  [15:0] v$INSTR$READ_10224_out0;
wire  [15:0] v$INSTR$READ_10225_out0;
wire  [15:0] v$INSTR$READ_4830_out0;
wire  [15:0] v$INSTR$READ_4831_out0;
wire  [15:0] v$IN_180_out0;
wire  [15:0] v$IN_181_out0;
wire  [15:0] v$IN_3016_out0;
wire  [15:0] v$IN_3017_out0;
wire  [15:0] v$IN_3018_out0;
wire  [15:0] v$IN_3019_out0;
wire  [15:0] v$IN_3020_out0;
wire  [15:0] v$IN_3021_out0;
wire  [15:0] v$IN_3022_out0;
wire  [15:0] v$IN_3023_out0;
wire  [15:0] v$IN_6532_out0;
wire  [15:0] v$IN_6533_out0;
wire  [15:0] v$IN_6534_out0;
wire  [15:0] v$IN_6535_out0;
wire  [15:0] v$IN_6536_out0;
wire  [15:0] v$IN_6537_out0;
wire  [15:0] v$IN_6538_out0;
wire  [15:0] v$IN_6539_out0;
wire  [15:0] v$IN_9132_out0;
wire  [15:0] v$IN_9133_out0;
wire  [15:0] v$IN_9134_out0;
wire  [15:0] v$IN_9136_out0;
wire  [15:0] v$IN_9137_out0;
wire  [15:0] v$IN_9138_out0;
wire  [15:0] v$IN_9140_out0;
wire  [15:0] v$IN_9141_out0;
wire  [15:0] v$IN_9142_out0;
wire  [15:0] v$IN_9144_out0;
wire  [15:0] v$IN_9145_out0;
wire  [15:0] v$IN_9146_out0;
wire  [15:0] v$IR$READ$IN$PREV$CYCLE_4206_out0;
wire  [15:0] v$IR$READ$IN$PREV$CYCLE_4207_out0;
wire  [15:0] v$IR1$VIEWER_5010_out0;
wire  [15:0] v$IR1$VIEWER_5011_out0;
wire  [15:0] v$IR1_11186_out0;
wire  [15:0] v$IR1_11187_out0;
wire  [15:0] v$IR1_11742_out0;
wire  [15:0] v$IR1_11743_out0;
wire  [15:0] v$IR1_12803_out0;
wire  [15:0] v$IR1_12804_out0;
wire  [15:0] v$IR1_24_out0;
wire  [15:0] v$IR1_25_out0;
wire  [15:0] v$IR1_2845_out0;
wire  [15:0] v$IR1_2846_out0;
wire  [15:0] v$IR1_370_out0;
wire  [15:0] v$IR1_371_out0;
wire  [15:0] v$IR1_5151_out0;
wire  [15:0] v$IR1_5152_out0;
wire  [15:0] v$IR1_8963_out0;
wire  [15:0] v$IR1_8964_out0;
wire  [15:0] v$IR2$VIEWER_11430_out0;
wire  [15:0] v$IR2$VIEWER_11431_out0;
wire  [15:0] v$IR2_1150_out0;
wire  [15:0] v$IR2_1151_out0;
wire  [15:0] v$IR2_11640_out0;
wire  [15:0] v$IR2_11641_out0;
wire  [15:0] v$IR2_12729_out0;
wire  [15:0] v$IR2_12730_out0;
wire  [15:0] v$IR2_1700_out0;
wire  [15:0] v$IR2_1701_out0;
wire  [15:0] v$IR2_1985_out0;
wire  [15:0] v$IR2_1986_out0;
wire  [15:0] v$IR2_2660_out0;
wire  [15:0] v$IR2_2661_out0;
wire  [15:0] v$IR2_5306_out0;
wire  [15:0] v$IR2_5307_out0;
wire  [15:0] v$IR2_929_out0;
wire  [15:0] v$IR2_930_out0;
wire  [15:0] v$LDST$RAMDOUT_453_out0;
wire  [15:0] v$LDST$RAMDOUT_454_out0;
wire  [15:0] v$LDST$RMN_5273_out0;
wire  [15:0] v$LDST$RMN_5274_out0;
wire  [15:0] v$LDSTN_1793_out0;
wire  [15:0] v$LDSTN_1794_out0;
wire  [15:0] v$LDSTRM_5177_out0;
wire  [15:0] v$LDSTRM_5178_out0;
wire  [15:0] v$LOAD$STORE$OUT_12382_out0;
wire  [15:0] v$LOAD$STORE$OUT_12383_out0;
wire  [15:0] v$LOWER$PART_5054_out0;
wire  [15:0] v$LOWER$PART_5055_out0;
wire  [15:0] v$MULTIPLY$DENORMALIZATION$16$BIT_7536_out0;
wire  [15:0] v$MULTIPLY$DENORMALIZATION$16$BIT_7537_out0;
wire  [15:0] v$MUX10_11878_out0;
wire  [15:0] v$MUX10_11879_out0;
wire  [15:0] v$MUX11_5920_out0;
wire  [15:0] v$MUX11_5921_out0;
wire  [15:0] v$MUX13_1458_out0;
wire  [15:0] v$MUX13_1459_out0;
wire  [15:0] v$MUX15_4768_out0;
wire  [15:0] v$MUX15_4769_out0;
wire  [15:0] v$MUX16_13179_out0;
wire  [15:0] v$MUX16_13180_out0;
wire  [15:0] v$MUX1_10579_out0;
wire  [15:0] v$MUX1_10580_out0;
wire  [15:0] v$MUX1_1139_out0;
wire  [15:0] v$MUX1_1140_out0;
wire  [15:0] v$MUX1_12538_out0;
wire  [15:0] v$MUX1_12539_out0;
wire  [15:0] v$MUX1_13028_out0;
wire  [15:0] v$MUX1_13029_out0;
wire  [15:0] v$MUX1_1505_out0;
wire  [15:0] v$MUX1_1506_out0;
wire  [15:0] v$MUX1_2758_out0;
wire  [15:0] v$MUX1_2759_out0;
wire  [15:0] v$MUX1_3839_out0;
wire  [15:0] v$MUX1_3840_out0;
wire  [15:0] v$MUX1_4667_out0;
wire  [15:0] v$MUX1_4668_out0;
wire  [15:0] v$MUX1_4669_out0;
wire  [15:0] v$MUX1_4670_out0;
wire  [15:0] v$MUX1_4671_out0;
wire  [15:0] v$MUX1_4672_out0;
wire  [15:0] v$MUX1_4673_out0;
wire  [15:0] v$MUX1_4674_out0;
wire  [15:0] v$MUX1_7566_out0;
wire  [15:0] v$MUX1_7567_out0;
wire  [15:0] v$MUX1_985_out0;
wire  [15:0] v$MUX1_986_out0;
wire  [15:0] v$MUX2_10495_out0;
wire  [15:0] v$MUX2_10496_out0;
wire  [15:0] v$MUX2_11061_out0;
wire  [15:0] v$MUX2_7000_out0;
wire  [15:0] v$MUX2_7001_out0;
wire  [15:0] v$MUX2_7752_out0;
wire  [15:0] v$MUX2_7753_out0;
wire  [15:0] v$MUX2_7822_out0;
wire  [15:0] v$MUX2_7823_out0;
wire  [15:0] v$MUX2_7824_out0;
wire  [15:0] v$MUX2_7825_out0;
wire  [15:0] v$MUX2_7826_out0;
wire  [15:0] v$MUX2_7827_out0;
wire  [15:0] v$MUX2_7828_out0;
wire  [15:0] v$MUX2_7829_out0;
wire  [15:0] v$MUX3_1098_out0;
wire  [15:0] v$MUX3_1099_out0;
wire  [15:0] v$MUX3_1100_out0;
wire  [15:0] v$MUX3_1101_out0;
wire  [15:0] v$MUX3_1102_out0;
wire  [15:0] v$MUX3_1103_out0;
wire  [15:0] v$MUX3_1104_out0;
wire  [15:0] v$MUX3_1105_out0;
wire  [15:0] v$MUX3_13078_out0;
wire  [15:0] v$MUX3_13079_out0;
wire  [15:0] v$MUX3_2588_out0;
wire  [15:0] v$MUX3_2589_out0;
wire  [15:0] v$MUX3_787_out0;
wire  [15:0] v$MUX3_788_out0;
wire  [15:0] v$MUX4_11178_out0;
wire  [15:0] v$MUX4_11179_out0;
wire  [15:0] v$MUX4_11180_out0;
wire  [15:0] v$MUX4_11181_out0;
wire  [15:0] v$MUX4_11182_out0;
wire  [15:0] v$MUX4_11183_out0;
wire  [15:0] v$MUX4_11184_out0;
wire  [15:0] v$MUX4_11185_out0;
wire  [15:0] v$MUX4_12532_out0;
wire  [15:0] v$MUX4_12533_out0;
wire  [15:0] v$MUX4_2551_out0;
wire  [15:0] v$MUX4_3947_out0;
wire  [15:0] v$MUX4_3948_out0;
wire  [15:0] v$MUX4_42_out0;
wire  [15:0] v$MUX4_43_out0;
wire  [15:0] v$MUX4_849_out0;
wire  [15:0] v$MUX4_850_out0;
wire  [15:0] v$MUX5_7180_out0;
wire  [15:0] v$MUX5_7734_out0;
wire  [15:0] v$MUX5_7735_out0;
wire  [15:0] v$MUX5_9474_out0;
wire  [15:0] v$MUX5_9475_out0;
wire  [15:0] v$MUX6_3439_out0;
wire  [15:0] v$MUX6_3440_out0;
wire  [15:0] v$MUX6_5016_out0;
wire  [15:0] v$MUX6_5017_out0;
wire  [15:0] v$MUX9_12717_out0;
wire  [15:0] v$MUX9_12718_out0;
wire  [15:0] v$NEXTENDED_1060_out0;
wire  [15:0] v$NEXTENDED_1061_out0;
wire  [15:0] v$NEXTENDED_9754_out0;
wire  [15:0] v$NEXTENDED_9755_out0;
wire  [15:0] v$OP1_10521_out0;
wire  [15:0] v$OP1_10522_out0;
wire  [15:0] v$OP1_3661_out0;
wire  [15:0] v$OP1_3662_out0;
wire  [15:0] v$OP2_10356_out0;
wire  [15:0] v$OP2_10357_out0;
wire  [15:0] v$OP2_5118_out0;
wire  [15:0] v$OP2_5119_out0;
wire  [15:0] v$OP2_6767_out0;
wire  [15:0] v$OP2_6768_out0;
wire  [15:0] v$OP2_9394_out0;
wire  [15:0] v$OP2_9395_out0;
wire  [15:0] v$OUT_1899_out0;
wire  [15:0] v$OUT_1900_out0;
wire  [15:0] v$OUT_1901_out0;
wire  [15:0] v$OUT_1902_out0;
wire  [15:0] v$OUT_1903_out0;
wire  [15:0] v$OUT_1904_out0;
wire  [15:0] v$OUT_1905_out0;
wire  [15:0] v$OUT_1906_out0;
wire  [15:0] v$OUT_3625_out0;
wire  [15:0] v$OUT_3626_out0;
wire  [15:0] v$OUT_551_out0;
wire  [15:0] v$OUT_552_out0;
wire  [15:0] v$OUT_8119_out0;
wire  [15:0] v$OUT_8121_out0;
wire  [15:0] v$OUT_9893_out0;
wire  [15:0] v$OUT_9894_out0;
wire  [15:0] v$PIN_1702_out0;
wire  [15:0] v$PIN_1703_out0;
wire  [15:0] v$R0TEST_5724_out0;
wire  [15:0] v$R0TEST_5725_out0;
wire  [15:0] v$R0TEST_9432_out0;
wire  [15:0] v$R0TEST_9433_out0;
wire  [15:0] v$R0_1977_out0;
wire  [15:0] v$R0_1978_out0;
wire  [15:0] v$R1TEST_10449_out0;
wire  [15:0] v$R1TEST_10450_out0;
wire  [15:0] v$R1TEST_5732_out0;
wire  [15:0] v$R1TEST_5733_out0;
wire  [15:0] v$R1_9296_out0;
wire  [15:0] v$R1_9297_out0;
wire  [15:0] v$R2TEST_10971_out0;
wire  [15:0] v$R2TEST_10972_out0;
wire  [15:0] v$R2TEST_11029_out0;
wire  [15:0] v$R2TEST_11030_out0;
wire  [15:0] v$R2_5454_out0;
wire  [15:0] v$R2_5455_out0;
wire  [15:0] v$R3TEST_5094_out0;
wire  [15:0] v$R3TEST_5095_out0;
wire  [15:0] v$R3TEST_7604_out0;
wire  [15:0] v$R3TEST_7605_out0;
wire  [15:0] v$R3_7072_out0;
wire  [15:0] v$R3_7073_out0;
wire  [15:0] v$RAM1_8558_out0;
wire  [15:0] v$RAMDIN_4792_out0;
wire  [15:0] v$RAMDIN_4793_out0;
wire  [15:0] v$RAMDOUT$DATAPATH_366_out0;
wire  [15:0] v$RAMDOUT$DATAPATH_367_out0;
wire  [15:0] v$RAMDOUT0_6338_out0;
wire  [15:0] v$RAMDOUT1_5788_out0;
wire  [15:0] v$RAMDOUT_11827_out0;
wire  [15:0] v$RAMDOUT_11828_out0;
wire  [15:0] v$RAMDOUT_3669_out0;
wire  [15:0] v$RAMDOUT_3670_out0;
wire  [15:0] v$RAMDOUT_5424_out0;
wire  [15:0] v$RAMDOUT_5425_out0;
wire  [15:0] v$RAMDOUT_66_out0;
wire  [15:0] v$RAMDOUT_67_out0;
wire  [15:0] v$RAMDOutOut_1911_out0;
wire  [15:0] v$RAMDOutOut_1912_out0;
wire  [15:0] v$RDOUT_6895_out0;
wire  [15:0] v$RDOUT_6896_out0;
wire  [15:0] v$RD_1154_out0;
wire  [15:0] v$RD_1155_out0;
wire  [15:0] v$REGDIN_11576_out0;
wire  [15:0] v$REGDIN_11577_out0;
wire  [15:0] v$REGDIN_13076_out0;
wire  [15:0] v$REGDIN_13077_out0;
wire  [15:0] v$RMN_4169_out0;
wire  [15:0] v$RMN_4170_out0;
wire  [15:0] v$RMORIGINAL_8617_out0;
wire  [15:0] v$RMORIGINAL_8618_out0;
wire  [15:0] v$RM_11349_out0;
wire  [15:0] v$RM_11350_out0;
wire  [15:0] v$RM_12933_out0;
wire  [15:0] v$RM_12934_out0;
wire  [15:0] v$RM_13239_out0;
wire  [15:0] v$RM_13240_out0;
wire  [15:0] v$RM_6421_out0;
wire  [15:0] v$RM_6422_out0;
wire  [15:0] v$RM_6813_out0;
wire  [15:0] v$RM_6814_out0;
wire  [15:0] v$ROM1_12254_out0;
wire  [15:0] v$ROM1_12255_out0;
wire  [15:0] v$R_13054_out0;
wire  [15:0] v$R_13055_out0;
wire  [15:0] v$R_56_out0;
wire  [15:0] v$R_57_out0;
wire  [15:0] v$SEL1_10679_out0;
wire  [15:0] v$SEL1_10683_out0;
wire  [15:0] v$SEL1_10689_out0;
wire  [15:0] v$SEL1_10696_out0;
wire  [15:0] v$SEL1_10701_out0;
wire  [15:0] v$SEL1_10706_out0;
wire  [15:0] v$SEL1_10711_out0;
wire  [15:0] v$SEL1_10715_out0;
wire  [15:0] v$SEL1_10721_out0;
wire  [15:0] v$SEL1_10728_out0;
wire  [15:0] v$SEL1_10733_out0;
wire  [15:0] v$SEL1_10738_out0;
wire  [15:0] v$SEL1_11746_out0;
wire  [15:0] v$SEL1_11750_out0;
wire  [15:0] v$SEL1_11754_out0;
wire  [15:0] v$SEL1_11758_out0;
wire  [15:0] v$SEL1_5935_out0;
wire  [15:0] v$SEL1_5939_out0;
wire  [15:0] v$SEL1_5945_out0;
wire  [15:0] v$SEL1_5952_out0;
wire  [15:0] v$SEL1_5957_out0;
wire  [15:0] v$SEL1_5962_out0;
wire  [15:0] v$SEL1_5967_out0;
wire  [15:0] v$SEL1_5971_out0;
wire  [15:0] v$SEL1_5977_out0;
wire  [15:0] v$SEL1_5984_out0;
wire  [15:0] v$SEL1_5989_out0;
wire  [15:0] v$SEL1_5994_out0;
wire  [15:0] v$SEL2_9368_out0;
wire  [15:0] v$SEL2_9372_out0;
wire  [15:0] v$SEL2_9376_out0;
wire  [15:0] v$SEL2_9380_out0;
wire  [15:0] v$SEL3_4957_out0;
wire  [15:0] v$SEL3_4961_out0;
wire  [15:0] v$SEL3_4965_out0;
wire  [15:0] v$SEL3_4969_out0;
wire  [15:0] v$SEL4_6522_out0;
wire  [15:0] v$SEL4_6523_out0;
wire  [15:0] v$SEL5_9159_out0;
wire  [15:0] v$SEL5_9160_out0;
wire  [15:0] v$SHIFT1OUT_5120_out0;
wire  [15:0] v$SHIFT1OUT_5121_out0;
wire  [15:0] v$SHIFT2OUT_10942_out0;
wire  [15:0] v$SHIFT2OUT_10943_out0;
wire  [15:0] v$SHIFT4OUT_3949_out0;
wire  [15:0] v$SHIFT4OUT_3950_out0;
wire  [15:0] v$SHIFT8OUT_5516_out0;
wire  [15:0] v$SHIFT8OUT_5517_out0;
wire  [15:0] v$SUM_6865_out0;
wire  [15:0] v$SUM_6866_out0;
wire  [15:0] v$THRESHOLD_10815_out0;
wire  [15:0] v$THRESHOLD_10816_out0;
wire  [15:0] v$UART$DOUT_12260_out0;
wire  [15:0] v$UART$DOUT_12261_out0;
wire  [15:0] v$XOR1_3455_out0;
wire  [15:0] v$XOR1_3456_out0;
wire  [15:0] v$XOR1_6518_out0;
wire  [15:0] v$XOR1_6519_out0;
wire  [15:0] v$_11477_out1;
wire  [15:0] v$_11478_out1;
wire  [15:0] v$_11479_out0;
wire  [15:0] v$_11480_out0;
wire  [15:0] v$_12276_out0;
wire  [15:0] v$_12277_out0;
wire  [15:0] v$_13103_out0;
wire  [15:0] v$_13105_out0;
wire  [15:0] v$_4688_out0;
wire  [15:0] v$_4689_out0;
wire  [15:0] v$_6441_out0;
wire  [15:0] v$_6442_out0;
wire  [15:0] v$_6443_out0;
wire  [15:0] v$_6444_out0;
wire  [15:0] v$_6445_out0;
wire  [15:0] v$_6446_out0;
wire  [15:0] v$_6447_out0;
wire  [15:0] v$_6448_out0;
wire  [15:0] v$_6656_out1;
wire  [15:0] v$_6657_out1;
wire  [15:0] v$_709_out0;
wire  [15:0] v$_710_out0;
wire  [15:0] v$_711_out0;
wire  [15:0] v$_712_out0;
wire  [15:0] v$_713_out0;
wire  [15:0] v$_714_out0;
wire  [15:0] v$_715_out0;
wire  [15:0] v$_716_out0;
wire  [15:0] v$_723_out0;
wire  [15:0] v$_724_out0;
wire  [15:0] v$_7486_out0;
wire  [15:0] v$_7487_out0;
wire  [15:0] v$_7572_out0;
wire  [15:0] v$_7573_out0;
wire  [15:0] v$_7608_out0;
wire  [15:0] v$_7609_out0;
wire  [15:0] v$_7610_out0;
wire  [15:0] v$_7611_out0;
wire  [15:0] v$_7612_out0;
wire  [15:0] v$_7613_out0;
wire  [15:0] v$_7614_out0;
wire  [15:0] v$_7615_out0;
wire  [15:0] v$_8000_out0;
wire  [15:0] v$_8001_out0;
wire  [15:0] v$_8877_out0;
wire  [15:0] v$_8878_out0;
wire  [15:0] v$_8879_out0;
wire  [15:0] v$_8880_out0;
wire  [15:0] v$_8881_out0;
wire  [15:0] v$_8882_out0;
wire  [15:0] v$_8883_out0;
wire  [15:0] v$_8884_out0;
wire  [19:0] v$SEL1_10681_out0;
wire  [19:0] v$SEL1_10698_out0;
wire  [19:0] v$SEL1_10703_out0;
wire  [19:0] v$SEL1_10708_out0;
wire  [19:0] v$SEL1_10713_out0;
wire  [19:0] v$SEL1_10730_out0;
wire  [19:0] v$SEL1_10735_out0;
wire  [19:0] v$SEL1_10740_out0;
wire  [19:0] v$SEL1_5937_out0;
wire  [19:0] v$SEL1_5954_out0;
wire  [19:0] v$SEL1_5959_out0;
wire  [19:0] v$SEL1_5964_out0;
wire  [19:0] v$SEL1_5969_out0;
wire  [19:0] v$SEL1_5986_out0;
wire  [19:0] v$SEL1_5991_out0;
wire  [19:0] v$SEL1_5996_out0;
wire  [1:0] v$2_8391_out0;
wire  [1:0] v$2_8392_out0;
wire  [1:0] v$5_5074_out0;
wire  [1:0] v$5_5075_out0;
wire  [1:0] v$7_9409_out0;
wire  [1:0] v$7_9410_out0;
wire  [1:0] v$8_481_out0;
wire  [1:0] v$8_482_out0;
wire  [1:0] v$AD1VIEWER_4770_out0;
wire  [1:0] v$AD1VIEWER_4771_out0;
wire  [1:0] v$AD1_1011_out0;
wire  [1:0] v$AD1_1012_out0;
wire  [1:0] v$AD1_13302_out0;
wire  [1:0] v$AD1_13303_out0;
wire  [1:0] v$AD1_4656_out0;
wire  [1:0] v$AD1_4657_out0;
wire  [1:0] v$AD1_5142_out0;
wire  [1:0] v$AD1_5143_out0;
wire  [1:0] v$AD2$viewer_10993_out0;
wire  [1:0] v$AD2$viewer_10994_out0;
wire  [1:0] v$AD2_10930_out0;
wire  [1:0] v$AD2_10931_out0;
wire  [1:0] v$AD2_2656_out0;
wire  [1:0] v$AD2_2657_out0;
wire  [1:0] v$AD2_4413_out0;
wire  [1:0] v$AD2_4414_out0;
wire  [1:0] v$AD2_6334_out0;
wire  [1:0] v$AD2_6335_out0;
wire  [1:0] v$AD3$VIEWER_5791_out0;
wire  [1:0] v$AD3$VIEWER_5792_out0;
wire  [1:0] v$AD3_10447_out0;
wire  [1:0] v$AD3_10448_out0;
wire  [1:0] v$AD3_8756_out0;
wire  [1:0] v$AD3_8757_out0;
wire  [1:0] v$C1_1779_out0;
wire  [1:0] v$C1_1780_out0;
wire  [1:0] v$C1_3967_out0;
wire  [1:0] v$C1_3970_out0;
wire  [1:0] v$C1_3976_out0;
wire  [1:0] v$C1_3984_out0;
wire  [1:0] v$C1_3989_out0;
wire  [1:0] v$C1_3994_out0;
wire  [1:0] v$C1_3999_out0;
wire  [1:0] v$C1_4002_out0;
wire  [1:0] v$C1_4008_out0;
wire  [1:0] v$C1_4016_out0;
wire  [1:0] v$C1_4021_out0;
wire  [1:0] v$C1_4026_out0;
wire  [1:0] v$C1_5267_out0;
wire  [1:0] v$C1_5268_out0;
wire  [1:0] v$C1_5479_out0;
wire  [1:0] v$C1_5483_out0;
wire  [1:0] v$C1_9650_out0;
wire  [1:0] v$C1_9651_out0;
wire  [1:0] v$C2_100_out0;
wire  [1:0] v$C2_103_out0;
wire  [1:0] v$C2_109_out0;
wire  [1:0] v$C2_117_out0;
wire  [1:0] v$C2_122_out0;
wire  [1:0] v$C2_127_out0;
wire  [1:0] v$C2_132_out0;
wire  [1:0] v$C2_135_out0;
wire  [1:0] v$C2_141_out0;
wire  [1:0] v$C2_149_out0;
wire  [1:0] v$C2_154_out0;
wire  [1:0] v$C2_159_out0;
wire  [1:0] v$C2_8960_out0;
wire  [1:0] v$C2_8961_out0;
wire  [1:0] v$C3_2001_out0;
wire  [1:0] v$C3_2002_out0;
wire  [1:0] v$C3_2003_out0;
wire  [1:0] v$C3_2004_out0;
wire  [1:0] v$C3_2005_out0;
wire  [1:0] v$C3_2006_out0;
wire  [1:0] v$C3_2007_out0;
wire  [1:0] v$C3_2008_out0;
wire  [1:0] v$C3_2009_out0;
wire  [1:0] v$C3_2010_out0;
wire  [1:0] v$C3_2011_out0;
wire  [1:0] v$C3_2012_out0;
wire  [1:0] v$C4_11432_out0;
wire  [1:0] v$C4_11433_out0;
wire  [1:0] v$C4_11588_out0;
wire  [1:0] v$C4_11589_out0;
wire  [1:0] v$C4_11590_out0;
wire  [1:0] v$C4_11591_out0;
wire  [1:0] v$C4_11592_out0;
wire  [1:0] v$C4_11593_out0;
wire  [1:0] v$C4_11594_out0;
wire  [1:0] v$C4_11595_out0;
wire  [1:0] v$C4_11596_out0;
wire  [1:0] v$C4_11597_out0;
wire  [1:0] v$C4_11598_out0;
wire  [1:0] v$C4_11599_out0;
wire  [1:0] v$C4_11600_out0;
wire  [1:0] v$C4_11601_out0;
wire  [1:0] v$C4_11602_out0;
wire  [1:0] v$C4_11603_out0;
wire  [1:0] v$C5_11957_out0;
wire  [1:0] v$C5_11958_out0;
wire  [1:0] v$C5_11959_out0;
wire  [1:0] v$C5_11960_out0;
wire  [1:0] v$C5_11961_out0;
wire  [1:0] v$C5_11962_out0;
wire  [1:0] v$C5_11963_out0;
wire  [1:0] v$C5_11964_out0;
wire  [1:0] v$C5_11965_out0;
wire  [1:0] v$C5_11966_out0;
wire  [1:0] v$C5_11967_out0;
wire  [1:0] v$C5_11968_out0;
wire  [1:0] v$C5_11969_out0;
wire  [1:0] v$C5_11970_out0;
wire  [1:0] v$C5_11971_out0;
wire  [1:0] v$C5_11972_out0;
wire  [1:0] v$C6_4536_out0;
wire  [1:0] v$C6_4537_out0;
wire  [1:0] v$C6_4538_out0;
wire  [1:0] v$C6_4539_out0;
wire  [1:0] v$C6_4540_out0;
wire  [1:0] v$C6_4541_out0;
wire  [1:0] v$C6_4542_out0;
wire  [1:0] v$C6_4543_out0;
wire  [1:0] v$C6_4544_out0;
wire  [1:0] v$C6_4545_out0;
wire  [1:0] v$C6_4546_out0;
wire  [1:0] v$C6_4547_out0;
wire  [1:0] v$C6_4548_out0;
wire  [1:0] v$C6_4549_out0;
wire  [1:0] v$C6_4550_out0;
wire  [1:0] v$C6_4551_out0;
wire  [1:0] v$END_317_out0;
wire  [1:0] v$END_318_out0;
wire  [1:0] v$FPU$OP_10984_out0;
wire  [1:0] v$FPU$OP_10985_out0;
wire  [1:0] v$FPU$OP_8416_out0;
wire  [1:0] v$FPU$OP_8417_out0;
wire  [1:0] v$FPU$OP_9460_out0;
wire  [1:0] v$FPU$OP_9461_out0;
wire  [1:0] v$INTERRUPTNUMBER_36_out0;
wire  [1:0] v$INTERRUPTNUMBER_37_out0;
wire  [1:0] v$IR1$D_10187_out0;
wire  [1:0] v$IR1$D_10188_out0;
wire  [1:0] v$IR1$D_2900_out0;
wire  [1:0] v$IR1$D_2901_out0;
wire  [1:0] v$IR1$FPU$OP$CODE_13016_out0;
wire  [1:0] v$IR1$FPU$OP$CODE_13017_out0;
wire  [1:0] v$IR1$FPU$OP_2545_out0;
wire  [1:0] v$IR1$FPU$OP_2546_out0;
wire  [1:0] v$IR1$M_8274_out0;
wire  [1:0] v$IR1$M_8275_out0;
wire  [1:0] v$IR1$M_8836_out0;
wire  [1:0] v$IR1$M_8837_out0;
wire  [1:0] v$IR1$RD$VIEWER_13072_out0;
wire  [1:0] v$IR1$RD$VIEWER_13073_out0;
wire  [1:0] v$IR1$RD_3732_out0;
wire  [1:0] v$IR1$RD_3733_out0;
wire  [1:0] v$IR1$RM$VIEWER_5422_out0;
wire  [1:0] v$IR1$RM$VIEWER_5423_out0;
wire  [1:0] v$IR1$RM_13011_out0;
wire  [1:0] v$IR1$RM_13012_out0;
wire  [1:0] v$IR1$RM_20_out0;
wire  [1:0] v$IR1$RM_21_out0;
wire  [1:0] v$IR2$D_3290_out0;
wire  [1:0] v$IR2$D_3291_out0;
wire  [1:0] v$IR2$D_9879_out0;
wire  [1:0] v$IR2$D_9880_out0;
wire  [1:0] v$IR2$FPU$OP_1657_out0;
wire  [1:0] v$IR2$FPU$OP_1658_out0;
wire  [1:0] v$IR2$FPU$OP_5098_out0;
wire  [1:0] v$IR2$FPU$OP_5099_out0;
wire  [1:0] v$IR2$FPU$OP_881_out0;
wire  [1:0] v$IR2$FPU$OP_882_out0;
wire  [1:0] v$IR2$M_6072_out0;
wire  [1:0] v$IR2$M_6073_out0;
wire  [1:0] v$IR2$M_8626_out0;
wire  [1:0] v$IR2$M_8627_out0;
wire  [1:0] v$IR2$RD$VIEWER_6358_out0;
wire  [1:0] v$IR2$RD$VIEWER_6359_out0;
wire  [1:0] v$IR2$RD_11468_out0;
wire  [1:0] v$IR2$RD_11469_out0;
wire  [1:0] v$IR2$RD_8874_out0;
wire  [1:0] v$IR2$RD_8875_out0;
wire  [1:0] v$MUX10_2334_out0;
wire  [1:0] v$MUX10_2335_out0;
wire  [1:0] v$MUX11_3121_out0;
wire  [1:0] v$MUX11_3122_out0;
wire  [1:0] v$MUX1_5804_out0;
wire  [1:0] v$MUX1_5805_out0;
wire  [1:0] v$MUX2_1661_out0;
wire  [1:0] v$MUX2_1662_out0;
wire  [1:0] v$MUX5_5450_out0;
wire  [1:0] v$MUX5_5451_out0;
wire  [1:0] v$MUX6_542_out0;
wire  [1:0] v$MUX6_543_out0;
wire  [1:0] v$MUX9_5181_out0;
wire  [1:0] v$MUX9_5182_out0;
wire  [1:0] v$NINTERRUPT_798_out0;
wire  [1:0] v$NINTERRUPT_799_out0;
wire  [1:0] v$NINT_1603_out0;
wire  [1:0] v$NINT_1604_out0;
wire  [1:0] v$OP_553_out0;
wire  [1:0] v$OP_554_out0;
wire  [1:0] v$S$REG_2143_out0;
wire  [1:0] v$S$REG_2144_out0;
wire  [1:0] v$SEL10_8472_out0;
wire  [1:0] v$SEL10_8473_out0;
wire  [1:0] v$SEL13_3246_out0;
wire  [1:0] v$SEL13_3247_out0;
wire  [1:0] v$SEL1_3611_out0;
wire  [1:0] v$SEL1_3612_out0;
wire  [1:0] v$SEL4_6439_out0;
wire  [1:0] v$SEL4_6440_out0;
wire  [1:0] v$SEL5_368_out0;
wire  [1:0] v$SEL5_369_out0;
wire  [1:0] v$SEL6_1769_out0;
wire  [1:0] v$SEL6_1770_out0;
wire  [1:0] v$SEL8_10430_out0;
wire  [1:0] v$SEL8_10431_out0;
wire  [1:0] v$SEL9_5490_out0;
wire  [1:0] v$SEL9_5491_out0;
wire  [1:0] v$SHIFT_4778_out0;
wire  [1:0] v$SHIFT_4779_out0;
wire  [1:0] v$SHIFT_5531_out0;
wire  [1:0] v$SHIFT_5532_out0;
wire  [1:0] v$SR_11838_out0;
wire  [1:0] v$SR_11839_out0;
wire  [1:0] v$SR_11840_out0;
wire  [1:0] v$SR_11841_out0;
wire  [1:0] v$SR_11842_out0;
wire  [1:0] v$SR_11843_out0;
wire  [1:0] v$SR_11844_out0;
wire  [1:0] v$SR_11845_out0;
wire  [1:0] v$SR_3024_out0;
wire  [1:0] v$SR_3025_out0;
wire  [1:0] v$SR_3026_out0;
wire  [1:0] v$SR_3027_out0;
wire  [1:0] v$SR_3028_out0;
wire  [1:0] v$SR_3029_out0;
wire  [1:0] v$SR_3030_out0;
wire  [1:0] v$SR_3031_out0;
wire  [1:0] v$SR_6654_out0;
wire  [1:0] v$SR_6655_out0;
wire  [1:0] v$XOR1_3401_out0;
wire  [1:0] v$XOR1_3402_out0;
wire  [1:0] v$XOR1_5800_out0;
wire  [1:0] v$XOR1_5801_out0;
wire  [1:0] v$XOR2_13161_out0;
wire  [1:0] v$XOR2_13162_out0;
wire  [1:0] v$XOR3_2754_out0;
wire  [1:0] v$XOR3_2755_out0;
wire  [1:0] v$Y_4474_out0;
wire  [1:0] v$Y_4475_out0;
wire  [1:0] v$Y_4476_out0;
wire  [1:0] v$Y_4477_out0;
wire  [1:0] v$Y_4478_out0;
wire  [1:0] v$Y_4479_out0;
wire  [1:0] v$Y_4480_out0;
wire  [1:0] v$Y_4481_out0;
wire  [1:0] v$Y_4482_out0;
wire  [1:0] v$Y_4483_out0;
wire  [1:0] v$Y_4484_out0;
wire  [1:0] v$Y_4485_out0;
wire  [1:0] v$Y_4486_out0;
wire  [1:0] v$Y_4487_out0;
wire  [1:0] v$Y_4488_out0;
wire  [1:0] v$Y_4489_out0;
wire  [1:0] v$Y_4490_out0;
wire  [1:0] v$Y_4491_out0;
wire  [1:0] v$Y_4492_out0;
wire  [1:0] v$Y_4493_out0;
wire  [1:0] v$Y_4494_out0;
wire  [1:0] v$Y_4495_out0;
wire  [1:0] v$Y_4496_out0;
wire  [1:0] v$Y_4497_out0;
wire  [1:0] v$Y_4498_out0;
wire  [1:0] v$Y_4499_out0;
wire  [1:0] v$Y_4500_out0;
wire  [1:0] v$Y_4501_out0;
wire  [1:0] v$Y_4502_out0;
wire  [1:0] v$Y_4503_out0;
wire  [1:0] v$Y_4504_out0;
wire  [1:0] v$Y_4505_out0;
wire  [1:0] v$Y_4506_out0;
wire  [1:0] v$Y_4507_out0;
wire  [1:0] v$Y_4508_out0;
wire  [1:0] v$Y_4509_out0;
wire  [1:0] v$Y_4510_out0;
wire  [1:0] v$Y_4511_out0;
wire  [1:0] v$Y_4512_out0;
wire  [1:0] v$Y_4513_out0;
wire  [1:0] v$Y_4514_out0;
wire  [1:0] v$Y_4515_out0;
wire  [1:0] v$Y_4516_out0;
wire  [1:0] v$Y_4517_out0;
wire  [1:0] v$Y_4518_out0;
wire  [1:0] v$Y_4519_out0;
wire  [1:0] v$Y_4520_out0;
wire  [1:0] v$Y_4521_out0;
wire  [1:0] v$Y_4522_out0;
wire  [1:0] v$Y_4523_out0;
wire  [1:0] v$Y_4524_out0;
wire  [1:0] v$Y_4525_out0;
wire  [1:0] v$Y_4526_out0;
wire  [1:0] v$Y_4527_out0;
wire  [1:0] v$Y_4528_out0;
wire  [1:0] v$Y_4529_out0;
wire  [1:0] v$Y_4530_out0;
wire  [1:0] v$Y_4531_out0;
wire  [1:0] v$Y_4532_out0;
wire  [1:0] v$Y_4533_out0;
wire  [1:0] v$_1005_out0;
wire  [1:0] v$_1006_out0;
wire  [1:0] v$_10125_out0;
wire  [1:0] v$_10126_out0;
wire  [1:0] v$_10228_out0;
wire  [1:0] v$_10229_out0;
wire  [1:0] v$_10329_out0;
wire  [1:0] v$_10329_out1;
wire  [1:0] v$_10330_out0;
wire  [1:0] v$_10330_out1;
wire  [1:0] v$_10615_out0;
wire  [1:0] v$_10616_out0;
wire  [1:0] v$_11128_out0;
wire  [1:0] v$_11129_out0;
wire  [1:0] v$_11152_out0;
wire  [1:0] v$_11153_out0;
wire  [1:0] v$_11188_out0;
wire  [1:0] v$_11189_out0;
wire  [1:0] v$_11300_out0;
wire  [1:0] v$_11301_out0;
wire  [1:0] v$_11387_out0;
wire  [1:0] v$_11387_out1;
wire  [1:0] v$_11388_out0;
wire  [1:0] v$_11388_out1;
wire  [1:0] v$_11788_out0;
wire  [1:0] v$_11789_out0;
wire  [1:0] v$_11823_out0;
wire  [1:0] v$_11824_out0;
wire  [1:0] v$_1185_out0;
wire  [1:0] v$_1186_out0;
wire  [1:0] v$_12106_out0;
wire  [1:0] v$_12107_out0;
wire  [1:0] v$_1213_out0;
wire  [1:0] v$_1213_out1;
wire  [1:0] v$_1214_out0;
wire  [1:0] v$_1214_out1;
wire  [1:0] v$_12735_out0;
wire  [1:0] v$_12736_out0;
wire  [1:0] v$_13007_out1;
wire  [1:0] v$_13008_out1;
wire  [1:0] v$_13026_out0;
wire  [1:0] v$_13027_out0;
wire  [1:0] v$_13097_out0;
wire  [1:0] v$_13098_out0;
wire  [1:0] v$_13175_out0;
wire  [1:0] v$_13176_out0;
wire  [1:0] v$_13213_out0;
wire  [1:0] v$_13214_out0;
wire  [1:0] v$_1571_out0;
wire  [1:0] v$_1572_out0;
wire  [1:0] v$_1879_out0;
wire  [1:0] v$_1880_out0;
wire  [1:0] v$_192_out0;
wire  [1:0] v$_192_out1;
wire  [1:0] v$_193_out0;
wire  [1:0] v$_193_out1;
wire  [1:0] v$_199_out0;
wire  [1:0] v$_199_out1;
wire  [1:0] v$_200_out0;
wire  [1:0] v$_200_out1;
wire  [1:0] v$_2415_out0;
wire  [1:0] v$_2415_out1;
wire  [1:0] v$_2416_out0;
wire  [1:0] v$_2416_out1;
wire  [1:0] v$_2493_out0;
wire  [1:0] v$_2494_out0;
wire  [1:0] v$_3459_out0;
wire  [1:0] v$_3460_out0;
wire  [1:0] v$_3516_out0;
wire  [1:0] v$_3516_out1;
wire  [1:0] v$_3517_out0;
wire  [1:0] v$_3517_out1;
wire  [1:0] v$_4077_out1;
wire  [1:0] v$_4078_out1;
wire  [1:0] v$_414_out0;
wire  [1:0] v$_415_out0;
wire  [1:0] v$_4200_out0;
wire  [1:0] v$_4201_out0;
wire  [1:0] v$_4267_out0;
wire  [1:0] v$_4268_out0;
wire  [1:0] v$_4269_out0;
wire  [1:0] v$_4270_out0;
wire  [1:0] v$_4271_out0;
wire  [1:0] v$_4272_out0;
wire  [1:0] v$_4273_out0;
wire  [1:0] v$_4274_out0;
wire  [1:0] v$_4275_out0;
wire  [1:0] v$_4276_out0;
wire  [1:0] v$_4277_out0;
wire  [1:0] v$_4278_out0;
wire  [1:0] v$_4279_out0;
wire  [1:0] v$_4280_out0;
wire  [1:0] v$_4281_out0;
wire  [1:0] v$_4282_out0;
wire  [1:0] v$_4283_out0;
wire  [1:0] v$_4284_out0;
wire  [1:0] v$_4285_out0;
wire  [1:0] v$_4286_out0;
wire  [1:0] v$_4287_out0;
wire  [1:0] v$_4288_out0;
wire  [1:0] v$_4289_out0;
wire  [1:0] v$_4290_out0;
wire  [1:0] v$_4291_out0;
wire  [1:0] v$_4292_out0;
wire  [1:0] v$_4293_out0;
wire  [1:0] v$_4294_out0;
wire  [1:0] v$_4295_out0;
wire  [1:0] v$_4296_out0;
wire  [1:0] v$_4297_out0;
wire  [1:0] v$_4298_out0;
wire  [1:0] v$_4299_out0;
wire  [1:0] v$_4300_out0;
wire  [1:0] v$_4301_out0;
wire  [1:0] v$_4302_out0;
wire  [1:0] v$_4303_out0;
wire  [1:0] v$_4304_out0;
wire  [1:0] v$_4305_out0;
wire  [1:0] v$_4306_out0;
wire  [1:0] v$_4307_out0;
wire  [1:0] v$_4308_out0;
wire  [1:0] v$_4309_out0;
wire  [1:0] v$_4310_out0;
wire  [1:0] v$_4311_out0;
wire  [1:0] v$_4312_out0;
wire  [1:0] v$_4313_out0;
wire  [1:0] v$_4314_out0;
wire  [1:0] v$_4315_out0;
wire  [1:0] v$_4316_out0;
wire  [1:0] v$_4317_out0;
wire  [1:0] v$_4318_out0;
wire  [1:0] v$_4319_out0;
wire  [1:0] v$_4320_out0;
wire  [1:0] v$_4321_out0;
wire  [1:0] v$_4322_out0;
wire  [1:0] v$_4323_out0;
wire  [1:0] v$_4324_out0;
wire  [1:0] v$_4325_out0;
wire  [1:0] v$_4326_out0;
wire  [1:0] v$_4973_out0;
wire  [1:0] v$_4973_out1;
wire  [1:0] v$_4974_out0;
wire  [1:0] v$_4974_out1;
wire  [1:0] v$_5044_out0;
wire  [1:0] v$_5044_out1;
wire  [1:0] v$_5045_out0;
wire  [1:0] v$_5045_out1;
wire  [1:0] v$_50_out0;
wire  [1:0] v$_50_out1;
wire  [1:0] v$_51_out0;
wire  [1:0] v$_51_out1;
wire  [1:0] v$_525_out0;
wire  [1:0] v$_526_out0;
wire  [1:0] v$_5279_out0;
wire  [1:0] v$_5280_out0;
wire  [1:0] v$_5700_out0;
wire  [1:0] v$_5700_out1;
wire  [1:0] v$_5701_out0;
wire  [1:0] v$_5701_out1;
wire  [1:0] v$_5908_out0;
wire  [1:0] v$_5908_out1;
wire  [1:0] v$_5909_out0;
wire  [1:0] v$_5909_out1;
wire  [1:0] v$_5910_out0;
wire  [1:0] v$_5910_out1;
wire  [1:0] v$_5911_out0;
wire  [1:0] v$_5911_out1;
wire  [1:0] v$_5912_out0;
wire  [1:0] v$_5912_out1;
wire  [1:0] v$_5913_out0;
wire  [1:0] v$_5913_out1;
wire  [1:0] v$_5914_out0;
wire  [1:0] v$_5914_out1;
wire  [1:0] v$_5915_out0;
wire  [1:0] v$_5915_out1;
wire  [1:0] v$_5916_out0;
wire  [1:0] v$_5916_out1;
wire  [1:0] v$_5917_out0;
wire  [1:0] v$_5917_out1;
wire  [1:0] v$_5918_out0;
wire  [1:0] v$_5918_out1;
wire  [1:0] v$_5919_out0;
wire  [1:0] v$_5919_out1;
wire  [1:0] v$_6415_out0;
wire  [1:0] v$_6415_out1;
wire  [1:0] v$_6416_out0;
wire  [1:0] v$_6416_out1;
wire  [1:0] v$_6431_out0;
wire  [1:0] v$_6432_out0;
wire  [1:0] v$_6453_out0;
wire  [1:0] v$_6454_out0;
wire  [1:0] v$_6643_out0;
wire  [1:0] v$_6644_out0;
wire  [1:0] v$_6649_out0;
wire  [1:0] v$_6650_out0;
wire  [1:0] v$_705_out0;
wire  [1:0] v$_705_out1;
wire  [1:0] v$_706_out0;
wire  [1:0] v$_706_out1;
wire  [1:0] v$_7098_out0;
wire  [1:0] v$_7099_out0;
wire  [1:0] v$_7112_out0;
wire  [1:0] v$_7112_out1;
wire  [1:0] v$_7113_out0;
wire  [1:0] v$_7113_out1;
wire  [1:0] v$_7233_out0;
wire  [1:0] v$_7234_out0;
wire  [1:0] v$_7616_out0;
wire  [1:0] v$_7616_out1;
wire  [1:0] v$_7617_out0;
wire  [1:0] v$_7617_out1;
wire  [1:0] v$_807_out0;
wire  [1:0] v$_807_out1;
wire  [1:0] v$_808_out0;
wire  [1:0] v$_808_out1;
wire  [1:0] v$_8484_out0;
wire  [1:0] v$_8484_out1;
wire  [1:0] v$_8485_out0;
wire  [1:0] v$_8485_out1;
wire  [1:0] v$_8486_out0;
wire  [1:0] v$_8486_out1;
wire  [1:0] v$_8487_out0;
wire  [1:0] v$_8487_out1;
wire  [1:0] v$_8488_out0;
wire  [1:0] v$_8488_out1;
wire  [1:0] v$_8489_out0;
wire  [1:0] v$_8489_out1;
wire  [1:0] v$_8490_out0;
wire  [1:0] v$_8490_out1;
wire  [1:0] v$_8491_out0;
wire  [1:0] v$_8491_out1;
wire  [1:0] v$_8492_out0;
wire  [1:0] v$_8492_out1;
wire  [1:0] v$_8493_out0;
wire  [1:0] v$_8493_out1;
wire  [1:0] v$_8494_out0;
wire  [1:0] v$_8494_out1;
wire  [1:0] v$_8495_out0;
wire  [1:0] v$_8495_out1;
wire  [1:0] v$_8688_out0;
wire  [1:0] v$_8689_out0;
wire  [1:0] v$_8764_out0;
wire  [1:0] v$_8764_out1;
wire  [1:0] v$_8765_out0;
wire  [1:0] v$_8765_out1;
wire  [1:0] v$_8810_out0;
wire  [1:0] v$_8811_out0;
wire  [1:0] v$_8844_out0;
wire  [1:0] v$_8844_out1;
wire  [1:0] v$_8845_out0;
wire  [1:0] v$_8845_out1;
wire  [1:0] v$_885_out0;
wire  [1:0] v$_885_out1;
wire  [1:0] v$_8866_out0;
wire  [1:0] v$_8866_out1;
wire  [1:0] v$_8867_out0;
wire  [1:0] v$_8867_out1;
wire  [1:0] v$_886_out0;
wire  [1:0] v$_886_out1;
wire  [1:0] v$_8872_out1;
wire  [1:0] v$_8873_out1;
wire  [1:0] v$_8980_out0;
wire  [1:0] v$_8981_out0;
wire  [1:0] v$_9552_out0;
wire  [1:0] v$_9553_out0;
wire  [1:0] v$_9554_out0;
wire  [1:0] v$_9555_out0;
wire  [1:0] v$_9609_out0;
wire  [1:0] v$_9610_out0;
wire  [1:0] v$_9984_out0;
wire  [1:0] v$_9985_out0;
wire  [21:0] v$SEL1_10682_out0;
wire  [21:0] v$SEL1_10699_out0;
wire  [21:0] v$SEL1_10704_out0;
wire  [21:0] v$SEL1_10709_out0;
wire  [21:0] v$SEL1_10714_out0;
wire  [21:0] v$SEL1_10731_out0;
wire  [21:0] v$SEL1_10736_out0;
wire  [21:0] v$SEL1_10741_out0;
wire  [21:0] v$SEL1_5938_out0;
wire  [21:0] v$SEL1_5955_out0;
wire  [21:0] v$SEL1_5960_out0;
wire  [21:0] v$SEL1_5965_out0;
wire  [21:0] v$SEL1_5970_out0;
wire  [21:0] v$SEL1_5987_out0;
wire  [21:0] v$SEL1_5992_out0;
wire  [21:0] v$SEL1_5997_out0;
wire  [22:0] v$A$MANTISA$MUL_1556_out0;
wire  [22:0] v$A$MANTISA$MUL_1557_out0;
wire  [22:0] v$A$MANTISA_12691_out0;
wire  [22:0] v$A$MANTISA_12692_out0;
wire  [22:0] v$A$MANTISA_7625_out0;
wire  [22:0] v$A$MANTISA_7626_out0;
wire  [22:0] v$A$MANTISA_9937_out0;
wire  [22:0] v$A$MANTISA_9938_out0;
wire  [22:0] v$B$MANTISA$MUL_5662_out0;
wire  [22:0] v$B$MANTISA$MUL_5663_out0;
wire  [22:0] v$B$MANTISA_1763_out0;
wire  [22:0] v$B$MANTISA_1764_out0;
wire  [22:0] v$B$MANTISA_2780_out0;
wire  [22:0] v$B$MANTISA_2781_out0;
wire  [22:0] v$B$MANTISA_3300_out0;
wire  [22:0] v$B$MANTISA_3301_out0;
wire  [22:0] v$C5_10888_out0;
wire  [22:0] v$C5_10889_out0;
wire  [22:0] v$MANTISA$ADDITION_8782_out0;
wire  [22:0] v$MANTISA$ADDITION_8783_out0;
wire  [22:0] v$MANTISA$RESULT$BEFORE$MERGE_13345_out0;
wire  [22:0] v$MANTISA$RESULT$BEFORE$MERGE_13346_out0;
wire  [22:0] v$MANTISA$RESULT$FPU$ADDER_7690_out0;
wire  [22:0] v$MANTISA$RESULT$FPU$ADDER_7691_out0;
wire  [22:0] v$MANTISA$RESULT_4552_out0;
wire  [22:0] v$MANTISA$RESULT_4553_out0;
wire  [22:0] v$MUX1_1084_out0;
wire  [22:0] v$MUX1_1085_out0;
wire  [22:0] v$MUX2_1734_out0;
wire  [22:0] v$MUX2_1735_out0;
wire  [22:0] v$MUX2_813_out0;
wire  [22:0] v$MUX2_814_out0;
wire  [22:0] v$MUX6_8424_out0;
wire  [22:0] v$MUX6_8425_out0;
wire  [22:0] v$MUX7_8395_out0;
wire  [22:0] v$MUX7_8396_out0;
wire  [22:0] v$MUX8_4811_out0;
wire  [22:0] v$MUX8_4812_out0;
wire  [22:0] v$OUT1_6958_out0;
wire  [22:0] v$OUT1_6959_out0;
wire  [22:0] v$SEL1_10680_out0;
wire  [22:0] v$SEL1_10697_out0;
wire  [22:0] v$SEL1_10702_out0;
wire  [22:0] v$SEL1_10707_out0;
wire  [22:0] v$SEL1_10712_out0;
wire  [22:0] v$SEL1_10729_out0;
wire  [22:0] v$SEL1_10734_out0;
wire  [22:0] v$SEL1_10739_out0;
wire  [22:0] v$SEL1_10991_out0;
wire  [22:0] v$SEL1_10992_out0;
wire  [22:0] v$SEL1_5936_out0;
wire  [22:0] v$SEL1_5953_out0;
wire  [22:0] v$SEL1_5958_out0;
wire  [22:0] v$SEL1_5963_out0;
wire  [22:0] v$SEL1_5968_out0;
wire  [22:0] v$SEL1_5985_out0;
wire  [22:0] v$SEL1_5990_out0;
wire  [22:0] v$SEL1_5995_out0;
wire  [22:0] v$SEL1_9750_out0;
wire  [22:0] v$SEL1_9751_out0;
wire  [22:0] v$SEL2_4035_out0;
wire  [22:0] v$SEL2_4036_out0;
wire  [22:0] v$SEL2_5606_out0;
wire  [22:0] v$SEL2_5608_out0;
wire  [22:0] v$SEL2_7265_out0;
wire  [22:0] v$SEL2_7266_out0;
wire  [22:0] v$SEL3_7684_out0;
wire  [22:0] v$SEL3_7685_out0;
wire  [22:0] v$SEL3_9646_out0;
wire  [22:0] v$SEL3_9647_out0;
wire  [22:0] v$SEL4_1201_out0;
wire  [22:0] v$SEL4_1202_out0;
wire  [22:0] v$SEL4_8615_out0;
wire  [22:0] v$SEL4_8616_out0;
wire  [22:0] v$SEL6_3085_out0;
wire  [22:0] v$SEL6_3086_out0;
wire  [22:0] v$SEL8_12288_out0;
wire  [22:0] v$SEL8_12289_out0;
wire  [22:0] v$SEL8_12465_out0;
wire  [22:0] v$SEL8_12466_out0;
wire  [22:0] v$SEL8_12467_out0;
wire  [22:0] v$SEL8_12468_out0;
wire  [22:0] v$SEL8_12469_out0;
wire  [22:0] v$SEL8_12470_out0;
wire  [22:0] v$SEL8_12471_out0;
wire  [22:0] v$SEL8_12472_out0;
wire  [22:0] v$SEL8_12473_out0;
wire  [22:0] v$SEL8_12474_out0;
wire  [22:0] v$SEL8_12475_out0;
wire  [22:0] v$SEL8_12476_out0;
wire  [22:0] v$SEL8_12477_out0;
wire  [22:0] v$SEL8_12478_out0;
wire  [22:0] v$SEL8_12479_out0;
wire  [22:0] v$SEL8_12480_out0;
wire  [22:0] v$SEL8_12481_out0;
wire  [22:0] v$SEL8_12482_out0;
wire  [22:0] v$SEL8_12483_out0;
wire  [22:0] v$SEL8_12484_out0;
wire  [22:0] v$SEL8_12485_out0;
wire  [22:0] v$SEL8_12486_out0;
wire  [22:0] v$SEL8_12487_out0;
wire  [22:0] v$SEL8_12488_out0;
wire  [22:0] v$SEL8_4873_out0;
wire  [22:0] v$SEL8_4874_out0;
wire  [22:0] v$_11393_out0;
wire  [22:0] v$_11394_out0;
wire  [22:0] v$_1158_out0;
wire  [22:0] v$_1159_out0;
wire  [22:0] v$_12839_out0;
wire  [22:0] v$_12840_out0;
wire  [22:0] v$_879_out0;
wire  [22:0] v$_880_out0;
wire  [23:0] v$A$MANTISA$COMPARATOR_5072_out0;
wire  [23:0] v$A$MANTISA$COMPARATOR_5073_out0;
wire  [23:0] v$A$MANTISA_2469_out0;
wire  [23:0] v$A$MANTISA_2470_out0;
wire  [23:0] v$A$MANTISSA_8789_out0;
wire  [23:0] v$A$MANTISSA_8790_out0;
wire  [23:0] v$A1_10523_out0;
wire  [23:0] v$A1_10524_out0;
wire  [23:0] v$A1_10525_out0;
wire  [23:0] v$A1_10526_out0;
wire  [23:0] v$A1_10527_out0;
wire  [23:0] v$A1_10528_out0;
wire  [23:0] v$A1_10529_out0;
wire  [23:0] v$A1_10530_out0;
wire  [23:0] v$A1_10531_out0;
wire  [23:0] v$A1_10532_out0;
wire  [23:0] v$A1_10533_out0;
wire  [23:0] v$A1_10534_out0;
wire  [23:0] v$A1_10535_out0;
wire  [23:0] v$A1_10536_out0;
wire  [23:0] v$A1_10537_out0;
wire  [23:0] v$A1_10538_out0;
wire  [23:0] v$A1_10539_out0;
wire  [23:0] v$A1_10540_out0;
wire  [23:0] v$A1_10541_out0;
wire  [23:0] v$A1_10542_out0;
wire  [23:0] v$A1_10543_out0;
wire  [23:0] v$A1_10544_out0;
wire  [23:0] v$A1_10545_out0;
wire  [23:0] v$A1_10546_out0;
wire  [23:0] v$A1_229_out0;
wire  [23:0] v$A1_230_out0;
wire  [23:0] v$A2_8371_out0;
wire  [23:0] v$A2_8372_out0;
wire  [23:0] v$ADDER$A_2411_out0;
wire  [23:0] v$ADDER$A_2412_out0;
wire  [23:0] v$ADDER$B_4449_out0;
wire  [23:0] v$ADDER$B_4450_out0;
wire  [23:0] v$A_10147_out0;
wire  [23:0] v$A_10148_out0;
wire  [23:0] v$A_3663_out0;
wire  [23:0] v$A_3664_out0;
wire  [23:0] v$B$MANTISA$COMPARATOR_11084_out0;
wire  [23:0] v$B$MANTISA$COMPARATOR_11085_out0;
wire  [23:0] v$B$MANTISA_10857_out0;
wire  [23:0] v$B$MANTISA_10858_out0;
wire  [23:0] v$B$MANTISSA_1575_out0;
wire  [23:0] v$B$MANTISSA_1576_out0;
wire  [23:0] v$B_1106_out0;
wire  [23:0] v$B_1107_out0;
wire  [23:0] v$B_5834_out0;
wire  [23:0] v$B_5835_out0;
wire  [23:0] v$C1_11389_out0;
wire  [23:0] v$C1_11390_out0;
wire  [23:0] v$C1_3093_out0;
wire  [23:0] v$C1_3094_out0;
wire  [23:0] v$C1_3095_out0;
wire  [23:0] v$C1_3096_out0;
wire  [23:0] v$C1_3097_out0;
wire  [23:0] v$C1_3098_out0;
wire  [23:0] v$C1_3099_out0;
wire  [23:0] v$C1_3100_out0;
wire  [23:0] v$C2_5340_out0;
wire  [23:0] v$C2_5341_out0;
wire  [23:0] v$C5_2672_out0;
wire  [23:0] v$C5_2673_out0;
wire  [23:0] v$C5_2674_out0;
wire  [23:0] v$C5_2675_out0;
wire  [23:0] v$C5_2676_out0;
wire  [23:0] v$C5_2677_out0;
wire  [23:0] v$C5_2678_out0;
wire  [23:0] v$C5_2679_out0;
wire  [23:0] v$C5_2680_out0;
wire  [23:0] v$C5_2681_out0;
wire  [23:0] v$C5_2682_out0;
wire  [23:0] v$C5_2683_out0;
wire  [23:0] v$C5_2684_out0;
wire  [23:0] v$C5_2685_out0;
wire  [23:0] v$C5_2686_out0;
wire  [23:0] v$C5_2687_out0;
wire  [23:0] v$C5_2688_out0;
wire  [23:0] v$C5_2689_out0;
wire  [23:0] v$C5_2690_out0;
wire  [23:0] v$C5_2691_out0;
wire  [23:0] v$C5_2692_out0;
wire  [23:0] v$C5_2693_out0;
wire  [23:0] v$C5_2694_out0;
wire  [23:0] v$C5_2695_out0;
wire  [23:0] v$C7_10012_out0;
wire  [23:0] v$C7_10013_out0;
wire  [23:0] v$C8_9178_out0;
wire  [23:0] v$C8_9179_out0;
wire  [23:0] v$C9_10581_out0;
wire  [23:0] v$C9_10582_out0;
wire  [23:0] v$IN_10872_out0;
wire  [23:0] v$IN_10875_out0;
wire  [23:0] v$IN_10876_out0;
wire  [23:0] v$IN_10877_out0;
wire  [23:0] v$IN_10878_out0;
wire  [23:0] v$IN_10881_out0;
wire  [23:0] v$IN_10882_out0;
wire  [23:0] v$IN_10883_out0;
wire  [23:0] v$IN_12747_out0;
wire  [23:0] v$IN_12748_out0;
wire  [23:0] v$IN_2566_out0;
wire  [23:0] v$IN_2573_out0;
wire  [23:0] v$IN_2574_out0;
wire  [23:0] v$IN_2575_out0;
wire  [23:0] v$IN_2576_out0;
wire  [23:0] v$IN_2583_out0;
wire  [23:0] v$IN_2584_out0;
wire  [23:0] v$IN_2585_out0;
wire  [23:0] v$IN_3411_out0;
wire  [23:0] v$IN_3412_out0;
wire  [23:0] v$IN_3415_out0;
wire  [23:0] v$IN_3416_out0;
wire  [23:0] v$IN_3417_out0;
wire  [23:0] v$IN_3418_out0;
wire  [23:0] v$IN_3419_out0;
wire  [23:0] v$IN_3420_out0;
wire  [23:0] v$IN_3421_out0;
wire  [23:0] v$IN_3422_out0;
wire  [23:0] v$IN_3425_out0;
wire  [23:0] v$IN_3426_out0;
wire  [23:0] v$IN_3427_out0;
wire  [23:0] v$IN_3428_out0;
wire  [23:0] v$IN_3429_out0;
wire  [23:0] v$IN_3430_out0;
wire  [23:0] v$IN_3521_out0;
wire  [23:0] v$IN_3522_out0;
wire  [23:0] v$IN_3523_out0;
wire  [23:0] v$IN_3524_out0;
wire  [23:0] v$IN_3525_out0;
wire  [23:0] v$IN_3538_out0;
wire  [23:0] v$IN_3539_out0;
wire  [23:0] v$IN_3540_out0;
wire  [23:0] v$IN_3541_out0;
wire  [23:0] v$IN_3542_out0;
wire  [23:0] v$IN_3543_out0;
wire  [23:0] v$IN_3544_out0;
wire  [23:0] v$IN_3545_out0;
wire  [23:0] v$IN_3546_out0;
wire  [23:0] v$IN_3547_out0;
wire  [23:0] v$IN_3548_out0;
wire  [23:0] v$IN_3549_out0;
wire  [23:0] v$IN_3550_out0;
wire  [23:0] v$IN_3551_out0;
wire  [23:0] v$IN_3552_out0;
wire  [23:0] v$IN_3553_out0;
wire  [23:0] v$IN_3554_out0;
wire  [23:0] v$IN_3555_out0;
wire  [23:0] v$IN_3556_out0;
wire  [23:0] v$IN_3557_out0;
wire  [23:0] v$IN_3570_out0;
wire  [23:0] v$IN_3571_out0;
wire  [23:0] v$IN_3572_out0;
wire  [23:0] v$IN_3573_out0;
wire  [23:0] v$IN_3574_out0;
wire  [23:0] v$IN_3575_out0;
wire  [23:0] v$IN_3576_out0;
wire  [23:0] v$IN_3577_out0;
wire  [23:0] v$IN_3578_out0;
wire  [23:0] v$IN_3579_out0;
wire  [23:0] v$IN_3580_out0;
wire  [23:0] v$IN_3581_out0;
wire  [23:0] v$IN_3582_out0;
wire  [23:0] v$IN_3583_out0;
wire  [23:0] v$IN_3584_out0;
wire  [23:0] v$IN_7582_out0;
wire  [23:0] v$IN_7585_out0;
wire  [23:0] v$IN_7586_out0;
wire  [23:0] v$IN_7587_out0;
wire  [23:0] v$IN_7588_out0;
wire  [23:0] v$IN_7591_out0;
wire  [23:0] v$IN_7592_out0;
wire  [23:0] v$IN_7593_out0;
wire  [23:0] v$IN_8774_out0;
wire  [23:0] v$IN_8775_out0;
wire  [23:0] v$IN_8776_out0;
wire  [23:0] v$IN_8777_out0;
wire  [23:0] v$IN_8778_out0;
wire  [23:0] v$IN_8779_out0;
wire  [23:0] v$IN_8780_out0;
wire  [23:0] v$IN_8781_out0;
wire  [23:0] v$LZD$INPUT_6076_out0;
wire  [23:0] v$LZD$INPUT_6077_out0;
wire  [23:0] v$MULTIPLIER_4366_out0;
wire  [23:0] v$MULTIPLIER_4367_out0;
wire  [23:0] v$MULTIPLIER_4368_out0;
wire  [23:0] v$MULTIPLIER_4369_out0;
wire  [23:0] v$MULTIPLIER_4370_out0;
wire  [23:0] v$MULTIPLIER_4371_out0;
wire  [23:0] v$MULTIPLIER_4372_out0;
wire  [23:0] v$MULTIPLIER_4373_out0;
wire  [23:0] v$MULTIPLIER_4374_out0;
wire  [23:0] v$MULTIPLIER_4375_out0;
wire  [23:0] v$MULTIPLIER_4376_out0;
wire  [23:0] v$MULTIPLIER_4377_out0;
wire  [23:0] v$MULTIPLIER_4378_out0;
wire  [23:0] v$MULTIPLIER_4379_out0;
wire  [23:0] v$MULTIPLIER_4380_out0;
wire  [23:0] v$MULTIPLIER_4381_out0;
wire  [23:0] v$MULTIPLIER_4382_out0;
wire  [23:0] v$MULTIPLIER_4383_out0;
wire  [23:0] v$MULTIPLIER_4384_out0;
wire  [23:0] v$MULTIPLIER_4385_out0;
wire  [23:0] v$MULTIPLIER_4386_out0;
wire  [23:0] v$MULTIPLIER_4387_out0;
wire  [23:0] v$MULTIPLIER_4388_out0;
wire  [23:0] v$MULTIPLIER_4389_out0;
wire  [23:0] v$MUX1_1283_out0;
wire  [23:0] v$MUX1_1284_out0;
wire  [23:0] v$MUX1_1285_out0;
wire  [23:0] v$MUX1_1286_out0;
wire  [23:0] v$MUX1_1287_out0;
wire  [23:0] v$MUX1_1300_out0;
wire  [23:0] v$MUX1_1301_out0;
wire  [23:0] v$MUX1_1302_out0;
wire  [23:0] v$MUX1_1303_out0;
wire  [23:0] v$MUX1_1304_out0;
wire  [23:0] v$MUX1_1305_out0;
wire  [23:0] v$MUX1_1306_out0;
wire  [23:0] v$MUX1_1307_out0;
wire  [23:0] v$MUX1_1308_out0;
wire  [23:0] v$MUX1_1309_out0;
wire  [23:0] v$MUX1_1310_out0;
wire  [23:0] v$MUX1_1311_out0;
wire  [23:0] v$MUX1_1312_out0;
wire  [23:0] v$MUX1_1313_out0;
wire  [23:0] v$MUX1_1314_out0;
wire  [23:0] v$MUX1_1315_out0;
wire  [23:0] v$MUX1_1316_out0;
wire  [23:0] v$MUX1_1317_out0;
wire  [23:0] v$MUX1_1318_out0;
wire  [23:0] v$MUX1_1319_out0;
wire  [23:0] v$MUX1_1332_out0;
wire  [23:0] v$MUX1_1333_out0;
wire  [23:0] v$MUX1_1334_out0;
wire  [23:0] v$MUX1_1335_out0;
wire  [23:0] v$MUX1_1336_out0;
wire  [23:0] v$MUX1_1337_out0;
wire  [23:0] v$MUX1_1338_out0;
wire  [23:0] v$MUX1_1339_out0;
wire  [23:0] v$MUX1_1340_out0;
wire  [23:0] v$MUX1_1341_out0;
wire  [23:0] v$MUX1_1342_out0;
wire  [23:0] v$MUX1_1343_out0;
wire  [23:0] v$MUX1_1344_out0;
wire  [23:0] v$MUX1_1345_out0;
wire  [23:0] v$MUX1_1346_out0;
wire  [23:0] v$MUX1_5806_out0;
wire  [23:0] v$MUX1_5807_out0;
wire  [23:0] v$MUX1_5808_out0;
wire  [23:0] v$MUX1_5809_out0;
wire  [23:0] v$MUX1_5810_out0;
wire  [23:0] v$MUX1_5811_out0;
wire  [23:0] v$MUX1_5812_out0;
wire  [23:0] v$MUX1_5813_out0;
wire  [23:0] v$MUX1_5814_out0;
wire  [23:0] v$MUX1_5815_out0;
wire  [23:0] v$MUX1_5816_out0;
wire  [23:0] v$MUX1_5817_out0;
wire  [23:0] v$MUX1_5818_out0;
wire  [23:0] v$MUX1_5819_out0;
wire  [23:0] v$MUX1_5820_out0;
wire  [23:0] v$MUX1_5821_out0;
wire  [23:0] v$MUX1_5822_out0;
wire  [23:0] v$MUX1_5823_out0;
wire  [23:0] v$MUX1_5824_out0;
wire  [23:0] v$MUX1_5825_out0;
wire  [23:0] v$MUX1_5826_out0;
wire  [23:0] v$MUX1_5827_out0;
wire  [23:0] v$MUX1_5828_out0;
wire  [23:0] v$MUX1_5829_out0;
wire  [23:0] v$MUX1_7471_out0;
wire  [23:0] v$MUX1_7472_out0;
wire  [23:0] v$MUX1_7473_out0;
wire  [23:0] v$MUX1_7474_out0;
wire  [23:0] v$MUX1_7475_out0;
wire  [23:0] v$MUX1_7476_out0;
wire  [23:0] v$MUX1_7477_out0;
wire  [23:0] v$MUX1_7478_out0;
wire  [23:0] v$MUX1_9571_out0;
wire  [23:0] v$MUX1_9572_out0;
wire  [23:0] v$MUX2_10555_out0;
wire  [23:0] v$MUX2_10558_out0;
wire  [23:0] v$MUX2_10559_out0;
wire  [23:0] v$MUX2_10560_out0;
wire  [23:0] v$MUX2_10561_out0;
wire  [23:0] v$MUX2_10564_out0;
wire  [23:0] v$MUX2_10565_out0;
wire  [23:0] v$MUX2_10566_out0;
wire  [23:0] v$MUX2_12807_out0;
wire  [23:0] v$MUX2_12808_out0;
wire  [23:0] v$MUX2_13217_out0;
wire  [23:0] v$MUX2_13224_out0;
wire  [23:0] v$MUX2_13225_out0;
wire  [23:0] v$MUX2_13226_out0;
wire  [23:0] v$MUX2_13227_out0;
wire  [23:0] v$MUX2_13234_out0;
wire  [23:0] v$MUX2_13235_out0;
wire  [23:0] v$MUX2_13236_out0;
wire  [23:0] v$MUX2_1393_out0;
wire  [23:0] v$MUX2_1396_out0;
wire  [23:0] v$MUX2_1397_out0;
wire  [23:0] v$MUX2_1398_out0;
wire  [23:0] v$MUX2_1399_out0;
wire  [23:0] v$MUX2_1402_out0;
wire  [23:0] v$MUX2_1403_out0;
wire  [23:0] v$MUX2_1404_out0;
wire  [23:0] v$MUX2_1405_out0;
wire  [23:0] v$MUX2_1406_out0;
wire  [23:0] v$MUX2_1409_out0;
wire  [23:0] v$MUX2_1410_out0;
wire  [23:0] v$MUX2_1411_out0;
wire  [23:0] v$MUX2_1412_out0;
wire  [23:0] v$MUX2_1413_out0;
wire  [23:0] v$MUX2_1414_out0;
wire  [23:0] v$MUX2_1415_out0;
wire  [23:0] v$MUX2_1416_out0;
wire  [23:0] v$MUX2_1419_out0;
wire  [23:0] v$MUX2_1420_out0;
wire  [23:0] v$MUX2_1421_out0;
wire  [23:0] v$MUX2_1422_out0;
wire  [23:0] v$MUX2_1423_out0;
wire  [23:0] v$MUX2_1424_out0;
wire  [23:0] v$MUX3_1862_out0;
wire  [23:0] v$MUX3_1863_out0;
wire  [23:0] v$MUX3_2479_out0;
wire  [23:0] v$MUX3_2480_out0;
wire  [23:0] v$MUX3_5173_out0;
wire  [23:0] v$MUX3_5174_out0;
wire  [23:0] v$MUX3_8454_out0;
wire  [23:0] v$MUX3_8455_out0;
wire  [23:0] v$MUX4_12976_out0;
wire  [23:0] v$MUX4_12977_out0;
wire  [23:0] v$MUX4_3912_out0;
wire  [23:0] v$MUX4_3913_out0;
wire  [23:0] v$MUX5_4229_out0;
wire  [23:0] v$MUX5_4230_out0;
wire  [23:0] v$MUX5_815_out0;
wire  [23:0] v$MUX5_816_out0;
wire  [23:0] v$MUX7_1979_out0;
wire  [23:0] v$MUX7_1980_out0;
wire  [23:0] v$MUX8_3643_out0;
wire  [23:0] v$MUX8_3644_out0;
wire  [23:0] v$MUX9_1381_out0;
wire  [23:0] v$MUX9_1382_out0;
wire  [23:0] v$OP1$MANTISA$ADDER_2346_out0;
wire  [23:0] v$OP1$MANTISA$ADDER_2347_out0;
wire  [23:0] v$OP1$MANTISA$MULTIPLY_7682_out0;
wire  [23:0] v$OP1$MANTISA$MULTIPLY_7683_out0;
wire  [23:0] v$OP1$MANTISA_2497_out0;
wire  [23:0] v$OP1$MANTISA_2498_out0;
wire  [23:0] v$OP1$MANTISA_6355_out0;
wire  [23:0] v$OP1$MANTISA_6356_out0;
wire  [23:0] v$OP1$MANTISA_7606_out0;
wire  [23:0] v$OP1$MANTISA_7607_out0;
wire  [23:0] v$OP1_2073_out0;
wire  [23:0] v$OP1_2074_out0;
wire  [23:0] v$OP1_2075_out0;
wire  [23:0] v$OP1_2076_out0;
wire  [23:0] v$OP1_2077_out0;
wire  [23:0] v$OP1_2078_out0;
wire  [23:0] v$OP1_2079_out0;
wire  [23:0] v$OP1_2080_out0;
wire  [23:0] v$OP1_2081_out0;
wire  [23:0] v$OP1_2082_out0;
wire  [23:0] v$OP1_2083_out0;
wire  [23:0] v$OP1_2084_out0;
wire  [23:0] v$OP1_2085_out0;
wire  [23:0] v$OP1_2086_out0;
wire  [23:0] v$OP1_2087_out0;
wire  [23:0] v$OP1_2088_out0;
wire  [23:0] v$OP1_2089_out0;
wire  [23:0] v$OP1_2090_out0;
wire  [23:0] v$OP1_2091_out0;
wire  [23:0] v$OP1_2092_out0;
wire  [23:0] v$OP1_2093_out0;
wire  [23:0] v$OP1_2094_out0;
wire  [23:0] v$OP1_2095_out0;
wire  [23:0] v$OP1_2096_out0;
wire  [23:0] v$OP1_2798_out0;
wire  [23:0] v$OP1_2799_out0;
wire  [23:0] v$OP1_9573_out0;
wire  [23:0] v$OP1_9574_out0;
wire  [23:0] v$OP1_9575_out0;
wire  [23:0] v$OP1_9576_out0;
wire  [23:0] v$OP1_9577_out0;
wire  [23:0] v$OP1_9578_out0;
wire  [23:0] v$OP1_9579_out0;
wire  [23:0] v$OP1_9580_out0;
wire  [23:0] v$OP1_9581_out0;
wire  [23:0] v$OP1_9582_out0;
wire  [23:0] v$OP1_9583_out0;
wire  [23:0] v$OP1_9584_out0;
wire  [23:0] v$OP1_9585_out0;
wire  [23:0] v$OP1_9586_out0;
wire  [23:0] v$OP1_9587_out0;
wire  [23:0] v$OP1_9588_out0;
wire  [23:0] v$OP1_9589_out0;
wire  [23:0] v$OP1_9590_out0;
wire  [23:0] v$OP1_9591_out0;
wire  [23:0] v$OP1_9592_out0;
wire  [23:0] v$OP1_9593_out0;
wire  [23:0] v$OP1_9594_out0;
wire  [23:0] v$OP1_9595_out0;
wire  [23:0] v$OP1_9596_out0;
wire  [23:0] v$OP2$MANTISA$ADDER_5066_out0;
wire  [23:0] v$OP2$MANTISA$ADDER_5067_out0;
wire  [23:0] v$OP2$MANTISA$MULTIPLY_1385_out0;
wire  [23:0] v$OP2$MANTISA$MULTIPLY_1386_out0;
wire  [23:0] v$OP2$MANTISA_1558_out0;
wire  [23:0] v$OP2$MANTISA_1559_out0;
wire  [23:0] v$OP2$MANTISA_2212_out0;
wire  [23:0] v$OP2$MANTISA_2213_out0;
wire  [23:0] v$OP2$MANTISA_6520_out0;
wire  [23:0] v$OP2$MANTISA_6521_out0;
wire  [23:0] v$OP2_2372_out0;
wire  [23:0] v$OP2_2373_out0;
wire  [23:0] v$OP2_2374_out0;
wire  [23:0] v$OP2_2375_out0;
wire  [23:0] v$OP2_2376_out0;
wire  [23:0] v$OP2_2377_out0;
wire  [23:0] v$OP2_2378_out0;
wire  [23:0] v$OP2_2379_out0;
wire  [23:0] v$OP2_2380_out0;
wire  [23:0] v$OP2_2381_out0;
wire  [23:0] v$OP2_2382_out0;
wire  [23:0] v$OP2_2383_out0;
wire  [23:0] v$OP2_2384_out0;
wire  [23:0] v$OP2_2385_out0;
wire  [23:0] v$OP2_2386_out0;
wire  [23:0] v$OP2_2387_out0;
wire  [23:0] v$OP2_2388_out0;
wire  [23:0] v$OP2_2389_out0;
wire  [23:0] v$OP2_2390_out0;
wire  [23:0] v$OP2_2391_out0;
wire  [23:0] v$OP2_2392_out0;
wire  [23:0] v$OP2_2393_out0;
wire  [23:0] v$OP2_2394_out0;
wire  [23:0] v$OP2_2395_out0;
wire  [23:0] v$OP2_2852_out0;
wire  [23:0] v$OP2_2853_out0;
wire  [23:0] v$OP2_6911_out0;
wire  [23:0] v$OP2_6912_out0;
wire  [23:0] v$OP2_6913_out0;
wire  [23:0] v$OP2_6914_out0;
wire  [23:0] v$OP2_6915_out0;
wire  [23:0] v$OP2_6916_out0;
wire  [23:0] v$OP2_6917_out0;
wire  [23:0] v$OP2_6918_out0;
wire  [23:0] v$OP2_6919_out0;
wire  [23:0] v$OP2_6920_out0;
wire  [23:0] v$OP2_6921_out0;
wire  [23:0] v$OP2_6922_out0;
wire  [23:0] v$OP2_6923_out0;
wire  [23:0] v$OP2_6924_out0;
wire  [23:0] v$OP2_6925_out0;
wire  [23:0] v$OP2_6926_out0;
wire  [23:0] v$OP2_6927_out0;
wire  [23:0] v$OP2_6928_out0;
wire  [23:0] v$OP2_6929_out0;
wire  [23:0] v$OP2_6930_out0;
wire  [23:0] v$OP2_6931_out0;
wire  [23:0] v$OP2_6932_out0;
wire  [23:0] v$OP2_6933_out0;
wire  [23:0] v$OP2_6934_out0;
wire  [23:0] v$OUT_10234_out0;
wire  [23:0] v$OUT_10235_out0;
wire  [23:0] v$OUT_10236_out0;
wire  [23:0] v$OUT_10237_out0;
wire  [23:0] v$OUT_10238_out0;
wire  [23:0] v$OUT_10251_out0;
wire  [23:0] v$OUT_10252_out0;
wire  [23:0] v$OUT_10253_out0;
wire  [23:0] v$OUT_10254_out0;
wire  [23:0] v$OUT_10255_out0;
wire  [23:0] v$OUT_10256_out0;
wire  [23:0] v$OUT_10257_out0;
wire  [23:0] v$OUT_10258_out0;
wire  [23:0] v$OUT_10259_out0;
wire  [23:0] v$OUT_10260_out0;
wire  [23:0] v$OUT_10261_out0;
wire  [23:0] v$OUT_10262_out0;
wire  [23:0] v$OUT_10263_out0;
wire  [23:0] v$OUT_10264_out0;
wire  [23:0] v$OUT_10265_out0;
wire  [23:0] v$OUT_10266_out0;
wire  [23:0] v$OUT_10267_out0;
wire  [23:0] v$OUT_10268_out0;
wire  [23:0] v$OUT_10269_out0;
wire  [23:0] v$OUT_10270_out0;
wire  [23:0] v$OUT_10283_out0;
wire  [23:0] v$OUT_10284_out0;
wire  [23:0] v$OUT_10285_out0;
wire  [23:0] v$OUT_10286_out0;
wire  [23:0] v$OUT_10287_out0;
wire  [23:0] v$OUT_10288_out0;
wire  [23:0] v$OUT_10289_out0;
wire  [23:0] v$OUT_10290_out0;
wire  [23:0] v$OUT_10291_out0;
wire  [23:0] v$OUT_10292_out0;
wire  [23:0] v$OUT_10293_out0;
wire  [23:0] v$OUT_10294_out0;
wire  [23:0] v$OUT_10295_out0;
wire  [23:0] v$OUT_10296_out0;
wire  [23:0] v$OUT_10297_out0;
wire  [23:0] v$OUT_6726_out0;
wire  [23:0] v$OUT_6727_out0;
wire  [23:0] v$OUT_6728_out0;
wire  [23:0] v$OUT_6729_out0;
wire  [23:0] v$OUT_6730_out0;
wire  [23:0] v$OUT_6731_out0;
wire  [23:0] v$OUT_6732_out0;
wire  [23:0] v$OUT_6733_out0;
wire  [23:0] v$SEL6_3784_out0;
wire  [23:0] v$SEL6_3785_out0;
wire  [23:0] v$SUM$EXEC1_13195_out0;
wire  [23:0] v$SUM$EXEC1_13196_out0;
wire  [23:0] v$SUM$HALF_1659_out0;
wire  [23:0] v$SUM$HALF_1660_out0;
wire  [23:0] v$SUM1_3677_out0;
wire  [23:0] v$SUM1_3678_out0;
wire  [23:0] v$SUM_10459_out0;
wire  [23:0] v$SUM_10460_out0;
wire  [23:0] v$SUM_10461_out0;
wire  [23:0] v$SUM_10462_out0;
wire  [23:0] v$SUM_10463_out0;
wire  [23:0] v$SUM_10464_out0;
wire  [23:0] v$SUM_10465_out0;
wire  [23:0] v$SUM_10466_out0;
wire  [23:0] v$SUM_10467_out0;
wire  [23:0] v$SUM_10468_out0;
wire  [23:0] v$SUM_10469_out0;
wire  [23:0] v$SUM_10470_out0;
wire  [23:0] v$SUM_10471_out0;
wire  [23:0] v$SUM_10472_out0;
wire  [23:0] v$SUM_10473_out0;
wire  [23:0] v$SUM_10474_out0;
wire  [23:0] v$SUM_10475_out0;
wire  [23:0] v$SUM_10476_out0;
wire  [23:0] v$SUM_10477_out0;
wire  [23:0] v$SUM_10478_out0;
wire  [23:0] v$SUM_10479_out0;
wire  [23:0] v$SUM_10480_out0;
wire  [23:0] v$SUM_10481_out0;
wire  [23:0] v$SUM_10482_out0;
wire  [23:0] v$SUM_1056_out0;
wire  [23:0] v$SUM_1057_out0;
wire  [23:0] v$SUM_2161_out0;
wire  [23:0] v$SUM_2162_out0;
wire  [23:0] v$SUM_2163_out0;
wire  [23:0] v$SUM_2164_out0;
wire  [23:0] v$SUM_2165_out0;
wire  [23:0] v$SUM_2166_out0;
wire  [23:0] v$SUM_2167_out0;
wire  [23:0] v$SUM_2168_out0;
wire  [23:0] v$SUM_2169_out0;
wire  [23:0] v$SUM_2170_out0;
wire  [23:0] v$SUM_2171_out0;
wire  [23:0] v$SUM_2172_out0;
wire  [23:0] v$SUM_2173_out0;
wire  [23:0] v$SUM_2174_out0;
wire  [23:0] v$SUM_2175_out0;
wire  [23:0] v$SUM_2176_out0;
wire  [23:0] v$SUM_2177_out0;
wire  [23:0] v$SUM_2178_out0;
wire  [23:0] v$SUM_2179_out0;
wire  [23:0] v$SUM_2180_out0;
wire  [23:0] v$SUM_2181_out0;
wire  [23:0] v$SUM_2182_out0;
wire  [23:0] v$SUM_2183_out0;
wire  [23:0] v$SUM_2184_out0;
wire  [23:0] v$SUM_396_out0;
wire  [23:0] v$SUM_397_out0;
wire  [23:0] v$XOR$IN_1172_out0;
wire  [23:0] v$XOR$IN_1173_out0;
wire  [23:0] v$XOR1_3645_out0;
wire  [23:0] v$XOR1_3646_out0;
wire  [23:0] v$XOR2_5376_out0;
wire  [23:0] v$XOR2_5377_out0;
wire  [23:0] v$_10645_out0;
wire  [23:0] v$_10646_out0;
wire  [23:0] v$_12560_out0;
wire  [23:0] v$_12561_out0;
wire  [23:0] v$_12755_out0;
wire  [23:0] v$_12756_out0;
wire  [23:0] v$_12757_out0;
wire  [23:0] v$_12758_out0;
wire  [23:0] v$_12759_out0;
wire  [23:0] v$_12760_out0;
wire  [23:0] v$_12761_out0;
wire  [23:0] v$_12762_out0;
wire  [23:0] v$_12763_out0;
wire  [23:0] v$_12764_out0;
wire  [23:0] v$_12765_out0;
wire  [23:0] v$_12766_out0;
wire  [23:0] v$_12767_out0;
wire  [23:0] v$_12768_out0;
wire  [23:0] v$_12769_out0;
wire  [23:0] v$_12770_out0;
wire  [23:0] v$_12771_out0;
wire  [23:0] v$_12772_out0;
wire  [23:0] v$_12773_out0;
wire  [23:0] v$_12774_out0;
wire  [23:0] v$_12775_out0;
wire  [23:0] v$_12776_out0;
wire  [23:0] v$_12777_out0;
wire  [23:0] v$_12778_out0;
wire  [23:0] v$_2920_out0;
wire  [23:0] v$_2921_out0;
wire  [23:0] v$_2922_out0;
wire  [23:0] v$_2923_out0;
wire  [23:0] v$_2924_out0;
wire  [23:0] v$_2937_out0;
wire  [23:0] v$_2938_out0;
wire  [23:0] v$_2939_out0;
wire  [23:0] v$_2940_out0;
wire  [23:0] v$_2941_out0;
wire  [23:0] v$_2942_out0;
wire  [23:0] v$_2943_out0;
wire  [23:0] v$_2944_out0;
wire  [23:0] v$_2945_out0;
wire  [23:0] v$_2946_out0;
wire  [23:0] v$_2947_out0;
wire  [23:0] v$_2948_out0;
wire  [23:0] v$_2949_out0;
wire  [23:0] v$_2950_out0;
wire  [23:0] v$_2951_out0;
wire  [23:0] v$_2952_out0;
wire  [23:0] v$_2953_out0;
wire  [23:0] v$_2954_out0;
wire  [23:0] v$_2955_out0;
wire  [23:0] v$_2956_out0;
wire  [23:0] v$_2969_out0;
wire  [23:0] v$_2970_out0;
wire  [23:0] v$_2971_out0;
wire  [23:0] v$_2972_out0;
wire  [23:0] v$_2973_out0;
wire  [23:0] v$_2974_out0;
wire  [23:0] v$_2975_out0;
wire  [23:0] v$_2976_out0;
wire  [23:0] v$_2977_out0;
wire  [23:0] v$_2978_out0;
wire  [23:0] v$_2979_out0;
wire  [23:0] v$_2980_out0;
wire  [23:0] v$_2981_out0;
wire  [23:0] v$_2982_out0;
wire  [23:0] v$_2983_out0;
wire  [23:0] v$_5001_out0;
wire  [23:0] v$_5002_out0;
wire  [23:0] v$_5153_out0;
wire  [23:0] v$_5154_out0;
wire  [23:0] v$_6227_out0;
wire  [23:0] v$_6228_out0;
wire  [23:0] v$_6229_out0;
wire  [23:0] v$_6230_out0;
wire  [23:0] v$_6231_out0;
wire  [23:0] v$_6244_out0;
wire  [23:0] v$_6245_out0;
wire  [23:0] v$_6246_out0;
wire  [23:0] v$_6247_out0;
wire  [23:0] v$_6248_out0;
wire  [23:0] v$_6249_out0;
wire  [23:0] v$_6250_out0;
wire  [23:0] v$_6251_out0;
wire  [23:0] v$_6252_out0;
wire  [23:0] v$_6253_out0;
wire  [23:0] v$_6254_out0;
wire  [23:0] v$_6255_out0;
wire  [23:0] v$_6256_out0;
wire  [23:0] v$_6257_out0;
wire  [23:0] v$_6258_out0;
wire  [23:0] v$_6259_out0;
wire  [23:0] v$_6260_out0;
wire  [23:0] v$_6261_out0;
wire  [23:0] v$_6262_out0;
wire  [23:0] v$_6263_out0;
wire  [23:0] v$_6276_out0;
wire  [23:0] v$_6277_out0;
wire  [23:0] v$_6278_out0;
wire  [23:0] v$_6279_out0;
wire  [23:0] v$_6280_out0;
wire  [23:0] v$_6281_out0;
wire  [23:0] v$_6282_out0;
wire  [23:0] v$_6283_out0;
wire  [23:0] v$_6284_out0;
wire  [23:0] v$_6285_out0;
wire  [23:0] v$_6286_out0;
wire  [23:0] v$_6287_out0;
wire  [23:0] v$_6288_out0;
wire  [23:0] v$_6289_out0;
wire  [23:0] v$_6290_out0;
wire  [23:0] v$_6744_out0;
wire  [23:0] v$_6745_out0;
wire  [23:0] v$_7269_out0;
wire  [23:0] v$_7270_out0;
wire  [23:0] v$_735_out0;
wire  [23:0] v$_736_out0;
wire  [23:0] v$_9480_out0;
wire  [23:0] v$_9481_out0;
wire  [23:0] v$_9986_out0;
wire  [23:0] v$_9987_out0;
wire  [24:0] v$_12837_out0;
wire  [24:0] v$_12838_out0;
wire  [24:0] v$_6994_out0;
wire  [24:0] v$_6995_out0;
wire  [25:0] v$_3302_out0;
wire  [25:0] v$_3303_out0;
wire  [25:0] v$_7574_out0;
wire  [25:0] v$_7575_out0;
wire  [26:0] v$_5159_out0;
wire  [26:0] v$_5160_out0;
wire  [26:0] v$_9388_out0;
wire  [26:0] v$_9389_out0;
wire  [27:0] v$_2847_out0;
wire  [27:0] v$_2848_out0;
wire  [27:0] v$_6656_out0;
wire  [27:0] v$_6657_out0;
wire  [27:0] v$_6742_out0;
wire  [27:0] v$_6743_out0;
wire  [28:0] v$_10424_out0;
wire  [28:0] v$_10425_out0;
wire  [28:0] v$_11466_out0;
wire  [28:0] v$_11467_out0;
wire  [29:0] v$_1113_out0;
wire  [29:0] v$_1114_out0;
wire  [29:0] v$_12212_out0;
wire  [29:0] v$_12213_out0;
wire  [2:0] v$9_9550_out0;
wire  [2:0] v$9_9551_out0;
wire  [2:0] v$ALU$OP_11875_out0;
wire  [2:0] v$ALU$OP_11876_out0;
wire  [2:0] v$C10_9110_out0;
wire  [2:0] v$C10_9111_out0;
wire  [2:0] v$C1_11890_out0;
wire  [2:0] v$C1_11891_out0;
wire  [2:0] v$C2_8899_out0;
wire  [2:0] v$C2_8900_out0;
wire  [2:0] v$C4_4630_out0;
wire  [2:0] v$C4_4631_out0;
wire  [2:0] v$IR1$OP_3762_out0;
wire  [2:0] v$IR1$OP_3763_out0;
wire  [2:0] v$IR2$OP_11080_out0;
wire  [2:0] v$IR2$OP_11081_out0;
wire  [2:0] v$IR2$OP_12789_out0;
wire  [2:0] v$IR2$OP_12790_out0;
wire  [2:0] v$MODE_6360_out0;
wire  [2:0] v$MODE_6361_out0;
wire  [2:0] v$MODE_821_out0;
wire  [2:0] v$MODE_822_out0;
wire  [2:0] v$MUX1_10052_out0;
wire  [2:0] v$MUX1_10053_out0;
wire  [2:0] v$MUX1_10054_out0;
wire  [2:0] v$MUX1_10055_out0;
wire  [2:0] v$MUX1_10056_out0;
wire  [2:0] v$MUX1_10057_out0;
wire  [2:0] v$Mode_7235_out0;
wire  [2:0] v$Mode_7236_out0;
wire  [2:0] v$Mode_8796_out0;
wire  [2:0] v$Mode_8797_out0;
wire  [2:0] v$NUPPER_12173_out0;
wire  [2:0] v$NUPPER_12174_out0;
wire  [2:0] v$NUPPER_12175_out0;
wire  [2:0] v$NUPPER_12176_out0;
wire  [2:0] v$OPCODE_5408_out0;
wire  [2:0] v$OPCODE_5409_out0;
wire  [2:0] v$OP_1032_out0;
wire  [2:0] v$OP_1033_out0;
wire  [2:0] v$OP_12461_out0;
wire  [2:0] v$OP_12462_out0;
wire  [2:0] v$SEL26_3242_out0;
wire  [2:0] v$SEL26_3243_out0;
wire  [2:0] v$SEL26_3244_out0;
wire  [2:0] v$SEL26_3245_out0;
wire  [2:0] v$Y_5296_out0;
wire  [2:0] v$Y_5297_out0;
wire  [2:0] v$Y_5298_out0;
wire  [2:0] v$Y_5299_out0;
wire  [2:0] v$Y_5300_out0;
wire  [2:0] v$Y_5301_out0;
wire  [2:0] v$_11744_out0;
wire  [2:0] v$_11745_out0;
wire  [2:0] v$_13197_out0;
wire  [2:0] v$_13198_out0;
wire  [2:0] v$_3288_out0;
wire  [2:0] v$_3289_out0;
wire  [2:0] v$_3390_out0;
wire  [2:0] v$_3391_out0;
wire  [2:0] v$_3712_out0;
wire  [2:0] v$_3713_out0;
wire  [2:0] v$_3714_out0;
wire  [2:0] v$_3715_out0;
wire  [2:0] v$_3716_out0;
wire  [2:0] v$_3717_out0;
wire  [2:0] v$_5609_out0;
wire  [2:0] v$_5610_out0;
wire  [2:0] v$_5652_out0;
wire  [2:0] v$_5653_out0;
wire  [2:0] v$_5654_out0;
wire  [2:0] v$_5655_out0;
wire  [2:0] v$_5656_out0;
wire  [2:0] v$_5657_out0;
wire  [30:0] v$C4_5740_out0;
wire  [30:0] v$C4_5742_out0;
wire  [30:0] v$MUX12_10443_out0;
wire  [30:0] v$MUX12_10444_out0;
wire  [30:0] v$MUX2_9188_out0;
wire  [30:0] v$MUX2_9190_out0;
wire  [30:0] v$MUX6_12238_out0;
wire  [30:0] v$MUX6_12239_out0;
wire  [30:0] v$SINGLE$MERGE_7895_out0;
wire  [30:0] v$SINGLE$MERGE_7896_out0;
wire  [30:0] v$_10647_out0;
wire  [30:0] v$_10648_out0;
wire  [30:0] v$_11065_out0;
wire  [30:0] v$_11067_out0;
wire  [30:0] v$_4780_out0;
wire  [30:0] v$_4781_out0;
wire  [30:0] v$_52_out0;
wire  [30:0] v$_53_out0;
wire  [30:0] v$_5743_out0;
wire  [30:0] v$_5744_out0;
wire  [30:0] v$_7631_out0;
wire  [30:0] v$_7632_out0;
wire  [30:0] v$_8292_out0;
wire  [30:0] v$_8293_out0;
wire  [31:0] v$A$32$BIT$MUL_2491_out0;
wire  [31:0] v$A$32$BIT$MUL_2492_out0;
wire  [31:0] v$A$32$BIT_13121_out0;
wire  [31:0] v$A$32$BIT_13122_out0;
wire  [31:0] v$A$32BIT_1751_out0;
wire  [31:0] v$A$32BIT_1752_out0;
wire  [31:0] v$A$FPU$ADDER$32$BIT_11102_out0;
wire  [31:0] v$A$FPU$ADDER$32$BIT_11103_out0;
wire  [31:0] v$A_9335_out0;
wire  [31:0] v$A_9337_out0;
wire  [31:0] v$A_9339_out0;
wire  [31:0] v$A_9341_out0;
wire  [31:0] v$B$32$BIT$FPU$ADDER_6765_out0;
wire  [31:0] v$B$32$BIT$FPU$ADDER_6766_out0;
wire  [31:0] v$B$32$BIT_1046_out0;
wire  [31:0] v$B$32$BIT_1047_out0;
wire  [31:0] v$B$32$MUL_8842_out0;
wire  [31:0] v$B$32$MUL_8843_out0;
wire  [31:0] v$B$32BIT_13139_out0;
wire  [31:0] v$B$32BIT_13140_out0;
wire  [31:0] v$B_3231_out0;
wire  [31:0] v$B_3233_out0;
wire  [31:0] v$B_3235_out0;
wire  [31:0] v$B_3237_out0;
wire  [31:0] v$C1_10547_out0;
wire  [31:0] v$C1_10548_out0;
wire  [31:0] v$C1_3968_out0;
wire  [31:0] v$C1_3974_out0;
wire  [31:0] v$C1_4000_out0;
wire  [31:0] v$C1_4006_out0;
wire  [31:0] v$C2_101_out0;
wire  [31:0] v$C2_107_out0;
wire  [31:0] v$C2_133_out0;
wire  [31:0] v$C2_139_out0;
wire  [31:0] v$C4_9419_out0;
wire  [31:0] v$C4_9420_out0;
wire  [31:0] v$C5_2811_out0;
wire  [31:0] v$C5_2812_out0;
wire  [31:0] v$FPU$ADDER$OUT_2726_out0;
wire  [31:0] v$FPU$ADDER$OUT_2727_out0;
wire  [31:0] v$FPU$MULTIPLIER$OUT_7195_out0;
wire  [31:0] v$FPU$MULTIPLIER$OUT_7196_out0;
wire  [31:0] v$HALF$PRECISION$32$BIT_10149_out0;
wire  [31:0] v$HALF$PRECISION$32$BIT_10150_out0;
wire  [31:0] v$HALF$PRECISION_6871_out0;
wire  [31:0] v$HALF$PRECISION_6872_out0;
wire  [31:0] v$MUX12_11834_out0;
wire  [31:0] v$MUX12_11835_out0;
wire  [31:0] v$MUX1_9125_out0;
wire  [31:0] v$MUX1_9126_out0;
wire  [31:0] v$MUX2_11385_out0;
wire  [31:0] v$MUX2_11386_out0;
wire  [31:0] v$MUX3_6217_out0;
wire  [31:0] v$MUX3_6218_out0;
wire  [31:0] v$MUX4_519_out0;
wire  [31:0] v$MUX4_520_out0;
wire  [31:0] v$MUX7_3262_out0;
wire  [31:0] v$MUX7_3263_out0;
wire  [31:0] v$OUT1_12605_out0;
wire  [31:0] v$OUT1_12606_out0;
wire  [31:0] v$OUT_2054_out0;
wire  [31:0] v$OUT_2055_out0;
wire  [31:0] v$OUT_8120_out0;
wire  [31:0] v$OUT_8122_out0;
wire  [31:0] v$SEL1_10686_out0;
wire  [31:0] v$SEL1_10692_out0;
wire  [31:0] v$SEL1_10718_out0;
wire  [31:0] v$SEL1_10724_out0;
wire  [31:0] v$SEL1_5942_out0;
wire  [31:0] v$SEL1_5948_out0;
wire  [31:0] v$SEL1_5974_out0;
wire  [31:0] v$SEL1_5980_out0;
wire  [31:0] v$SINGLE$PRECISION_5416_out0;
wire  [31:0] v$SINGLE$PRECISION_5417_out0;
wire  [31:0] v$_1024_out0;
wire  [31:0] v$_1025_out0;
wire  [31:0] v$_11044_out0;
wire  [31:0] v$_11045_out0;
wire  [31:0] v$_11279_out0;
wire  [31:0] v$_11280_out0;
wire  [31:0] v$_11586_out0;
wire  [31:0] v$_11587_out0;
wire  [31:0] v$_11836_out0;
wire  [31:0] v$_11837_out0;
wire  [31:0] v$_12090_out0;
wire  [31:0] v$_12091_out0;
wire  [31:0] v$_12980_out0;
wire  [31:0] v$_12981_out0;
wire  [31:0] v$_13104_out0;
wire  [31:0] v$_13106_out0;
wire  [31:0] v$_3734_out0;
wire  [31:0] v$_3735_out0;
wire  [31:0] v$_8159_out0;
wire  [31:0] v$_8160_out0;
wire  [32:0] v$_6479_out0;
wire  [32:0] v$_6480_out0;
wire  [32:0] v$_8624_out0;
wire  [32:0] v$_8625_out0;
wire  [33:0] v$_11078_out0;
wire  [33:0] v$_11079_out0;
wire  [33:0] v$_11582_out0;
wire  [33:0] v$_11583_out0;
wire  [34:0] v$_1003_out0;
wire  [34:0] v$_1004_out0;
wire  [34:0] v$_11454_out0;
wire  [34:0] v$_11455_out0;
wire  [35:0] v$MULTIPLIER$TO$SAVE_11792_out0;
wire  [35:0] v$MULTIPLIER$TO$SAVE_11793_out0;
wire  [35:0] v$SAVED_10674_out0;
wire  [35:0] v$SAVED_10675_out0;
wire  [35:0] v$_809_out0;
wire  [35:0] v$_810_out0;
wire  [35:0] v$_8889_out0;
wire  [35:0] v$_8890_out0;
wire  [39:0] v$SEL1_10684_out0;
wire  [39:0] v$SEL1_10690_out0;
wire  [39:0] v$SEL1_10716_out0;
wire  [39:0] v$SEL1_10722_out0;
wire  [39:0] v$SEL1_5940_out0;
wire  [39:0] v$SEL1_5946_out0;
wire  [39:0] v$SEL1_5972_out0;
wire  [39:0] v$SEL1_5978_out0;
wire  [3:0] v$3_8971_out0;
wire  [3:0] v$3_8972_out0;
wire  [3:0] v$9_9707_out0;
wire  [3:0] v$9_9708_out0;
wire  [3:0] v$ADDRMSB_10339_out0;
wire  [3:0] v$ADDRMSB_10340_out0;
wire  [3:0] v$A_7352_out0;
wire  [3:0] v$A_7353_out0;
wire  [3:0] v$A_7354_out0;
wire  [3:0] v$A_7356_out0;
wire  [3:0] v$A_7357_out0;
wire  [3:0] v$A_7358_out0;
wire  [3:0] v$A_7360_out0;
wire  [3:0] v$A_7361_out0;
wire  [3:0] v$A_7364_out0;
wire  [3:0] v$A_7365_out0;
wire  [3:0] v$A_7368_out0;
wire  [3:0] v$A_7369_out0;
wire  [3:0] v$A_7370_out0;
wire  [3:0] v$A_7372_out0;
wire  [3:0] v$A_7373_out0;
wire  [3:0] v$A_7374_out0;
wire  [3:0] v$A_7376_out0;
wire  [3:0] v$A_7377_out0;
wire  [3:0] v$A_7380_out0;
wire  [3:0] v$A_7381_out0;
wire  [3:0] v$B_2417_out0;
wire  [3:0] v$B_2418_out0;
wire  [3:0] v$B_5789_out0;
wire  [3:0] v$B_5790_out0;
wire  [3:0] v$B_8806_out0;
wire  [3:0] v$B_8807_out0;
wire  [3:0] v$B_9809_out0;
wire  [3:0] v$B_9810_out0;
wire  [3:0] v$B_9811_out0;
wire  [3:0] v$B_9813_out0;
wire  [3:0] v$B_9814_out0;
wire  [3:0] v$B_9815_out0;
wire  [3:0] v$B_9817_out0;
wire  [3:0] v$B_9818_out0;
wire  [3:0] v$B_9821_out0;
wire  [3:0] v$B_9822_out0;
wire  [3:0] v$B_9825_out0;
wire  [3:0] v$B_9826_out0;
wire  [3:0] v$B_9827_out0;
wire  [3:0] v$B_9829_out0;
wire  [3:0] v$B_9830_out0;
wire  [3:0] v$B_9831_out0;
wire  [3:0] v$B_9833_out0;
wire  [3:0] v$B_9834_out0;
wire  [3:0] v$B_9837_out0;
wire  [3:0] v$B_9838_out0;
wire  [3:0] v$B_9992_out0;
wire  [3:0] v$B_9993_out0;
wire  [3:0] v$C0_190_out0;
wire  [3:0] v$C0_191_out0;
wire  [3:0] v$C12_1981_out0;
wire  [3:0] v$C12_1982_out0;
wire  [3:0] v$C1_3657_out0;
wire  [3:0] v$C1_3658_out0;
wire  [3:0] v$C1_3966_out0;
wire  [3:0] v$C1_3973_out0;
wire  [3:0] v$C1_3979_out0;
wire  [3:0] v$C1_3983_out0;
wire  [3:0] v$C1_3988_out0;
wire  [3:0] v$C1_3993_out0;
wire  [3:0] v$C1_3998_out0;
wire  [3:0] v$C1_4005_out0;
wire  [3:0] v$C1_4011_out0;
wire  [3:0] v$C1_4015_out0;
wire  [3:0] v$C1_4020_out0;
wire  [3:0] v$C1_4025_out0;
wire  [3:0] v$C1_5480_out0;
wire  [3:0] v$C1_5484_out0;
wire  [3:0] v$C1_8474_out0;
wire  [3:0] v$C1_8475_out0;
wire  [3:0] v$C2_106_out0;
wire  [3:0] v$C2_112_out0;
wire  [3:0] v$C2_116_out0;
wire  [3:0] v$C2_121_out0;
wire  [3:0] v$C2_126_out0;
wire  [3:0] v$C2_131_out0;
wire  [3:0] v$C2_138_out0;
wire  [3:0] v$C2_144_out0;
wire  [3:0] v$C2_148_out0;
wire  [3:0] v$C2_153_out0;
wire  [3:0] v$C2_158_out0;
wire  [3:0] v$C2_99_out0;
wire  [3:0] v$C4_7090_out0;
wire  [3:0] v$C4_7091_out0;
wire  [3:0] v$C8_4879_out0;
wire  [3:0] v$C8_4880_out0;
wire  [3:0] v$C8_5798_out0;
wire  [3:0] v$C8_5799_out0;
wire  [3:0] v$IN_10358_out0;
wire  [3:0] v$IN_10359_out0;
wire  [3:0] v$IN_10360_out0;
wire  [3:0] v$IN_10361_out0;
wire  [3:0] v$IN_10362_out0;
wire  [3:0] v$IN_10363_out0;
wire  [3:0] v$IN_10364_out0;
wire  [3:0] v$IN_10365_out0;
wire  [3:0] v$IN_10366_out0;
wire  [3:0] v$IN_10367_out0;
wire  [3:0] v$IN_10368_out0;
wire  [3:0] v$IN_10369_out0;
wire  [3:0] v$IN_10370_out0;
wire  [3:0] v$IN_10371_out0;
wire  [3:0] v$IN_10372_out0;
wire  [3:0] v$IN_10373_out0;
wire  [3:0] v$IN_10374_out0;
wire  [3:0] v$IN_10375_out0;
wire  [3:0] v$IN_10376_out0;
wire  [3:0] v$IN_10377_out0;
wire  [3:0] v$IN_10378_out0;
wire  [3:0] v$IN_10379_out0;
wire  [3:0] v$IN_10380_out0;
wire  [3:0] v$IN_10381_out0;
wire  [3:0] v$IN_10382_out0;
wire  [3:0] v$IN_10383_out0;
wire  [3:0] v$IN_10384_out0;
wire  [3:0] v$IN_10385_out0;
wire  [3:0] v$IN_10386_out0;
wire  [3:0] v$IN_10387_out0;
wire  [3:0] v$IN_10388_out0;
wire  [3:0] v$IN_10389_out0;
wire  [3:0] v$IN_10390_out0;
wire  [3:0] v$IN_10391_out0;
wire  [3:0] v$IN_10392_out0;
wire  [3:0] v$IN_10393_out0;
wire  [3:0] v$IN_10394_out0;
wire  [3:0] v$IN_10395_out0;
wire  [3:0] v$IN_10396_out0;
wire  [3:0] v$IN_10397_out0;
wire  [3:0] v$IN_10398_out0;
wire  [3:0] v$IN_10399_out0;
wire  [3:0] v$IN_10400_out0;
wire  [3:0] v$IN_10401_out0;
wire  [3:0] v$IN_10402_out0;
wire  [3:0] v$IN_10403_out0;
wire  [3:0] v$IN_10404_out0;
wire  [3:0] v$IN_10405_out0;
wire  [3:0] v$IN_10406_out0;
wire  [3:0] v$IN_10407_out0;
wire  [3:0] v$IN_10408_out0;
wire  [3:0] v$IN_10409_out0;
wire  [3:0] v$IN_10410_out0;
wire  [3:0] v$IN_10411_out0;
wire  [3:0] v$IN_10412_out0;
wire  [3:0] v$IN_10413_out0;
wire  [3:0] v$IN_10414_out0;
wire  [3:0] v$IN_10415_out0;
wire  [3:0] v$IN_10416_out0;
wire  [3:0] v$IN_10417_out0;
wire  [3:0] v$IR1$FULL$OP$CODE_12104_out0;
wire  [3:0] v$IR1$FULL$OP$CODE_12105_out0;
wire  [3:0] v$IR1$N_11003_out0;
wire  [3:0] v$IR1$N_11004_out0;
wire  [3:0] v$IR1$OPCODE_1671_out0;
wire  [3:0] v$IR1$OPCODE_1672_out0;
wire  [3:0] v$IR1$OPCODE_6530_out0;
wire  [3:0] v$IR1$OPCODE_6531_out0;
wire  [3:0] v$IR2$FULL$OP$CODE_7620_out0;
wire  [3:0] v$IR2$FULL$OP$CODE_7621_out0;
wire  [3:0] v$IR2$N_1745_out0;
wire  [3:0] v$IR2$N_1746_out0;
wire  [3:0] v$IR2$OPCODE_1482_out0;
wire  [3:0] v$IR2$OPCODE_1483_out0;
wire  [3:0] v$LSBS_10623_out0;
wire  [3:0] v$LSBS_10624_out0;
wire  [3:0] v$MUX3_12264_out0;
wire  [3:0] v$MUX3_12265_out0;
wire  [3:0] v$MUX3_12266_out0;
wire  [3:0] v$MUX3_12267_out0;
wire  [3:0] v$MUX3_12268_out0;
wire  [3:0] v$MUX3_12269_out0;
wire  [3:0] v$MUX3_12270_out0;
wire  [3:0] v$MUX3_12271_out0;
wire  [3:0] v$MUX3_12272_out0;
wire  [3:0] v$MUX3_12273_out0;
wire  [3:0] v$MUX3_12274_out0;
wire  [3:0] v$MUX3_12275_out0;
wire  [3:0] v$MUX4_1642_out0;
wire  [3:0] v$MUX4_1643_out0;
wire  [3:0] v$MUX4_1644_out0;
wire  [3:0] v$MUX4_1646_out0;
wire  [3:0] v$MUX4_1647_out0;
wire  [3:0] v$MUX4_1648_out0;
wire  [3:0] v$MUX4_1650_out0;
wire  [3:0] v$MUX4_1651_out0;
wire  [3:0] v$MUX4_1652_out0;
wire  [3:0] v$MUX4_1654_out0;
wire  [3:0] v$MUX4_1655_out0;
wire  [3:0] v$MUX4_1656_out0;
wire  [3:0] v$MUX5_2765_out0;
wire  [3:0] v$MUX5_2766_out0;
wire  [3:0] v$MUX5_2767_out0;
wire  [3:0] v$MUX5_2769_out0;
wire  [3:0] v$MUX5_2770_out0;
wire  [3:0] v$MUX5_2771_out0;
wire  [3:0] v$MUX5_2773_out0;
wire  [3:0] v$MUX5_2774_out0;
wire  [3:0] v$MUX5_2775_out0;
wire  [3:0] v$MUX5_2777_out0;
wire  [3:0] v$MUX5_2778_out0;
wire  [3:0] v$MUX5_2779_out0;
wire  [3:0] v$MUX5_9877_out0;
wire  [3:0] v$MUX5_9878_out0;
wire  [3:0] v$MUX6_1605_out0;
wire  [3:0] v$MUX6_1606_out0;
wire  [3:0] v$OPCODE_12815_out0;
wire  [3:0] v$OPCODE_12816_out0;
wire  [3:0] v$OP_10131_out0;
wire  [3:0] v$OP_10132_out0;
wire  [3:0] v$OP_12599_out0;
wire  [3:0] v$OP_12600_out0;
wire  [3:0] v$OP_2405_out0;
wire  [3:0] v$OP_2406_out0;
wire  [3:0] v$OP_3431_out0;
wire  [3:0] v$OP_3432_out0;
wire  [3:0] v$OP_7246_out0;
wire  [3:0] v$OP_7247_out0;
wire  [3:0] v$OUT_6200_out0;
wire  [3:0] v$OUT_6201_out0;
wire  [3:0] v$OUT_6202_out0;
wire  [3:0] v$OUT_6204_out0;
wire  [3:0] v$OUT_6205_out0;
wire  [3:0] v$OUT_6206_out0;
wire  [3:0] v$OUT_6208_out0;
wire  [3:0] v$OUT_6209_out0;
wire  [3:0] v$OUT_6210_out0;
wire  [3:0] v$OUT_6212_out0;
wire  [3:0] v$OUT_6213_out0;
wire  [3:0] v$OUT_6214_out0;
wire  [3:0] v$QP_13189_out0;
wire  [3:0] v$QP_13190_out0;
wire  [3:0] v$Q_4167_out0;
wire  [3:0] v$Q_4168_out0;
wire  [3:0] v$Q_8619_out0;
wire  [3:0] v$Q_8620_out0;
wire  [3:0] v$RXFSMQP_6740_out0;
wire  [3:0] v$RXFSMQP_6741_out0;
wire  [3:0] v$RXFSMQ_7116_out0;
wire  [3:0] v$RXFSMQ_7117_out0;
wire  [3:0] v$SEL12_8456_out0;
wire  [3:0] v$SEL12_8457_out0;
wire  [3:0] v$SEL1_11535_out0;
wire  [3:0] v$SEL1_11536_out0;
wire  [3:0] v$SEL1_11537_out0;
wire  [3:0] v$SEL1_11538_out0;
wire  [3:0] v$SEL1_11539_out0;
wire  [3:0] v$SEL1_11540_out0;
wire  [3:0] v$SEL1_11747_out0;
wire  [3:0] v$SEL1_11748_out0;
wire  [3:0] v$SEL1_11749_out0;
wire  [3:0] v$SEL1_11751_out0;
wire  [3:0] v$SEL1_11752_out0;
wire  [3:0] v$SEL1_11753_out0;
wire  [3:0] v$SEL1_11755_out0;
wire  [3:0] v$SEL1_11756_out0;
wire  [3:0] v$SEL1_11757_out0;
wire  [3:0] v$SEL1_11759_out0;
wire  [3:0] v$SEL1_11760_out0;
wire  [3:0] v$SEL1_11761_out0;
wire  [3:0] v$SEL1_12970_out0;
wire  [3:0] v$SEL1_12971_out0;
wire  [3:0] v$SEL1_6041_out0;
wire  [3:0] v$SEL1_6042_out0;
wire  [3:0] v$SEL1_6851_out0;
wire  [3:0] v$SEL1_6852_out0;
wire  [3:0] v$SEL1_6853_out0;
wire  [3:0] v$SEL1_6854_out0;
wire  [3:0] v$SEL1_6855_out0;
wire  [3:0] v$SEL1_6856_out0;
wire  [3:0] v$SEL1_6857_out0;
wire  [3:0] v$SEL1_6858_out0;
wire  [3:0] v$SEL2_12242_out0;
wire  [3:0] v$SEL2_12243_out0;
wire  [3:0] v$SEL2_12244_out0;
wire  [3:0] v$SEL2_12245_out0;
wire  [3:0] v$SEL2_12246_out0;
wire  [3:0] v$SEL2_12247_out0;
wire  [3:0] v$SEL2_12248_out0;
wire  [3:0] v$SEL2_12249_out0;
wire  [3:0] v$SEL2_1361_out0;
wire  [3:0] v$SEL2_1362_out0;
wire  [3:0] v$SEL2_1785_out0;
wire  [3:0] v$SEL2_1786_out0;
wire  [3:0] v$SEL2_1787_out0;
wire  [3:0] v$SEL2_1788_out0;
wire  [3:0] v$SEL2_1789_out0;
wire  [3:0] v$SEL2_1790_out0;
wire  [3:0] v$SEL2_9369_out0;
wire  [3:0] v$SEL2_9370_out0;
wire  [3:0] v$SEL2_9371_out0;
wire  [3:0] v$SEL2_9373_out0;
wire  [3:0] v$SEL2_9374_out0;
wire  [3:0] v$SEL2_9375_out0;
wire  [3:0] v$SEL2_9377_out0;
wire  [3:0] v$SEL2_9378_out0;
wire  [3:0] v$SEL2_9379_out0;
wire  [3:0] v$SEL2_9381_out0;
wire  [3:0] v$SEL2_9382_out0;
wire  [3:0] v$SEL2_9383_out0;
wire  [3:0] v$SEL3_11722_out0;
wire  [3:0] v$SEL3_11723_out0;
wire  [3:0] v$SEL3_13253_out0;
wire  [3:0] v$SEL3_13254_out0;
wire  [3:0] v$SEL3_13255_out0;
wire  [3:0] v$SEL3_13256_out0;
wire  [3:0] v$SEL3_4958_out0;
wire  [3:0] v$SEL3_4959_out0;
wire  [3:0] v$SEL3_4960_out0;
wire  [3:0] v$SEL3_4962_out0;
wire  [3:0] v$SEL3_4963_out0;
wire  [3:0] v$SEL3_4964_out0;
wire  [3:0] v$SEL3_4966_out0;
wire  [3:0] v$SEL3_4967_out0;
wire  [3:0] v$SEL3_4968_out0;
wire  [3:0] v$SEL3_4970_out0;
wire  [3:0] v$SEL3_4971_out0;
wire  [3:0] v$SEL3_4972_out0;
wire  [3:0] v$SEL3_6295_out0;
wire  [3:0] v$SEL3_6296_out0;
wire  [3:0] v$SEL3_6297_out0;
wire  [3:0] v$SEL3_6298_out0;
wire  [3:0] v$SEL3_6299_out0;
wire  [3:0] v$SEL3_6300_out0;
wire  [3:0] v$SEL3_6301_out0;
wire  [3:0] v$SEL3_6302_out0;
wire  [3:0] v$SEL4_12149_out0;
wire  [3:0] v$SEL4_12150_out0;
wire  [3:0] v$SEL4_12151_out0;
wire  [3:0] v$SEL4_12152_out0;
wire  [3:0] v$SEL4_12153_out0;
wire  [3:0] v$SEL4_12154_out0;
wire  [3:0] v$SEL4_12155_out0;
wire  [3:0] v$SEL4_12156_out0;
wire  [3:0] v$SEL4_2058_out0;
wire  [3:0] v$SEL4_2059_out0;
wire  [3:0] v$SEL4_2060_out0;
wire  [3:0] v$SEL4_2061_out0;
wire  [3:0] v$SEL4_2062_out0;
wire  [3:0] v$SEL4_2063_out0;
wire  [3:0] v$SEL4_2064_out0;
wire  [3:0] v$SEL4_2065_out0;
wire  [3:0] v$SEL4_2066_out0;
wire  [3:0] v$SEL4_2067_out0;
wire  [3:0] v$SEL4_2068_out0;
wire  [3:0] v$SEL4_2069_out0;
wire  [3:0] v$SEL4_6540_out0;
wire  [3:0] v$SEL4_6541_out0;
wire  [3:0] v$SEL4_6542_out0;
wire  [3:0] v$SEL4_6543_out0;
wire  [3:0] v$TXFSMQP_6013_out0;
wire  [3:0] v$TXFSMQP_6014_out0;
wire  [3:0] v$TXFSMQ_4224_out0;
wire  [3:0] v$TXFSMQ_4225_out0;
wire  [3:0] v$USELESS_10774_out0;
wire  [3:0] v$_1009_out0;
wire  [3:0] v$_1010_out0;
wire  [3:0] v$_11221_out0;
wire  [3:0] v$_11222_out0;
wire  [3:0] v$_11296_out0;
wire  [3:0] v$_11297_out0;
wire  [3:0] v$_11935_out0;
wire  [3:0] v$_11936_out0;
wire  [3:0] v$_12218_out0;
wire  [3:0] v$_12219_out0;
wire  [3:0] v$_1279_out0;
wire  [3:0] v$_1279_out1;
wire  [3:0] v$_1280_out0;
wire  [3:0] v$_1280_out1;
wire  [3:0] v$_12972_out0;
wire  [3:0] v$_12973_out0;
wire  [3:0] v$_13131_out0;
wire  [3:0] v$_13131_out1;
wire  [3:0] v$_13132_out0;
wire  [3:0] v$_13132_out1;
wire  [3:0] v$_13249_out0;
wire  [3:0] v$_13250_out0;
wire  [3:0] v$_1673_out0;
wire  [3:0] v$_1673_out1;
wire  [3:0] v$_1674_out0;
wire  [3:0] v$_1674_out1;
wire  [3:0] v$_223_out0;
wire  [3:0] v$_224_out0;
wire  [3:0] v$_2419_out0;
wire  [3:0] v$_2420_out0;
wire  [3:0] v$_2507_out0;
wire  [3:0] v$_2508_out0;
wire  [3:0] v$_256_out0;
wire  [3:0] v$_257_out0;
wire  [3:0] v$_2700_out0;
wire  [3:0] v$_2701_out0;
wire  [3:0] v$_2702_out0;
wire  [3:0] v$_2703_out0;
wire  [3:0] v$_2704_out0;
wire  [3:0] v$_2705_out0;
wire  [3:0] v$_2706_out0;
wire  [3:0] v$_2707_out0;
wire  [3:0] v$_2708_out0;
wire  [3:0] v$_2709_out0;
wire  [3:0] v$_2710_out0;
wire  [3:0] v$_2711_out0;
wire  [3:0] v$_2854_out0;
wire  [3:0] v$_2855_out0;
wire  [3:0] v$_3462_out0;
wire  [3:0] v$_3463_out0;
wire  [3:0] v$_3464_out0;
wire  [3:0] v$_3466_out0;
wire  [3:0] v$_3467_out0;
wire  [3:0] v$_3468_out0;
wire  [3:0] v$_3470_out0;
wire  [3:0] v$_3471_out0;
wire  [3:0] v$_3472_out0;
wire  [3:0] v$_3474_out0;
wire  [3:0] v$_3475_out0;
wire  [3:0] v$_3476_out0;
wire  [3:0] v$_3609_out0;
wire  [3:0] v$_3610_out0;
wire  [3:0] v$_3718_out0;
wire  [3:0] v$_3719_out0;
wire  [3:0] v$_3760_out0;
wire  [3:0] v$_3761_out0;
wire  [3:0] v$_392_out0;
wire  [3:0] v$_393_out0;
wire  [3:0] v$_4355_out0;
wire  [3:0] v$_4356_out0;
wire  [3:0] v$_4458_out0;
wire  [3:0] v$_4458_out1;
wire  [3:0] v$_4459_out0;
wire  [3:0] v$_4459_out1;
wire  [3:0] v$_4751_out0;
wire  [3:0] v$_4752_out0;
wire  [3:0] v$_4782_out0;
wire  [3:0] v$_4783_out0;
wire  [3:0] v$_4875_out0;
wire  [3:0] v$_4977_out0;
wire  [3:0] v$_4978_out0;
wire  [3:0] v$_500_out0;
wire  [3:0] v$_501_out0;
wire  [3:0] v$_5102_out0;
wire  [3:0] v$_5103_out0;
wire  [3:0] v$_5706_out0;
wire  [3:0] v$_5706_out1;
wire  [3:0] v$_5707_out0;
wire  [3:0] v$_5707_out1;
wire  [3:0] v$_5874_out0;
wire  [3:0] v$_5874_out1;
wire  [3:0] v$_5875_out0;
wire  [3:0] v$_5875_out1;
wire  [3:0] v$_5930_out0;
wire  [3:0] v$_5931_out0;
wire  [3:0] v$_6022_out0;
wire  [3:0] v$_6023_out0;
wire  [3:0] v$_6024_out0;
wire  [3:0] v$_6026_out0;
wire  [3:0] v$_6027_out0;
wire  [3:0] v$_6028_out0;
wire  [3:0] v$_6030_out0;
wire  [3:0] v$_6031_out0;
wire  [3:0] v$_6032_out0;
wire  [3:0] v$_6034_out0;
wire  [3:0] v$_6035_out0;
wire  [3:0] v$_6036_out0;
wire  [3:0] v$_6148_out0;
wire  [3:0] v$_6149_out0;
wire  [3:0] v$_6150_out0;
wire  [3:0] v$_6152_out0;
wire  [3:0] v$_6153_out0;
wire  [3:0] v$_6154_out0;
wire  [3:0] v$_6156_out0;
wire  [3:0] v$_6157_out0;
wire  [3:0] v$_6158_out0;
wire  [3:0] v$_6160_out0;
wire  [3:0] v$_6161_out0;
wire  [3:0] v$_6162_out0;
wire  [3:0] v$_6183_out0;
wire  [3:0] v$_6184_out0;
wire  [3:0] v$_6427_out0;
wire  [3:0] v$_6428_out0;
wire  [3:0] v$_6821_out0;
wire  [3:0] v$_6822_out0;
wire  [3:0] v$_8504_out0;
wire  [3:0] v$_8504_out1;
wire  [3:0] v$_8505_out0;
wire  [3:0] v$_8505_out1;
wire  [3:0] v$_8506_out0;
wire  [3:0] v$_8506_out1;
wire  [3:0] v$_8507_out0;
wire  [3:0] v$_8507_out1;
wire  [3:0] v$_8508_out0;
wire  [3:0] v$_8508_out1;
wire  [3:0] v$_8509_out0;
wire  [3:0] v$_8509_out1;
wire  [3:0] v$_8510_out0;
wire  [3:0] v$_8510_out1;
wire  [3:0] v$_8511_out0;
wire  [3:0] v$_8511_out1;
wire  [3:0] v$_8512_out0;
wire  [3:0] v$_8512_out1;
wire  [3:0] v$_8513_out0;
wire  [3:0] v$_8513_out1;
wire  [3:0] v$_8514_out0;
wire  [3:0] v$_8514_out1;
wire  [3:0] v$_8515_out0;
wire  [3:0] v$_8515_out1;
wire  [3:0] v$_8546_out0;
wire  [3:0] v$_8547_out0;
wire  [3:0] v$_8636_out0;
wire  [3:0] v$_8637_out0;
wire  [3:0] v$_8853_out0;
wire  [3:0] v$_8856_out0;
wire  [3:0] v$_9417_out1;
wire  [3:0] v$_9418_out1;
wire  [43:0] v$AROM1_11322_out0;
wire  [43:0] v$AROM1_11323_out0;
wire  [43:0] v$SEL1_10688_out0;
wire  [43:0] v$SEL1_10694_out0;
wire  [43:0] v$SEL1_10720_out0;
wire  [43:0] v$SEL1_10726_out0;
wire  [43:0] v$SEL1_5944_out0;
wire  [43:0] v$SEL1_5950_out0;
wire  [43:0] v$SEL1_5976_out0;
wire  [43:0] v$SEL1_5982_out0;
wire  [45:0] v$SEL1_10685_out0;
wire  [45:0] v$SEL1_10691_out0;
wire  [45:0] v$SEL1_10717_out0;
wire  [45:0] v$SEL1_10723_out0;
wire  [45:0] v$SEL1_5941_out0;
wire  [45:0] v$SEL1_5947_out0;
wire  [45:0] v$SEL1_5973_out0;
wire  [45:0] v$SEL1_5979_out0;
wire  [46:0] v$SEL1_10687_out0;
wire  [46:0] v$SEL1_10693_out0;
wire  [46:0] v$SEL1_10719_out0;
wire  [46:0] v$SEL1_10725_out0;
wire  [46:0] v$SEL1_5943_out0;
wire  [46:0] v$SEL1_5949_out0;
wire  [46:0] v$SEL1_5975_out0;
wire  [46:0] v$SEL1_5981_out0;
wire  [47:0] v$IN_10873_out0;
wire  [47:0] v$IN_10874_out0;
wire  [47:0] v$IN_10879_out0;
wire  [47:0] v$IN_10880_out0;
wire  [47:0] v$IN_12982_out0;
wire  [47:0] v$IN_12983_out0;
wire  [47:0] v$IN_12984_out0;
wire  [47:0] v$IN_12985_out0;
wire  [47:0] v$IN_2567_out0;
wire  [47:0] v$IN_2568_out0;
wire  [47:0] v$IN_2569_out0;
wire  [47:0] v$IN_2570_out0;
wire  [47:0] v$IN_2571_out0;
wire  [47:0] v$IN_2572_out0;
wire  [47:0] v$IN_2577_out0;
wire  [47:0] v$IN_2578_out0;
wire  [47:0] v$IN_2579_out0;
wire  [47:0] v$IN_2580_out0;
wire  [47:0] v$IN_2581_out0;
wire  [47:0] v$IN_2582_out0;
wire  [47:0] v$IN_2880_out0;
wire  [47:0] v$IN_2881_out0;
wire  [47:0] v$IN_2882_out0;
wire  [47:0] v$IN_2883_out0;
wire  [47:0] v$IN_3413_out0;
wire  [47:0] v$IN_3414_out0;
wire  [47:0] v$IN_3423_out0;
wire  [47:0] v$IN_3424_out0;
wire  [47:0] v$IN_3526_out0;
wire  [47:0] v$IN_3527_out0;
wire  [47:0] v$IN_3528_out0;
wire  [47:0] v$IN_3529_out0;
wire  [47:0] v$IN_3530_out0;
wire  [47:0] v$IN_3531_out0;
wire  [47:0] v$IN_3532_out0;
wire  [47:0] v$IN_3533_out0;
wire  [47:0] v$IN_3534_out0;
wire  [47:0] v$IN_3535_out0;
wire  [47:0] v$IN_3536_out0;
wire  [47:0] v$IN_3537_out0;
wire  [47:0] v$IN_3558_out0;
wire  [47:0] v$IN_3559_out0;
wire  [47:0] v$IN_3560_out0;
wire  [47:0] v$IN_3561_out0;
wire  [47:0] v$IN_3562_out0;
wire  [47:0] v$IN_3563_out0;
wire  [47:0] v$IN_3564_out0;
wire  [47:0] v$IN_3565_out0;
wire  [47:0] v$IN_3566_out0;
wire  [47:0] v$IN_3567_out0;
wire  [47:0] v$IN_3568_out0;
wire  [47:0] v$IN_3569_out0;
wire  [47:0] v$IN_5768_out0;
wire  [47:0] v$IN_5769_out0;
wire  [47:0] v$IN_5770_out0;
wire  [47:0] v$IN_5771_out0;
wire  [47:0] v$IN_7304_out0;
wire  [47:0] v$IN_7305_out0;
wire  [47:0] v$IN_7306_out0;
wire  [47:0] v$IN_7307_out0;
wire  [47:0] v$IN_7482_out0;
wire  [47:0] v$IN_7483_out0;
wire  [47:0] v$IN_7484_out0;
wire  [47:0] v$IN_7485_out0;
wire  [47:0] v$IN_7583_out0;
wire  [47:0] v$IN_7584_out0;
wire  [47:0] v$IN_7589_out0;
wire  [47:0] v$IN_7590_out0;
wire  [47:0] v$IN_9131_out0;
wire  [47:0] v$IN_9135_out0;
wire  [47:0] v$IN_9139_out0;
wire  [47:0] v$IN_9143_out0;
wire  [47:0] v$MULTIPLIER$OUT_3807_out0;
wire  [47:0] v$MULTIPLIER$OUT_3808_out0;
wire  [47:0] v$MULTIPLIER$OUT_6372_out0;
wire  [47:0] v$MULTIPLIER$OUT_6373_out0;
wire  [47:0] v$MUX1_1288_out0;
wire  [47:0] v$MUX1_1289_out0;
wire  [47:0] v$MUX1_1290_out0;
wire  [47:0] v$MUX1_1291_out0;
wire  [47:0] v$MUX1_1292_out0;
wire  [47:0] v$MUX1_1293_out0;
wire  [47:0] v$MUX1_1294_out0;
wire  [47:0] v$MUX1_1295_out0;
wire  [47:0] v$MUX1_1296_out0;
wire  [47:0] v$MUX1_1297_out0;
wire  [47:0] v$MUX1_1298_out0;
wire  [47:0] v$MUX1_1299_out0;
wire  [47:0] v$MUX1_1320_out0;
wire  [47:0] v$MUX1_1321_out0;
wire  [47:0] v$MUX1_1322_out0;
wire  [47:0] v$MUX1_1323_out0;
wire  [47:0] v$MUX1_1324_out0;
wire  [47:0] v$MUX1_1325_out0;
wire  [47:0] v$MUX1_1326_out0;
wire  [47:0] v$MUX1_1327_out0;
wire  [47:0] v$MUX1_1328_out0;
wire  [47:0] v$MUX1_1329_out0;
wire  [47:0] v$MUX1_1330_out0;
wire  [47:0] v$MUX1_1331_out0;
wire  [47:0] v$MUX2_10556_out0;
wire  [47:0] v$MUX2_10557_out0;
wire  [47:0] v$MUX2_10562_out0;
wire  [47:0] v$MUX2_10563_out0;
wire  [47:0] v$MUX2_13218_out0;
wire  [47:0] v$MUX2_13219_out0;
wire  [47:0] v$MUX2_13220_out0;
wire  [47:0] v$MUX2_13221_out0;
wire  [47:0] v$MUX2_13222_out0;
wire  [47:0] v$MUX2_13223_out0;
wire  [47:0] v$MUX2_13228_out0;
wire  [47:0] v$MUX2_13229_out0;
wire  [47:0] v$MUX2_13230_out0;
wire  [47:0] v$MUX2_13231_out0;
wire  [47:0] v$MUX2_13232_out0;
wire  [47:0] v$MUX2_13233_out0;
wire  [47:0] v$MUX2_1394_out0;
wire  [47:0] v$MUX2_1395_out0;
wire  [47:0] v$MUX2_1400_out0;
wire  [47:0] v$MUX2_1401_out0;
wire  [47:0] v$MUX2_1407_out0;
wire  [47:0] v$MUX2_1408_out0;
wire  [47:0] v$MUX2_1417_out0;
wire  [47:0] v$MUX2_1418_out0;
wire  [47:0] v$OUT_10239_out0;
wire  [47:0] v$OUT_10240_out0;
wire  [47:0] v$OUT_10241_out0;
wire  [47:0] v$OUT_10242_out0;
wire  [47:0] v$OUT_10243_out0;
wire  [47:0] v$OUT_10244_out0;
wire  [47:0] v$OUT_10245_out0;
wire  [47:0] v$OUT_10246_out0;
wire  [47:0] v$OUT_10247_out0;
wire  [47:0] v$OUT_10248_out0;
wire  [47:0] v$OUT_10249_out0;
wire  [47:0] v$OUT_10250_out0;
wire  [47:0] v$OUT_10271_out0;
wire  [47:0] v$OUT_10272_out0;
wire  [47:0] v$OUT_10273_out0;
wire  [47:0] v$OUT_10274_out0;
wire  [47:0] v$OUT_10275_out0;
wire  [47:0] v$OUT_10276_out0;
wire  [47:0] v$OUT_10277_out0;
wire  [47:0] v$OUT_10278_out0;
wire  [47:0] v$OUT_10279_out0;
wire  [47:0] v$OUT_10280_out0;
wire  [47:0] v$OUT_10281_out0;
wire  [47:0] v$OUT_10282_out0;
wire  [47:0] v$OUT_3306_out0;
wire  [47:0] v$OUT_3307_out0;
wire  [47:0] v$OUT_3308_out0;
wire  [47:0] v$OUT_3309_out0;
wire  [47:0] v$OUT_5704_out0;
wire  [47:0] v$OUT_5705_out0;
wire  [47:0] v$_1441_out0;
wire  [47:0] v$_1442_out0;
wire  [47:0] v$_2925_out0;
wire  [47:0] v$_2926_out0;
wire  [47:0] v$_2927_out0;
wire  [47:0] v$_2928_out0;
wire  [47:0] v$_2929_out0;
wire  [47:0] v$_2930_out0;
wire  [47:0] v$_2931_out0;
wire  [47:0] v$_2932_out0;
wire  [47:0] v$_2933_out0;
wire  [47:0] v$_2934_out0;
wire  [47:0] v$_2935_out0;
wire  [47:0] v$_2936_out0;
wire  [47:0] v$_2957_out0;
wire  [47:0] v$_2958_out0;
wire  [47:0] v$_2959_out0;
wire  [47:0] v$_2960_out0;
wire  [47:0] v$_2961_out0;
wire  [47:0] v$_2962_out0;
wire  [47:0] v$_2963_out0;
wire  [47:0] v$_2964_out0;
wire  [47:0] v$_2965_out0;
wire  [47:0] v$_2966_out0;
wire  [47:0] v$_2967_out0;
wire  [47:0] v$_2968_out0;
wire  [47:0] v$_6232_out0;
wire  [47:0] v$_6233_out0;
wire  [47:0] v$_6234_out0;
wire  [47:0] v$_6235_out0;
wire  [47:0] v$_6236_out0;
wire  [47:0] v$_6237_out0;
wire  [47:0] v$_6238_out0;
wire  [47:0] v$_6239_out0;
wire  [47:0] v$_6240_out0;
wire  [47:0] v$_6241_out0;
wire  [47:0] v$_6242_out0;
wire  [47:0] v$_6243_out0;
wire  [47:0] v$_6264_out0;
wire  [47:0] v$_6265_out0;
wire  [47:0] v$_6266_out0;
wire  [47:0] v$_6267_out0;
wire  [47:0] v$_6268_out0;
wire  [47:0] v$_6269_out0;
wire  [47:0] v$_6270_out0;
wire  [47:0] v$_6271_out0;
wire  [47:0] v$_6272_out0;
wire  [47:0] v$_6273_out0;
wire  [47:0] v$_6274_out0;
wire  [47:0] v$_6275_out0;
wire  [4:0] v$A$EXP_236_out0;
wire  [4:0] v$A$EXP_238_out0;
wire  [4:0] v$A$EXP_240_out0;
wire  [4:0] v$A$EXP_242_out0;
wire  [4:0] v$A1_1564_out0;
wire  [4:0] v$A1_1566_out0;
wire  [4:0] v$A1_3809_out0;
wire  [4:0] v$A1_3811_out0;
wire  [4:0] v$A1_3813_out0;
wire  [4:0] v$A1_3815_out0;
wire  [4:0] v$A1_5275_out0;
wire  [4:0] v$A1_5276_out0;
wire  [4:0] v$A1_7602_out0;
wire  [4:0] v$A1_7603_out0;
wire  [4:0] v$A2_6750_out0;
wire  [4:0] v$A2_6752_out0;
wire  [4:0] v$A_7350_out0;
wire  [4:0] v$A_7362_out0;
wire  [4:0] v$A_7366_out0;
wire  [4:0] v$A_7378_out0;
wire  [4:0] v$B$EXP_11734_out0;
wire  [4:0] v$B$EXP_11736_out0;
wire  [4:0] v$B$EXP_11738_out0;
wire  [4:0] v$B$EXP_11740_out0;
wire  [4:0] v$B_9807_out0;
wire  [4:0] v$B_9819_out0;
wire  [4:0] v$B_9823_out0;
wire  [4:0] v$B_9835_out0;
wire  [4:0] v$C1_10982_out0;
wire  [4:0] v$C1_10983_out0;
wire  [4:0] v$C1_3957_out0;
wire  [4:0] v$C1_3959_out0;
wire  [4:0] v$C1_5006_out0;
wire  [4:0] v$C1_5007_out0;
wire  [4:0] v$C1_9147_out0;
wire  [4:0] v$C1_9149_out0;
wire  [4:0] v$C1_9151_out0;
wire  [4:0] v$C1_9153_out0;
wire  [4:0] v$DIFF_6326_out0;
wire  [4:0] v$DIFF_6328_out0;
wire  [4:0] v$DIFF_6330_out0;
wire  [4:0] v$DIFF_6332_out0;
wire  [4:0] v$EXPONENT_11194_out0;
wire  [4:0] v$EXPONENT_11195_out0;
wire  [4:0] v$EXPONENT_11500_out0;
wire  [4:0] v$EXPONENT_11501_out0;
wire  [4:0] v$EXPONENT_12831_out0;
wire  [4:0] v$EXPONENT_12832_out0;
wire  [4:0] v$HALF$PRECISION$EXPONENT$DENORM_4143_out0;
wire  [4:0] v$HALF$PRECISION$EXPONENT$DENORM_4144_out0;
wire  [4:0] v$HALF$PRECISION$EXPONENT_10032_out0;
wire  [4:0] v$HALF$PRECISION$EXPONENT_10033_out0;
wire  [4:0] v$HALF$PRECISION$EXPONENT_4401_out0;
wire  [4:0] v$HALF$PRECISION$EXPONENT_4402_out0;
wire  [4:0] v$HALF$PRECISSION$ADDITION$IN_447_out0;
wire  [4:0] v$HALF$PRECISSION$ADDITION$IN_448_out0;
wire  [4:0] v$K_253_out0;
wire  [4:0] v$K_254_out0;
wire  [4:0] v$LARGER$EXP_6839_out0;
wire  [4:0] v$LARGER$EXP_6841_out0;
wire  [4:0] v$MUX1_10603_out0;
wire  [4:0] v$MUX1_10604_out0;
wire  [4:0] v$MUX1_12699_out0;
wire  [4:0] v$MUX1_12701_out0;
wire  [4:0] v$MUX1_12703_out0;
wire  [4:0] v$MUX1_12705_out0;
wire  [4:0] v$MUX2_9114_out0;
wire  [4:0] v$MUX2_9115_out0;
wire  [4:0] v$MUX3_2097_out0;
wire  [4:0] v$MUX3_2099_out0;
wire  [4:0] v$MUX3_2101_out0;
wire  [4:0] v$MUX3_2103_out0;
wire  [4:0] v$NORMALIZATION$SHIFT_1000_out0;
wire  [4:0] v$NORMALIZATION$SHIFT_3052_out0;
wire  [4:0] v$NORMALIZATION$SHIFT_3053_out0;
wire  [4:0] v$NORMALIZATION$SHIFT_999_out0;
wire  [4:0] v$N_11398_out0;
wire  [4:0] v$N_11399_out0;
wire  [4:0] v$N_11400_out0;
wire  [4:0] v$N_11401_out0;
wire  [4:0] v$OUT_164_out0;
wire  [4:0] v$OUT_165_out0;
wire  [4:0] v$OUT_4211_out0;
wire  [4:0] v$OUT_4212_out0;
wire  [4:0] v$OUT_6175_out0;
wire  [4:0] v$OUT_6176_out0;
wire  [4:0] v$SEL10_1771_out0;
wire  [4:0] v$SEL10_1772_out0;
wire  [4:0] v$SEL14_6339_out0;
wire  [4:0] v$SEL14_6340_out0;
wire  [4:0] v$SEL18_12974_out0;
wire  [4:0] v$SEL18_12975_out0;
wire  [4:0] v$SEL1_5086_out0;
wire  [4:0] v$SEL1_5088_out0;
wire  [4:0] v$SEL1_5090_out0;
wire  [4:0] v$SEL1_5092_out0;
wire  [4:0] v$SEL1_6461_out0;
wire  [4:0] v$SEL1_6462_out0;
wire  [4:0] v$SEL25_9020_out0;
wire  [4:0] v$SEL25_9021_out0;
wire  [4:0] v$SEL25_9022_out0;
wire  [4:0] v$SEL25_9023_out0;
wire  [4:0] v$SEL2_4733_out0;
wire  [4:0] v$SEL2_4735_out0;
wire  [4:0] v$SEL2_4737_out0;
wire  [4:0] v$SEL2_4739_out0;
wire  [4:0] v$SEL9_2481_out0;
wire  [4:0] v$SEL9_2482_out0;
wire  [4:0] v$SMALLER$EXP_1707_out0;
wire  [4:0] v$SMALLER$EXP_1709_out0;
wire  [4:0] v$XOR1_5128_out0;
wire  [4:0] v$XOR1_5130_out0;
wire  [4:0] v$XOR1_5132_out0;
wire  [4:0] v$XOR1_5134_out0;
wire  [4:0] v$XOR1_7199_out0;
wire  [4:0] v$XOR1_7200_out0;
wire  [4:0] v$_1577_out0;
wire  [4:0] v$_1578_out0;
wire  [4:0] v$_2021_out0;
wire  [4:0] v$_2022_out0;
wire  [4:0] v$_4353_out0;
wire  [4:0] v$_4354_out0;
wire  [4:0] v$_4871_out0;
wire  [4:0] v$_4872_out0;
wire  [4:0] v$_555_out0;
wire  [4:0] v$_556_out0;
wire  [5:0] v$A1_2728_out0;
wire  [5:0] v$A1_2729_out0;
wire  [5:0] v$A2_10173_out0;
wire  [5:0] v$A2_10174_out0;
wire  [5:0] v$ADDRESS_9958_out0;
wire  [5:0] v$ADDRESS_9959_out0;
wire  [5:0] v$AMOUNT$OF$SHIFT_6455_out0;
wire  [5:0] v$AMOUNT$OF$SHIFT_6456_out0;
wire  [5:0] v$AMOUNT$OF$SHIFT_6457_out0;
wire  [5:0] v$AMOUNT$OF$SHIFT_6458_out0;
wire  [5:0] v$C2_11174_out0;
wire  [5:0] v$C2_11175_out0;
wire  [5:0] v$C3_8772_out0;
wire  [5:0] v$C3_8773_out0;
wire  [5:0] v$C6_5555_out0;
wire  [5:0] v$C6_5556_out0;
wire  [5:0] v$MUX1_6647_out0;
wire  [5:0] v$MUX1_6648_out0;
wire  [5:0] v$MUX4_1641_out0;
wire  [5:0] v$MUX4_1645_out0;
wire  [5:0] v$MUX4_1649_out0;
wire  [5:0] v$MUX4_1653_out0;
wire  [5:0] v$MUX5_2764_out0;
wire  [5:0] v$MUX5_2768_out0;
wire  [5:0] v$MUX5_2772_out0;
wire  [5:0] v$MUX5_2776_out0;
wire  [5:0] v$OUT_6199_out0;
wire  [5:0] v$OUT_6203_out0;
wire  [5:0] v$OUT_6207_out0;
wire  [5:0] v$OUT_6211_out0;
wire  [5:0] v$_3461_out0;
wire  [5:0] v$_3465_out0;
wire  [5:0] v$_3469_out0;
wire  [5:0] v$_3473_out0;
wire  [5:0] v$_6021_out0;
wire  [5:0] v$_6025_out0;
wire  [5:0] v$_6029_out0;
wire  [5:0] v$_6033_out0;
wire  [5:0] v$_6147_out0;
wire  [5:0] v$_6151_out0;
wire  [5:0] v$_6155_out0;
wire  [5:0] v$_6159_out0;
wire  [7:0] v$8LSB_5144_out0;
wire  [7:0] v$8LSB_5145_out0;
wire  [7:0] v$A$EXP_237_out0;
wire  [7:0] v$A$EXP_239_out0;
wire  [7:0] v$A$EXP_241_out0;
wire  [7:0] v$A$EXP_243_out0;
wire  [7:0] v$A1_11001_out0;
wire  [7:0] v$A1_11002_out0;
wire  [7:0] v$A1_1565_out0;
wire  [7:0] v$A1_1567_out0;
wire  [7:0] v$A1_362_out0;
wire  [7:0] v$A1_363_out0;
wire  [7:0] v$A1_3810_out0;
wire  [7:0] v$A1_3812_out0;
wire  [7:0] v$A1_3814_out0;
wire  [7:0] v$A1_3816_out0;
wire  [7:0] v$A2_6751_out0;
wire  [7:0] v$A2_6753_out0;
wire  [7:0] v$A_7351_out0;
wire  [7:0] v$A_7355_out0;
wire  [7:0] v$A_7359_out0;
wire  [7:0] v$A_7363_out0;
wire  [7:0] v$A_7367_out0;
wire  [7:0] v$A_7371_out0;
wire  [7:0] v$A_7375_out0;
wire  [7:0] v$A_7379_out0;
wire  [7:0] v$B$EXP_11735_out0;
wire  [7:0] v$B$EXP_11737_out0;
wire  [7:0] v$B$EXP_11739_out0;
wire  [7:0] v$B$EXP_11741_out0;
wire  [7:0] v$B_9808_out0;
wire  [7:0] v$B_9812_out0;
wire  [7:0] v$B_9816_out0;
wire  [7:0] v$B_9820_out0;
wire  [7:0] v$B_9824_out0;
wire  [7:0] v$B_9828_out0;
wire  [7:0] v$B_9832_out0;
wire  [7:0] v$B_9836_out0;
wire  [7:0] v$C1_10160_out0;
wire  [7:0] v$C1_10161_out0;
wire  [7:0] v$C1_3958_out0;
wire  [7:0] v$C1_3960_out0;
wire  [7:0] v$C1_3964_out0;
wire  [7:0] v$C1_3969_out0;
wire  [7:0] v$C1_3975_out0;
wire  [7:0] v$C1_3981_out0;
wire  [7:0] v$C1_3986_out0;
wire  [7:0] v$C1_3991_out0;
wire  [7:0] v$C1_3996_out0;
wire  [7:0] v$C1_4001_out0;
wire  [7:0] v$C1_4007_out0;
wire  [7:0] v$C1_4013_out0;
wire  [7:0] v$C1_4018_out0;
wire  [7:0] v$C1_4023_out0;
wire  [7:0] v$C1_5481_out0;
wire  [7:0] v$C1_5485_out0;
wire  [7:0] v$C1_767_out0;
wire  [7:0] v$C1_768_out0;
wire  [7:0] v$C1_9014_out0;
wire  [7:0] v$C1_9015_out0;
wire  [7:0] v$C1_9148_out0;
wire  [7:0] v$C1_9150_out0;
wire  [7:0] v$C1_9152_out0;
wire  [7:0] v$C1_9154_out0;
wire  [7:0] v$C1_9390_out0;
wire  [7:0] v$C1_9391_out0;
wire  [7:0] v$C2_102_out0;
wire  [7:0] v$C2_108_out0;
wire  [7:0] v$C2_114_out0;
wire  [7:0] v$C2_119_out0;
wire  [7:0] v$C2_124_out0;
wire  [7:0] v$C2_129_out0;
wire  [7:0] v$C2_134_out0;
wire  [7:0] v$C2_140_out0;
wire  [7:0] v$C2_146_out0;
wire  [7:0] v$C2_151_out0;
wire  [7:0] v$C2_156_out0;
wire  [7:0] v$C2_97_out0;
wire  [7:0] v$DIFF$VIEW$MANTISA$ADDER_8380_out0;
wire  [7:0] v$DIFF$VIEW$MANTISA$ADDER_8381_out0;
wire  [7:0] v$DIFF_11134_out0;
wire  [7:0] v$DIFF_11135_out0;
wire  [7:0] v$DIFF_12292_out0;
wire  [7:0] v$DIFF_12293_out0;
wire  [7:0] v$DIFF_12294_out0;
wire  [7:0] v$DIFF_12295_out0;
wire  [7:0] v$DIFF_1587_out0;
wire  [7:0] v$DIFF_1588_out0;
wire  [7:0] v$DIFF_244_out0;
wire  [7:0] v$DIFF_245_out0;
wire  [7:0] v$DIFF_6327_out0;
wire  [7:0] v$DIFF_6329_out0;
wire  [7:0] v$DIFF_6331_out0;
wire  [7:0] v$DIFF_6333_out0;
wire  [7:0] v$DIFF_8303_out0;
wire  [7:0] v$DIFF_8304_out0;
wire  [7:0] v$EDGEMODE_1663_out0;
wire  [7:0] v$EDGEMODE_1664_out0;
wire  [7:0] v$END_8367_out0;
wire  [7:0] v$END_8368_out0;
wire  [7:0] v$EXP$DIFF_12503_out0;
wire  [7:0] v$EXP$DIFF_12504_out0;
wire  [7:0] v$EXP$DIFF_8111_out0;
wire  [7:0] v$EXP$DIFF_8112_out0;
wire  [7:0] v$EXP$DIFF_9312_out0;
wire  [7:0] v$EXP$DIFF_9313_out0;
wire  [7:0] v$EXP$DIFF_9717_out0;
wire  [7:0] v$EXP$DIFF_9718_out0;
wire  [7:0] v$EXPONENT_583_out0;
wire  [7:0] v$EXPONENT_584_out0;
wire  [7:0] v$EXPONENT_9232_out0;
wire  [7:0] v$EXPONENT_9233_out0;
wire  [7:0] v$IN_10194_out0;
wire  [7:0] v$IN_10195_out0;
wire  [7:0] v$IN_10196_out0;
wire  [7:0] v$IN_10197_out0;
wire  [7:0] v$IN_10198_out0;
wire  [7:0] v$IN_10199_out0;
wire  [7:0] v$LARGER$EXP_6840_out0;
wire  [7:0] v$LARGER$EXP_6842_out0;
wire  [7:0] v$LSBS_5438_out0;
wire  [7:0] v$LSBS_5439_out0;
wire  [7:0] v$MODEIN_3801_out0;
wire  [7:0] v$MODEIN_3802_out0;
wire  [7:0] v$MODE_12630_out0;
wire  [7:0] v$MODE_12631_out0;
wire  [7:0] v$MODE_44_out0;
wire  [7:0] v$MODE_45_out0;
wire  [7:0] v$MODE_7108_out0;
wire  [7:0] v$MODE_7109_out0;
wire  [7:0] v$MUX13_6905_out0;
wire  [7:0] v$MUX13_6906_out0;
wire  [7:0] v$MUX1_12700_out0;
wire  [7:0] v$MUX1_12702_out0;
wire  [7:0] v$MUX1_12704_out0;
wire  [7:0] v$MUX1_12706_out0;
wire  [7:0] v$MUX2_12550_out0;
wire  [7:0] v$MUX2_12551_out0;
wire  [7:0] v$MUX3_2098_out0;
wire  [7:0] v$MUX3_2100_out0;
wire  [7:0] v$MUX3_2102_out0;
wire  [7:0] v$MUX3_2104_out0;
wire  [7:0] v$MUX5_8784_out0;
wire  [7:0] v$MUX5_8785_out0;
wire  [7:0] v$MUX6_5444_out0;
wire  [7:0] v$MUX6_5445_out0;
wire  [7:0] v$MUX6_9251_out0;
wire  [7:0] v$MUX6_9252_out0;
wire  [7:0] v$NORMALIZATION$SHIFT$WHOLE_4662_out0;
wire  [7:0] v$NORMALIZATION$SHIFT$WHOLE_4663_out0;
wire  [7:0] v$NORMALIZATION$SHIFT_13257_out0;
wire  [7:0] v$NORMALIZATION$SHIFT_13258_out0;
wire  [7:0] v$NORMALIZATION$SHIFT_1957_out0;
wire  [7:0] v$NORMALIZATION$SHIFT_1958_out0;
wire  [7:0] v$NORMALIZATION$SHIFT_459_out0;
wire  [7:0] v$NORMALIZATION$SHIFT_460_out0;
wire  [7:0] v$NORMALIZATION$SHIFT_7068_out0;
wire  [7:0] v$NORMALIZATION$SHIFT_7069_out0;
wire  [7:0] v$N_9462_out0;
wire  [7:0] v$N_9463_out0;
wire  [7:0] v$N_9464_out0;
wire  [7:0] v$N_9465_out0;
wire  [7:0] v$OUT_10129_out0;
wire  [7:0] v$OUT_10130_out0;
wire  [7:0] v$OUT_11281_out0;
wire  [7:0] v$OUT_11282_out0;
wire  [7:0] v$PIN_4634_out0;
wire  [7:0] v$PIN_4635_out0;
wire  [7:0] v$PIN_4636_out0;
wire  [7:0] v$PIN_4637_out0;
wire  [7:0] v$PIN_4638_out0;
wire  [7:0] v$PIN_4639_out0;
wire  [7:0] v$PIN_4640_out0;
wire  [7:0] v$PIN_4641_out0;
wire  [7:0] v$PIN_4642_out0;
wire  [7:0] v$PIN_4643_out0;
wire  [7:0] v$PIN_4644_out0;
wire  [7:0] v$PIN_4645_out0;
wire  [7:0] v$POUT_6903_out0;
wire  [7:0] v$POUT_6904_out0;
wire  [7:0] v$POut_9234_out0;
wire  [7:0] v$POut_9235_out0;
wire  [7:0] v$RXBYTE_13082_out0;
wire  [7:0] v$RXBYTE_13083_out0;
wire  [7:0] v$RXBYTE_6584_out0;
wire  [7:0] v$RXBYTE_6585_out0;
wire  [7:0] v$SEL17_3633_out0;
wire  [7:0] v$SEL17_3634_out0;
wire  [7:0] v$SEL1_10678_out0;
wire  [7:0] v$SEL1_10695_out0;
wire  [7:0] v$SEL1_10700_out0;
wire  [7:0] v$SEL1_10705_out0;
wire  [7:0] v$SEL1_10710_out0;
wire  [7:0] v$SEL1_10727_out0;
wire  [7:0] v$SEL1_10732_out0;
wire  [7:0] v$SEL1_10737_out0;
wire  [7:0] v$SEL1_12232_out0;
wire  [7:0] v$SEL1_12233_out0;
wire  [7:0] v$SEL1_282_out0;
wire  [7:0] v$SEL1_283_out0;
wire  [7:0] v$SEL1_5087_out0;
wire  [7:0] v$SEL1_5089_out0;
wire  [7:0] v$SEL1_5091_out0;
wire  [7:0] v$SEL1_5093_out0;
wire  [7:0] v$SEL1_5590_out0;
wire  [7:0] v$SEL1_5591_out0;
wire  [7:0] v$SEL1_5592_out0;
wire  [7:0] v$SEL1_5593_out0;
wire  [7:0] v$SEL1_5934_out0;
wire  [7:0] v$SEL1_5951_out0;
wire  [7:0] v$SEL1_5956_out0;
wire  [7:0] v$SEL1_5961_out0;
wire  [7:0] v$SEL1_5966_out0;
wire  [7:0] v$SEL1_5983_out0;
wire  [7:0] v$SEL1_5988_out0;
wire  [7:0] v$SEL1_5993_out0;
wire  [7:0] v$SEL2_12179_out0;
wire  [7:0] v$SEL2_12180_out0;
wire  [7:0] v$SEL2_12312_out0;
wire  [7:0] v$SEL2_12313_out0;
wire  [7:0] v$SEL2_12314_out0;
wire  [7:0] v$SEL2_12315_out0;
wire  [7:0] v$SEL2_4734_out0;
wire  [7:0] v$SEL2_4736_out0;
wire  [7:0] v$SEL2_4738_out0;
wire  [7:0] v$SEL2_4740_out0;
wire  [7:0] v$SEL3_12563_out0;
wire  [7:0] v$SEL3_12564_out0;
wire  [7:0] v$SEL3_12613_out0;
wire  [7:0] v$SEL3_12614_out0;
wire  [7:0] v$SEL4_7649_out0;
wire  [7:0] v$SEL4_7650_out0;
wire  [7:0] v$SEL4_7972_out0;
wire  [7:0] v$SEL4_7973_out0;
wire  [7:0] v$SHIFT$AMOUNT_4980_out0;
wire  [7:0] v$SHIFT$AMOUNT_4981_out0;
wire  [7:0] v$SHIFT$AMOUNT_4982_out0;
wire  [7:0] v$SHIFT$AMOUNT_4983_out0;
wire  [7:0] v$SHIFT$AMOUNT_4984_out0;
wire  [7:0] v$SHIFT$AMOUNT_4985_out0;
wire  [7:0] v$SHIFT$AMOUNT_4986_out0;
wire  [7:0] v$SHIFT$AMOUNT_4987_out0;
wire  [7:0] v$SINGLE$EXPONENT_4815_out0;
wire  [7:0] v$SINGLE$EXPONENT_4816_out0;
wire  [7:0] v$SINGLE$PRECISION$EXPONENT_7284_out0;
wire  [7:0] v$SINGLE$PRECISION$EXPONENT_7285_out0;
wire  [7:0] v$SMALLER$EXP_1708_out0;
wire  [7:0] v$SMALLER$EXP_1710_out0;
wire  [7:0] v$STATUS_28_out0;
wire  [7:0] v$STATUS_29_out0;
wire  [7:0] v$STATUS_6055_out0;
wire  [7:0] v$STATUS_6056_out0;
wire  [7:0] v$Status_2499_out0;
wire  [7:0] v$Status_2500_out0;
wire  [7:0] v$XOR1_5129_out0;
wire  [7:0] v$XOR1_5131_out0;
wire  [7:0] v$XOR1_5133_out0;
wire  [7:0] v$XOR1_5135_out0;
wire  [7:0] v$XOR1_9935_out0;
wire  [7:0] v$XOR1_9936_out0;
wire  [7:0] v$_10005_out0;
wire  [7:0] v$_10009_out0;
wire  [7:0] v$_10020_out0;
wire  [7:0] v$_10021_out0;
wire  [7:0] v$_10934_out0;
wire  [7:0] v$_10935_out0;
wire  [7:0] v$_11334_out0;
wire  [7:0] v$_11335_out0;
wire  [7:0] v$_11797_out0;
wire  [7:0] v$_11801_out0;
wire  [7:0] v$_11807_out0;
wire  [7:0] v$_11807_out1;
wire  [7:0] v$_11808_out0;
wire  [7:0] v$_11808_out1;
wire  [7:0] v$_12214_out0;
wire  [7:0] v$_12215_out0;
wire  [7:0] v$_2402_out0;
wire  [7:0] v$_2403_out0;
wire  [7:0] v$_3212_out0;
wire  [7:0] v$_3216_out0;
wire  [7:0] v$_4875_out1;
wire  [7:0] v$_5148_out0;
wire  [7:0] v$_5149_out0;
wire  [7:0] v$_5418_out0;
wire  [7:0] v$_5418_out1;
wire  [7:0] v$_5419_out0;
wire  [7:0] v$_5419_out1;
wire  [7:0] v$_6223_out0;
wire  [7:0] v$_6223_out1;
wire  [7:0] v$_6224_out0;
wire  [7:0] v$_6224_out1;
wire  [7:0] v$_6291_out0;
wire  [7:0] v$_6292_out0;
wire  [7:0] v$_6907_out0;
wire  [7:0] v$_6908_out0;
wire  [7:0] v$_749_out0;
wire  [7:0] v$_749_out1;
wire  [7:0] v$_750_out0;
wire  [7:0] v$_750_out1;
wire  [7:0] v$_8546_out1;
wire  [7:0] v$_8547_out1;
wire  [7:0] v$_863_out0;
wire  [7:0] v$_864_out0;
wire  [7:0] v$_865_out0;
wire  [7:0] v$_865_out1;
wire  [7:0] v$_866_out0;
wire  [7:0] v$_866_out1;
wire  [7:0] v$_8854_out0;
wire  [7:0] v$_8857_out0;
wire  [7:0] v$_9482_out0;
wire  [7:0] v$_9483_out0;
wire  [7:0] v$_9705_out0;
wire  [7:0] v$_9706_out0;
wire  [7:0] v$_9979_out0;
wire  [7:0] v$_9983_out0;
wire  [9:0] v$HALF$PRECISION$MANTISA$DENORM_9885_out0;
wire  [9:0] v$HALF$PRECISION$MANTISA$DENORM_9886_out0;
wire  [9:0] v$SEL10_1921_out0;
wire  [9:0] v$SEL10_1922_out0;
wire  [9:0] v$SEL12_18_out0;
wire  [9:0] v$SEL12_19_out0;
wire  [9:0] v$SEL2_5605_out0;
wire  [9:0] v$SEL2_5607_out0;
wire  [9:0] v$SEL5_5338_out0;
wire  [9:0] v$SEL5_5339_out0;
wire  [9:0] v$SEL7_1973_out0;
wire  [9:0] v$SEL7_1974_out0;
wire  [9:0] v$SEL7_8117_out0;
wire  [9:0] v$SEL7_8118_out0;
wire  [9:0] v$SEL9_6684_out0;
wire  [9:0] v$SEL9_6685_out0;
wire v$1_755_out0;
wire v$1_756_out0;
wire v$2StopBits_2191_out0;
wire v$2StopBits_2192_out0;
wire v$32BIT_11086_out0;
wire v$32BIT_11087_out0;
wire v$32BIT_7201_out0;
wire v$32BIT_7202_out0;
wire v$4_10457_out0;
wire v$4_10458_out0;
wire v$5_8062_out0;
wire v$5_8063_out0;
wire v$6_1094_out0;
wire v$6_1095_out0;
wire v$6_6615_out0;
wire v$6_6616_out0;
wire v$7_10649_out0;
wire v$7_10650_out0;
wire v$8_10817_out0;
wire v$8_10818_out0;
wire v$A$EXP$LARGER_12280_out0;
wire v$A$EXP$LARGER_12281_out0;
wire v$A$EXP$LARGER_12968_out0;
wire v$A$EXP$LARGER_12969_out0;
wire v$A$EXP$LARGER_6437_out0;
wire v$A$EXP$LARGER_6438_out0;
wire v$A$IS$OP1_3397_out0;
wire v$A$IS$OP1_3398_out0;
wire v$A$MANTISA$LARGER_10068_out0;
wire v$A$MANTISA$LARGER_10069_out0;
wire v$A$MANTISA$LARGER_11207_out0;
wire v$A$MANTISA$LARGER_11208_out0;
wire v$A0$COMP$B0_5492_out0;
wire v$A0$COMP$B0_5493_out0;
wire v$A0$COMP$B0_5494_out0;
wire v$A0$COMP$B0_5495_out0;
wire v$A0$COMP$B0_5496_out0;
wire v$A0$COMP$B0_5497_out0;
wire v$A0$COMP$B0_5498_out0;
wire v$A0$COMP$B0_5499_out0;
wire v$A0$COMP$B0_5500_out0;
wire v$A0$COMP$B0_5501_out0;
wire v$A0$COMP$B0_5502_out0;
wire v$A0$COMP$B0_5503_out0;
wire v$A0$COMP$B0_5504_out0;
wire v$A0$COMP$B0_5505_out0;
wire v$A0$COMP$B0_5506_out0;
wire v$A0$COMP$B0_5507_out0;
wire v$A0$COMP$B0_5508_out0;
wire v$A0$COMP$B0_5509_out0;
wire v$A0$COMP$B0_5510_out0;
wire v$A0$COMP$B0_5511_out0;
wire v$A0$COMP$B0_5512_out0;
wire v$A0$COMP$B0_5513_out0;
wire v$A0$COMP$B0_5514_out0;
wire v$A0$COMP$B0_5515_out0;
wire v$A0XNORB0_669_out0;
wire v$A0XNORB0_670_out0;
wire v$A0XNORB0_671_out0;
wire v$A0XNORB0_672_out0;
wire v$A0XNORB0_673_out0;
wire v$A0XNORB0_674_out0;
wire v$A0XNORB0_675_out0;
wire v$A0XNORB0_676_out0;
wire v$A0XNORB0_677_out0;
wire v$A0XNORB0_678_out0;
wire v$A0XNORB0_679_out0;
wire v$A0XNORB0_680_out0;
wire v$A0XNORB0_681_out0;
wire v$A0XNORB0_682_out0;
wire v$A0XNORB0_683_out0;
wire v$A0XNORB0_684_out0;
wire v$A0XNORB0_685_out0;
wire v$A0XNORB0_686_out0;
wire v$A0XNORB0_687_out0;
wire v$A0XNORB0_688_out0;
wire v$A0XNORB0_689_out0;
wire v$A0XNORB0_690_out0;
wire v$A0XNORB0_691_out0;
wire v$A0XNORB0_692_out0;
wire v$A0_905_out0;
wire v$A0_906_out0;
wire v$A0_907_out0;
wire v$A0_908_out0;
wire v$A0_909_out0;
wire v$A0_910_out0;
wire v$A0_911_out0;
wire v$A0_912_out0;
wire v$A0_913_out0;
wire v$A0_914_out0;
wire v$A0_915_out0;
wire v$A0_916_out0;
wire v$A0_917_out0;
wire v$A0_918_out0;
wire v$A0_919_out0;
wire v$A0_920_out0;
wire v$A0_921_out0;
wire v$A0_922_out0;
wire v$A0_923_out0;
wire v$A0_924_out0;
wire v$A0_925_out0;
wire v$A0_926_out0;
wire v$A0_927_out0;
wire v$A0_928_out0;
wire v$A1$COMP$B1_8127_out0;
wire v$A1$COMP$B1_8128_out0;
wire v$A1$COMP$B1_8129_out0;
wire v$A1$COMP$B1_8130_out0;
wire v$A1$COMP$B1_8131_out0;
wire v$A1$COMP$B1_8132_out0;
wire v$A1$COMP$B1_8133_out0;
wire v$A1$COMP$B1_8134_out0;
wire v$A1$COMP$B1_8135_out0;
wire v$A1$COMP$B1_8136_out0;
wire v$A1$COMP$B1_8137_out0;
wire v$A1$COMP$B1_8138_out0;
wire v$A1$COMP$B1_8139_out0;
wire v$A1$COMP$B1_8140_out0;
wire v$A1$COMP$B1_8141_out0;
wire v$A1$COMP$B1_8142_out0;
wire v$A1$COMP$B1_8143_out0;
wire v$A1$COMP$B1_8144_out0;
wire v$A1$COMP$B1_8145_out0;
wire v$A1$COMP$B1_8146_out0;
wire v$A1$COMP$B1_8147_out0;
wire v$A1$COMP$B1_8148_out0;
wire v$A1$COMP$B1_8149_out0;
wire v$A1$COMP$B1_8150_out0;
wire v$A1XNORB1_11225_out0;
wire v$A1XNORB1_11226_out0;
wire v$A1XNORB1_11227_out0;
wire v$A1XNORB1_11228_out0;
wire v$A1XNORB1_11229_out0;
wire v$A1XNORB1_11230_out0;
wire v$A1XNORB1_11231_out0;
wire v$A1XNORB1_11232_out0;
wire v$A1XNORB1_11233_out0;
wire v$A1XNORB1_11234_out0;
wire v$A1XNORB1_11235_out0;
wire v$A1XNORB1_11236_out0;
wire v$A1XNORB1_11237_out0;
wire v$A1XNORB1_11238_out0;
wire v$A1XNORB1_11239_out0;
wire v$A1XNORB1_11240_out0;
wire v$A1XNORB1_11241_out0;
wire v$A1XNORB1_11242_out0;
wire v$A1XNORB1_11243_out0;
wire v$A1XNORB1_11244_out0;
wire v$A1XNORB1_11245_out0;
wire v$A1XNORB1_11246_out0;
wire v$A1XNORB1_11247_out0;
wire v$A1XNORB1_11248_out0;
wire v$A1_10168_out1;
wire v$A1_10169_out1;
wire v$A1_10523_out1;
wire v$A1_10524_out1;
wire v$A1_10525_out1;
wire v$A1_10526_out1;
wire v$A1_10527_out1;
wire v$A1_10528_out1;
wire v$A1_10529_out1;
wire v$A1_10530_out1;
wire v$A1_10531_out1;
wire v$A1_10532_out1;
wire v$A1_10533_out1;
wire v$A1_10534_out1;
wire v$A1_10535_out1;
wire v$A1_10536_out1;
wire v$A1_10537_out1;
wire v$A1_10538_out1;
wire v$A1_10539_out1;
wire v$A1_10540_out1;
wire v$A1_10541_out1;
wire v$A1_10542_out1;
wire v$A1_10543_out1;
wire v$A1_10544_out1;
wire v$A1_10545_out1;
wire v$A1_10546_out1;
wire v$A1_11001_out1;
wire v$A1_11002_out1;
wire v$A1_1564_out1;
wire v$A1_1565_out1;
wire v$A1_1566_out1;
wire v$A1_1567_out1;
wire v$A1_229_out1;
wire v$A1_230_out1;
wire v$A1_2728_out1;
wire v$A1_2729_out1;
wire v$A1_362_out1;
wire v$A1_363_out1;
wire v$A1_3809_out1;
wire v$A1_3810_out1;
wire v$A1_3811_out1;
wire v$A1_3812_out1;
wire v$A1_3813_out1;
wire v$A1_3814_out1;
wire v$A1_3815_out1;
wire v$A1_3816_out1;
wire v$A1_4421_out1;
wire v$A1_4422_out1;
wire v$A1_5275_out1;
wire v$A1_5276_out1;
wire v$A1_6425_out1;
wire v$A1_6426_out1;
wire v$A1_7602_out1;
wire v$A1_7603_out1;
wire v$A1_9247_out1;
wire v$A1_9248_out1;
wire v$A1_9726_out0;
wire v$A1_9727_out0;
wire v$A1_9728_out0;
wire v$A1_9729_out0;
wire v$A1_9730_out0;
wire v$A1_9731_out0;
wire v$A1_9732_out0;
wire v$A1_9733_out0;
wire v$A1_9734_out0;
wire v$A1_9735_out0;
wire v$A1_9736_out0;
wire v$A1_9737_out0;
wire v$A1_9738_out0;
wire v$A1_9739_out0;
wire v$A1_9740_out0;
wire v$A1_9741_out0;
wire v$A1_9742_out0;
wire v$A1_9743_out0;
wire v$A1_9744_out0;
wire v$A1_9745_out0;
wire v$A1_9746_out0;
wire v$A1_9747_out0;
wire v$A1_9748_out0;
wire v$A1_9749_out0;
wire v$A2$COMP$B2_1115_out0;
wire v$A2$COMP$B2_1116_out0;
wire v$A2$COMP$B2_1117_out0;
wire v$A2$COMP$B2_1118_out0;
wire v$A2$COMP$B2_1119_out0;
wire v$A2$COMP$B2_1120_out0;
wire v$A2$COMP$B2_1121_out0;
wire v$A2$COMP$B2_1122_out0;
wire v$A2$COMP$B2_1123_out0;
wire v$A2$COMP$B2_1124_out0;
wire v$A2$COMP$B2_1125_out0;
wire v$A2$COMP$B2_1126_out0;
wire v$A2$COMP$B2_1127_out0;
wire v$A2$COMP$B2_1128_out0;
wire v$A2$COMP$B2_1129_out0;
wire v$A2$COMP$B2_1130_out0;
wire v$A2$COMP$B2_1131_out0;
wire v$A2$COMP$B2_1132_out0;
wire v$A2$COMP$B2_1133_out0;
wire v$A2$COMP$B2_1134_out0;
wire v$A2$COMP$B2_1135_out0;
wire v$A2$COMP$B2_1136_out0;
wire v$A2$COMP$B2_1137_out0;
wire v$A2$COMP$B2_1138_out0;
wire v$A2XNORB2_3125_out0;
wire v$A2XNORB2_3126_out0;
wire v$A2XNORB2_3127_out0;
wire v$A2XNORB2_3128_out0;
wire v$A2XNORB2_3129_out0;
wire v$A2XNORB2_3130_out0;
wire v$A2XNORB2_3131_out0;
wire v$A2XNORB2_3132_out0;
wire v$A2XNORB2_3133_out0;
wire v$A2XNORB2_3134_out0;
wire v$A2XNORB2_3135_out0;
wire v$A2XNORB2_3136_out0;
wire v$A2XNORB2_3137_out0;
wire v$A2XNORB2_3138_out0;
wire v$A2XNORB2_3139_out0;
wire v$A2XNORB2_3140_out0;
wire v$A2XNORB2_3141_out0;
wire v$A2XNORB2_3142_out0;
wire v$A2XNORB2_3143_out0;
wire v$A2XNORB2_3144_out0;
wire v$A2XNORB2_3145_out0;
wire v$A2XNORB2_3146_out0;
wire v$A2XNORB2_3147_out0;
wire v$A2XNORB2_3148_out0;
wire v$A2_10173_out1;
wire v$A2_10174_out1;
wire v$A2_5564_out0;
wire v$A2_5565_out0;
wire v$A2_5566_out0;
wire v$A2_5567_out0;
wire v$A2_5568_out0;
wire v$A2_5569_out0;
wire v$A2_5570_out0;
wire v$A2_5571_out0;
wire v$A2_5572_out0;
wire v$A2_5573_out0;
wire v$A2_5574_out0;
wire v$A2_5575_out0;
wire v$A2_5576_out0;
wire v$A2_5577_out0;
wire v$A2_5578_out0;
wire v$A2_5579_out0;
wire v$A2_5580_out0;
wire v$A2_5581_out0;
wire v$A2_5582_out0;
wire v$A2_5583_out0;
wire v$A2_5584_out0;
wire v$A2_5585_out0;
wire v$A2_5586_out0;
wire v$A2_5587_out0;
wire v$A2_6750_out1;
wire v$A2_6751_out1;
wire v$A2_6752_out1;
wire v$A2_6753_out1;
wire v$A2_8371_out1;
wire v$A2_8372_out1;
wire v$A3$COMP$B3_3338_out0;
wire v$A3$COMP$B3_3339_out0;
wire v$A3$COMP$B3_3340_out0;
wire v$A3$COMP$B3_3341_out0;
wire v$A3$COMP$B3_3342_out0;
wire v$A3$COMP$B3_3343_out0;
wire v$A3$COMP$B3_3344_out0;
wire v$A3$COMP$B3_3345_out0;
wire v$A3$COMP$B3_3346_out0;
wire v$A3$COMP$B3_3347_out0;
wire v$A3$COMP$B3_3348_out0;
wire v$A3$COMP$B3_3349_out0;
wire v$A3$COMP$B3_3350_out0;
wire v$A3$COMP$B3_3351_out0;
wire v$A3$COMP$B3_3352_out0;
wire v$A3$COMP$B3_3353_out0;
wire v$A3$COMP$B3_3354_out0;
wire v$A3$COMP$B3_3355_out0;
wire v$A3$COMP$B3_3356_out0;
wire v$A3$COMP$B3_3357_out0;
wire v$A3$COMP$B3_3358_out0;
wire v$A3$COMP$B3_3359_out0;
wire v$A3$COMP$B3_3360_out0;
wire v$A3$COMP$B3_3361_out0;
wire v$A3XNORB3_10072_out0;
wire v$A3XNORB3_10073_out0;
wire v$A3XNORB3_10074_out0;
wire v$A3XNORB3_10075_out0;
wire v$A3XNORB3_10076_out0;
wire v$A3XNORB3_10077_out0;
wire v$A3XNORB3_10078_out0;
wire v$A3XNORB3_10079_out0;
wire v$A3XNORB3_10080_out0;
wire v$A3XNORB3_10081_out0;
wire v$A3XNORB3_10082_out0;
wire v$A3XNORB3_10083_out0;
wire v$A3XNORB3_10084_out0;
wire v$A3XNORB3_10085_out0;
wire v$A3XNORB3_10086_out0;
wire v$A3XNORB3_10087_out0;
wire v$A3XNORB3_10088_out0;
wire v$A3XNORB3_10089_out0;
wire v$A3XNORB3_10090_out0;
wire v$A3XNORB3_10091_out0;
wire v$A3XNORB3_10092_out0;
wire v$A3XNORB3_10093_out0;
wire v$A3XNORB3_10094_out0;
wire v$A3XNORB3_10095_out0;
wire v$A3_7018_out0;
wire v$A3_7019_out0;
wire v$A3_7020_out0;
wire v$A3_7021_out0;
wire v$A3_7022_out0;
wire v$A3_7023_out0;
wire v$A3_7024_out0;
wire v$A3_7025_out0;
wire v$A3_7026_out0;
wire v$A3_7027_out0;
wire v$A3_7028_out0;
wire v$A3_7029_out0;
wire v$A3_7030_out0;
wire v$A3_7031_out0;
wire v$A3_7032_out0;
wire v$A3_7033_out0;
wire v$A3_7034_out0;
wire v$A3_7035_out0;
wire v$A3_7036_out0;
wire v$A3_7037_out0;
wire v$A3_7038_out0;
wire v$A3_7039_out0;
wire v$A3_7040_out0;
wire v$A3_7041_out0;
wire v$A4$COMP$B4_4997_out0;
wire v$A4$COMP$B4_4998_out0;
wire v$A4$COMP$B4_4999_out0;
wire v$A4$COMP$B4_5000_out0;
wire v$A4XNORB4_597_out0;
wire v$A4XNORB4_598_out0;
wire v$A4XNORB4_599_out0;
wire v$A4XNORB4_600_out0;
wire v$A4_10323_out0;
wire v$A4_10324_out0;
wire v$A4_10325_out0;
wire v$A4_10326_out0;
wire v$AD3$EQUALS$AD2_9945_out0;
wire v$AD3$EQUALS$AD2_9946_out0;
wire v$ADD_5712_out0;
wire v$ADD_5713_out0;
wire v$ARBHALT0_1685_out0;
wire v$ARBHALT1_3700_out0;
wire v$ARR0_7237_out0;
wire v$ARR1_6305_out0;
wire v$AUTODISABLE_12944_out0;
wire v$AUTODISABLE_12945_out0;
wire v$AWR0_972_out0;
wire v$AWR1_11104_out0;
wire v$B$IS$RD_9476_out0;
wire v$B$IS$RD_9477_out0;
wire v$B0_2348_out0;
wire v$B0_2349_out0;
wire v$B0_2350_out0;
wire v$B0_2351_out0;
wire v$B0_2352_out0;
wire v$B0_2353_out0;
wire v$B0_2354_out0;
wire v$B0_2355_out0;
wire v$B0_2356_out0;
wire v$B0_2357_out0;
wire v$B0_2358_out0;
wire v$B0_2359_out0;
wire v$B0_2360_out0;
wire v$B0_2361_out0;
wire v$B0_2362_out0;
wire v$B0_2363_out0;
wire v$B0_2364_out0;
wire v$B0_2365_out0;
wire v$B0_2366_out0;
wire v$B0_2367_out0;
wire v$B0_2368_out0;
wire v$B0_2369_out0;
wire v$B0_2370_out0;
wire v$B0_2371_out0;
wire v$B1_9617_out0;
wire v$B1_9618_out0;
wire v$B1_9619_out0;
wire v$B1_9620_out0;
wire v$B1_9621_out0;
wire v$B1_9622_out0;
wire v$B1_9623_out0;
wire v$B1_9624_out0;
wire v$B1_9625_out0;
wire v$B1_9626_out0;
wire v$B1_9627_out0;
wire v$B1_9628_out0;
wire v$B1_9629_out0;
wire v$B1_9630_out0;
wire v$B1_9631_out0;
wire v$B1_9632_out0;
wire v$B1_9633_out0;
wire v$B1_9634_out0;
wire v$B1_9635_out0;
wire v$B1_9636_out0;
wire v$B1_9637_out0;
wire v$B1_9638_out0;
wire v$B1_9639_out0;
wire v$B1_9640_out0;
wire v$B2_11696_out0;
wire v$B2_11697_out0;
wire v$B2_11698_out0;
wire v$B2_11699_out0;
wire v$B2_11700_out0;
wire v$B2_11701_out0;
wire v$B2_11702_out0;
wire v$B2_11703_out0;
wire v$B2_11704_out0;
wire v$B2_11705_out0;
wire v$B2_11706_out0;
wire v$B2_11707_out0;
wire v$B2_11708_out0;
wire v$B2_11709_out0;
wire v$B2_11710_out0;
wire v$B2_11711_out0;
wire v$B2_11712_out0;
wire v$B2_11713_out0;
wire v$B2_11714_out0;
wire v$B2_11715_out0;
wire v$B2_11716_out0;
wire v$B2_11717_out0;
wire v$B2_11718_out0;
wire v$B2_11719_out0;
wire v$B3_12638_out0;
wire v$B3_12639_out0;
wire v$B3_12640_out0;
wire v$B3_12641_out0;
wire v$B3_12642_out0;
wire v$B3_12643_out0;
wire v$B3_12644_out0;
wire v$B3_12645_out0;
wire v$B3_12646_out0;
wire v$B3_12647_out0;
wire v$B3_12648_out0;
wire v$B3_12649_out0;
wire v$B3_12650_out0;
wire v$B3_12651_out0;
wire v$B3_12652_out0;
wire v$B3_12653_out0;
wire v$B3_12654_out0;
wire v$B3_12655_out0;
wire v$B3_12656_out0;
wire v$B3_12657_out0;
wire v$B3_12658_out0;
wire v$B3_12659_out0;
wire v$B3_12660_out0;
wire v$B3_12661_out0;
wire v$B4_11979_out0;
wire v$B4_11980_out0;
wire v$B4_11981_out0;
wire v$B4_11982_out0;
wire v$C11_2340_out0;
wire v$C11_2341_out0;
wire v$C1_10973_out0;
wire v$C1_10974_out0;
wire v$C1_10975_out0;
wire v$C1_10976_out0;
wire v$C1_11126_out0;
wire v$C1_11127_out0;
wire v$C1_12157_out0;
wire v$C1_12158_out0;
wire v$C1_12159_out0;
wire v$C1_12160_out0;
wire v$C1_12492_out0;
wire v$C1_12493_out0;
wire v$C1_12494_out0;
wire v$C1_12495_out0;
wire v$C1_12496_out0;
wire v$C1_12497_out0;
wire v$C1_1535_out0;
wire v$C1_1536_out0;
wire v$C1_1537_out0;
wire v$C1_1538_out0;
wire v$C1_1539_out0;
wire v$C1_1540_out0;
wire v$C1_1541_out0;
wire v$C1_1542_out0;
wire v$C1_1543_out0;
wire v$C1_1544_out0;
wire v$C1_1545_out0;
wire v$C1_1546_out0;
wire v$C1_3012_out0;
wire v$C1_3013_out0;
wire v$C1_3681_out0;
wire v$C1_3682_out0;
wire v$C1_3965_out0;
wire v$C1_3972_out0;
wire v$C1_3978_out0;
wire v$C1_3982_out0;
wire v$C1_3987_out0;
wire v$C1_3992_out0;
wire v$C1_3997_out0;
wire v$C1_4004_out0;
wire v$C1_4010_out0;
wire v$C1_4014_out0;
wire v$C1_4019_out0;
wire v$C1_4024_out0;
wire v$C1_4454_out0;
wire v$C1_4455_out0;
wire v$C1_5478_out0;
wire v$C1_5482_out0;
wire v$C1_703_out0;
wire v$C1_704_out0;
wire v$C1_739_out0;
wire v$C1_740_out0;
wire v$C1_8496_out0;
wire v$C1_8497_out0;
wire v$C2_10483_out0;
wire v$C2_10484_out0;
wire v$C2_10485_out0;
wire v$C2_10486_out0;
wire v$C2_105_out0;
wire v$C2_111_out0;
wire v$C2_11391_out0;
wire v$C2_11392_out0;
wire v$C2_11416_out0;
wire v$C2_11417_out0;
wire v$C2_11418_out0;
wire v$C2_11419_out0;
wire v$C2_11444_out0;
wire v$C2_11445_out0;
wire v$C2_11446_out0;
wire v$C2_11447_out0;
wire v$C2_115_out0;
wire v$C2_12078_out0;
wire v$C2_12079_out0;
wire v$C2_120_out0;
wire v$C2_125_out0;
wire v$C2_13020_out0;
wire v$C2_13021_out0;
wire v$C2_130_out0;
wire v$C2_137_out0;
wire v$C2_143_out0;
wire v$C2_147_out0;
wire v$C2_152_out0;
wire v$C2_1568_out0;
wire v$C2_1569_out0;
wire v$C2_157_out0;
wire v$C2_1736_out0;
wire v$C2_1737_out0;
wire v$C2_2336_out0;
wire v$C2_2337_out0;
wire v$C2_465_out0;
wire v$C2_466_out0;
wire v$C2_5163_out0;
wire v$C2_5164_out0;
wire v$C2_5165_out0;
wire v$C2_5166_out0;
wire v$C2_5167_out0;
wire v$C2_5168_out0;
wire v$C2_693_out0;
wire v$C2_694_out0;
wire v$C2_9087_out0;
wire v$C2_9088_out0;
wire v$C2_98_out0;
wire v$C3_12863_out0;
wire v$C3_12864_out0;
wire v$C3_13205_out0;
wire v$C3_13206_out0;
wire v$C3_3631_out0;
wire v$C3_3632_out0;
wire v$C3_587_out0;
wire v$C3_588_out0;
wire v$C3_7504_out0;
wire v$C3_7505_out0;
wire v$C3_9093_out0;
wire v$C3_9094_out0;
wire v$C3_9095_out0;
wire v$C3_9096_out0;
wire v$C4_10175_out0;
wire v$C4_10176_out0;
wire v$C4_10177_out0;
wire v$C4_10178_out0;
wire v$C4_1692_out0;
wire v$C4_1693_out0;
wire v$C4_2467_out0;
wire v$C4_2468_out0;
wire v$C4_4391_out0;
wire v$C4_4392_out0;
wire v$C5_6002_out0;
wire v$C5_6003_out0;
wire v$C5_6004_out0;
wire v$C5_6005_out0;
wire v$C6_1357_out0;
wire v$C6_1358_out0;
wire v$C6_1359_out0;
wire v$C6_1360_out0;
wire v$C6_7384_out0;
wire v$C6_7385_out0;
wire v$C6_7386_out0;
wire v$C6_7387_out0;
wire v$C6_7388_out0;
wire v$C6_7389_out0;
wire v$C6_7390_out0;
wire v$C6_7391_out0;
wire v$C6_7392_out0;
wire v$C6_7393_out0;
wire v$C6_7394_out0;
wire v$C6_7395_out0;
wire v$C6_7396_out0;
wire v$C6_7397_out0;
wire v$C6_7398_out0;
wire v$C6_7399_out0;
wire v$C6_7400_out0;
wire v$C6_7401_out0;
wire v$C6_7402_out0;
wire v$C6_7403_out0;
wire v$C6_7404_out0;
wire v$C6_7405_out0;
wire v$C6_7406_out0;
wire v$C6_7407_out0;
wire v$C6_775_out0;
wire v$C6_776_out0;
wire v$C6_8186_out0;
wire v$C6_8187_out0;
wire v$C7_274_out0;
wire v$C7_275_out0;
wire v$CAPTURE_207_out0;
wire v$CAPTURE_208_out0;
wire v$CARRY_3395_out0;
wire v$CARRY_3396_out0;
wire v$CARRY_7187_out0;
wire v$CARRY_7188_out0;
wire v$CARRY_9008_out0;
wire v$CARRY_9009_out0;
wire v$CHECKPARITY_557_out0;
wire v$CHECKPARITY_558_out0;
wire v$CIN$EXEC1_792_out0;
wire v$CIN$EXEC1_793_out0;
wire v$CIN_11849_out0;
wire v$CIN_11850_out0;
wire v$CIN_11851_out0;
wire v$CIN_11852_out0;
wire v$CIN_11853_out0;
wire v$CIN_11854_out0;
wire v$CIN_11855_out0;
wire v$CIN_11856_out0;
wire v$CIN_11857_out0;
wire v$CIN_11858_out0;
wire v$CIN_11859_out0;
wire v$CIN_11860_out0;
wire v$CIN_11861_out0;
wire v$CIN_11862_out0;
wire v$CIN_11863_out0;
wire v$CIN_11864_out0;
wire v$CIN_11865_out0;
wire v$CIN_11866_out0;
wire v$CIN_11867_out0;
wire v$CIN_11868_out0;
wire v$CIN_11869_out0;
wire v$CIN_11870_out0;
wire v$CIN_11871_out0;
wire v$CIN_11872_out0;
wire v$CIN_12952_out0;
wire v$CIN_12953_out0;
wire v$CIN_12954_out0;
wire v$CIN_12955_out0;
wire v$CIN_12956_out0;
wire v$CIN_12957_out0;
wire v$CIN_12958_out0;
wire v$CIN_12959_out0;
wire v$CIN_2594_out0;
wire v$CIN_2595_out0;
wire v$CIN_2596_out0;
wire v$CIN_2597_out0;
wire v$CIN_2598_out0;
wire v$CIN_2599_out0;
wire v$CIN_2600_out0;
wire v$CIN_2601_out0;
wire v$CIN_2602_out0;
wire v$CIN_2603_out0;
wire v$CIN_2604_out0;
wire v$CIN_2605_out0;
wire v$CIN_2606_out0;
wire v$CIN_2607_out0;
wire v$CIN_2608_out0;
wire v$CIN_2609_out0;
wire v$CIN_2610_out0;
wire v$CIN_2611_out0;
wire v$CIN_2612_out0;
wire v$CIN_2613_out0;
wire v$CIN_2614_out0;
wire v$CIN_2615_out0;
wire v$CIN_2616_out0;
wire v$CIN_2617_out0;
wire v$CLEAR_13091_out0;
wire v$CLEAR_13092_out0;
wire v$CLK4_11784_out0;
wire v$CLK4_11785_out0;
wire v$CLK4_12743_out0;
wire v$CLK4_12744_out0;
wire v$CLK4_1439_out0;
wire v$CLK4_1440_out0;
wire v$CLK4_2409_out0;
wire v$CLK4_2410_out0;
wire v$CLK4_4804_out0;
wire v$CLK4_4805_out0;
wire v$CLK4_6074_out0;
wire v$CLK4_6075_out0;
wire v$CLK4_7986_out0;
wire v$CLK4_7987_out0;
wire v$CLRINTERRUPTS_276_out0;
wire v$CLRINTERRUPTS_277_out0;
wire v$CLR_3083_out0;
wire v$CLR_3084_out0;
wire v$COMP$H$OUT_4646_out0;
wire v$COMP$H$OUT_4647_out0;
wire v$COMP$L$OUT_7515_out0;
wire v$COMP$L$OUT_7516_out0;
wire v$COUNTEREN_828_out0;
wire v$COUNTEREN_829_out0;
wire v$COUNTEREN_9016_out0;
wire v$COUNTEREN_9017_out0;
wire v$COUNTERINTERRUPT_10189_out0;
wire v$COUNTERINTERRUPT_10190_out0;
wire v$COUT$EXEC1_796_out0;
wire v$COUT$EXEC1_797_out0;
wire v$COUT$HALF_70_out0;
wire v$COUT$HALF_71_out0;
wire v$COUT_3407_out0;
wire v$COUT_3408_out0;
wire v$COUT_5613_out0;
wire v$COUT_5614_out0;
wire v$COUT_5615_out0;
wire v$COUT_5616_out0;
wire v$COUT_5617_out0;
wire v$COUT_5618_out0;
wire v$COUT_5619_out0;
wire v$COUT_5620_out0;
wire v$COUT_5621_out0;
wire v$COUT_5622_out0;
wire v$COUT_5623_out0;
wire v$COUT_5624_out0;
wire v$COUT_5625_out0;
wire v$COUT_5626_out0;
wire v$COUT_5627_out0;
wire v$COUT_5628_out0;
wire v$COUT_5629_out0;
wire v$COUT_5630_out0;
wire v$COUT_5631_out0;
wire v$COUT_5632_out0;
wire v$COUT_5633_out0;
wire v$COUT_5634_out0;
wire v$COUT_5635_out0;
wire v$COUT_5636_out0;
wire v$COUT_5766_out0;
wire v$COUT_5767_out0;
wire v$COUT_7042_out0;
wire v$COUT_7043_out0;
wire v$COUT_7044_out0;
wire v$COUT_7045_out0;
wire v$COUT_7046_out0;
wire v$COUT_7047_out0;
wire v$COUT_7048_out0;
wire v$COUT_7049_out0;
wire v$COUT_7050_out0;
wire v$COUT_7051_out0;
wire v$COUT_7052_out0;
wire v$COUT_7053_out0;
wire v$COUT_7054_out0;
wire v$COUT_7055_out0;
wire v$COUT_7056_out0;
wire v$COUT_7057_out0;
wire v$COUT_7058_out0;
wire v$COUT_7059_out0;
wire v$COUT_7060_out0;
wire v$COUT_7061_out0;
wire v$COUT_7062_out0;
wire v$COUT_7063_out0;
wire v$COUT_7064_out0;
wire v$COUT_7065_out0;
wire v$C_11110_out0;
wire v$C_11111_out0;
wire v$C_1917_out0;
wire v$C_1918_out0;
wire v$C_2344_out0;
wire v$C_2345_out0;
wire v$C_4069_out0;
wire v$C_4070_out0;
wire v$C_6570_out0;
wire v$C_6571_out0;
wire v$CheckParity_13308_out0;
wire v$CheckParity_13309_out0;
wire v$Clear_10010_out0;
wire v$Clear_10011_out0;
wire v$Clear_8404_out0;
wire v$Clear_8405_out0;
wire v$D1_9486_out0;
wire v$D1_9486_out1;
wire v$D1_9486_out2;
wire v$D1_9486_out3;
wire v$D1_9487_out0;
wire v$D1_9487_out1;
wire v$D1_9487_out2;
wire v$D1_9487_out3;
wire v$DATA$DEPENDENCY_4171_out0;
wire v$DATA$DEPENDENCY_4172_out0;
wire v$DATA$PROCESS$WB_12623_out0;
wire v$DATA$PROCESS$WB_12624_out0;
wire v$DISABLEINTERRUPTS_10305_out0;
wire v$DISABLEINTERRUPTS_10306_out0;
wire v$DM1_11395_out0;
wire v$DM1_11395_out1;
wire v$EDGE0_2712_out0;
wire v$EDGE0_2713_out0;
wire v$EDGE0_3772_out0;
wire v$EDGE0_3773_out0;
wire v$EDGE1_10589_out0;
wire v$EDGE1_10590_out0;
wire v$EDGE1_12216_out0;
wire v$EDGE1_12217_out0;
wire v$EDGE2_12853_out0;
wire v$EDGE2_12854_out0;
wire v$EDGE2_4761_out0;
wire v$EDGE2_4762_out0;
wire v$EDGE3_1168_out0;
wire v$EDGE3_1169_out0;
wire v$EDGE3_7278_out0;
wire v$EDGE3_7279_out0;
wire v$ENABLEINTERRUPTS_12084_out0;
wire v$ENABLEINTERRUPTS_12085_out0;
wire v$ENABLEINTERRUPTS_8182_out0;
wire v$ENABLEINTERRUPTS_8183_out0;
wire v$ENCODED0_9415_out0;
wire v$ENCODED0_9416_out0;
wire v$ENCODED1_6496_out0;
wire v$ENCODED1_6497_out0;
wire v$END1_4730_out0;
wire v$END1_4731_out0;
wire v$END1_4747_out0;
wire v$END1_4748_out0;
wire v$END4_1971_out0;
wire v$END4_1972_out0;
wire v$END4_5637_out0;
wire v$END4_5638_out0;
wire v$END6_5096_out0;
wire v$END6_5097_out0;
wire v$END_10986_out0;
wire v$END_10987_out0;
wire v$END_12098_out0;
wire v$END_12099_out0;
wire v$END_5603_out0;
wire v$END_5604_out0;
wire v$ENMODE_5281_out0;
wire v$ENMODE_5282_out0;
wire v$ENMODE_9952_out0;
wire v$ENMODE_9953_out0;
wire v$EN_11112_out0;
wire v$EN_11113_out0;
wire v$EN_11490_out0;
wire v$EN_11491_out0;
wire v$EN_11492_out0;
wire v$EN_11493_out0;
wire v$EN_11494_out0;
wire v$EN_11495_out0;
wire v$EN_11496_out0;
wire v$EN_11497_out0;
wire v$EN_12029_out0;
wire v$EN_12030_out0;
wire v$EN_12031_out0;
wire v$EN_12032_out0;
wire v$EN_12033_out0;
wire v$EN_12034_out0;
wire v$EN_12035_out0;
wire v$EN_12036_out0;
wire v$EN_3165_out0;
wire v$EN_3166_out0;
wire v$EN_3167_out0;
wire v$EN_3168_out0;
wire v$EN_3169_out0;
wire v$EN_3170_out0;
wire v$EN_3171_out0;
wire v$EN_3172_out0;
wire v$EN_3173_out0;
wire v$EN_3174_out0;
wire v$EN_3175_out0;
wire v$EN_3176_out0;
wire v$EN_3585_out0;
wire v$EN_3586_out0;
wire v$EN_3587_out0;
wire v$EN_3588_out0;
wire v$EN_3589_out0;
wire v$EN_3590_out0;
wire v$EN_3591_out0;
wire v$EN_3592_out0;
wire v$EN_3593_out0;
wire v$EN_3594_out0;
wire v$EN_3595_out0;
wire v$EN_3596_out0;
wire v$EN_3597_out0;
wire v$EN_3598_out0;
wire v$EN_3599_out0;
wire v$EN_3600_out0;
wire v$EN_3601_out0;
wire v$EN_3602_out0;
wire v$EN_3603_out0;
wire v$EN_3604_out0;
wire v$EN_5389_out0;
wire v$EN_5390_out0;
wire v$EN_5391_out0;
wire v$EN_5392_out0;
wire v$EN_5393_out0;
wire v$EN_5394_out0;
wire v$EN_5395_out0;
wire v$EN_5396_out0;
wire v$EN_5397_out0;
wire v$EN_5398_out0;
wire v$EN_5399_out0;
wire v$EN_5400_out0;
wire v$EN_561_out0;
wire v$EN_562_out0;
wire v$EN_563_out0;
wire v$EN_564_out0;
wire v$EN_565_out0;
wire v$EN_566_out0;
wire v$EN_567_out0;
wire v$EN_568_out0;
wire v$EN_569_out0;
wire v$EN_570_out0;
wire v$EN_571_out0;
wire v$EN_572_out0;
wire v$EN_573_out0;
wire v$EN_574_out0;
wire v$EN_575_out0;
wire v$EN_576_out0;
wire v$EN_577_out0;
wire v$EN_578_out0;
wire v$EN_579_out0;
wire v$EN_580_out0;
wire v$EN_6318_out0;
wire v$EN_6319_out0;
wire v$EPARITY_13014_out0;
wire v$EPARITY_13015_out0;
wire v$EQ$LDST_12234_out0;
wire v$EQ$LDST_12235_out0;
wire v$EQ10_3914_out0;
wire v$EQ10_3915_out0;
wire v$EQ10_3916_out0;
wire v$EQ10_3917_out0;
wire v$EQ10_6613_out0;
wire v$EQ10_6614_out0;
wire v$EQ10_8978_out0;
wire v$EQ10_8979_out0;
wire v$EQ11_4157_out0;
wire v$EQ11_4158_out0;
wire v$EQ11_4159_out0;
wire v$EQ11_4160_out0;
wire v$EQ11_7677_out0;
wire v$EQ11_7678_out0;
wire v$EQ11_9167_out0;
wire v$EQ11_9168_out0;
wire v$EQ12_10420_out0;
wire v$EQ12_10421_out0;
wire v$EQ12_761_out0;
wire v$EQ12_762_out0;
wire v$EQ12_8848_out0;
wire v$EQ12_8849_out0;
wire v$EQ12_9356_out0;
wire v$EQ12_9357_out0;
wire v$EQ12_9358_out0;
wire v$EQ12_9359_out0;
wire v$EQ13_13201_out0;
wire v$EQ13_13202_out0;
wire v$EQ13_3617_out0;
wire v$EQ13_3618_out0;
wire v$EQ13_6370_out0;
wire v$EQ13_6371_out0;
wire v$EQ13_6491_out0;
wire v$EQ13_6492_out0;
wire v$EQ13_6493_out0;
wire v$EQ13_6494_out0;
wire v$EQ14_3647_out0;
wire v$EQ14_3648_out0;
wire v$EQ14_3649_out0;
wire v$EQ14_3650_out0;
wire v$EQ14_3730_out0;
wire v$EQ14_3731_out0;
wire v$EQ14_7897_out0;
wire v$EQ14_7898_out0;
wire v$EQ15_11158_out0;
wire v$EQ15_11159_out0;
wire v$EQ15_11160_out0;
wire v$EQ15_11161_out0;
wire v$EQ15_12096_out0;
wire v$EQ15_12097_out0;
wire v$EQ16_5760_out0;
wire v$EQ16_5761_out0;
wire v$EQ16_5762_out0;
wire v$EQ16_5763_out0;
wire v$EQ16_785_out0;
wire v$EQ16_786_out0;
wire v$EQ17_3906_out0;
wire v$EQ17_3907_out0;
wire v$EQ17_3908_out0;
wire v$EQ17_3909_out0;
wire v$EQ18_8460_out0;
wire v$EQ18_8461_out0;
wire v$EQ18_8462_out0;
wire v$EQ18_8463_out0;
wire v$EQ19_3689_out0;
wire v$EQ19_3690_out0;
wire v$EQ19_3691_out0;
wire v$EQ19_3692_out0;
wire v$EQ1_10605_out0;
wire v$EQ1_10606_out0;
wire v$EQ1_10629_out0;
wire v$EQ1_10630_out0;
wire v$EQ1_11291_out0;
wire v$EQ1_11292_out0;
wire v$EQ1_11375_out0;
wire v$EQ1_11376_out0;
wire v$EQ1_11412_out0;
wire v$EQ1_11413_out0;
wire v$EQ1_13237_out0;
wire v$EQ1_13238_out0;
wire v$EQ1_1429_out0;
wire v$EQ1_1430_out0;
wire v$EQ1_1585_out0;
wire v$EQ1_1586_out0;
wire v$EQ1_1719_out0;
wire v$EQ1_1720_out0;
wire v$EQ1_1925_out0;
wire v$EQ1_1926_out0;
wire v$EQ1_2809_out0;
wire v$EQ1_2810_out0;
wire v$EQ1_3449_out0;
wire v$EQ1_3450_out0;
wire v$EQ1_3457_out0;
wire v$EQ1_3458_out0;
wire v$EQ1_4702_out0;
wire v$EQ1_4703_out0;
wire v$EQ1_5014_out0;
wire v$EQ1_5015_out0;
wire v$EQ1_6960_out0;
wire v$EQ1_6961_out0;
wire v$EQ1_7467_out0;
wire v$EQ1_7468_out0;
wire v$EQ1_8585_out0;
wire v$EQ1_8586_out0;
wire v$EQ1_8927_out0;
wire v$EQ1_8928_out0;
wire v$EQ1_8984_out0;
wire v$EQ1_8985_out0;
wire v$EQ1_8986_out0;
wire v$EQ1_8987_out0;
wire v$EQ1_9709_out0;
wire v$EQ1_9710_out0;
wire v$EQ20_6666_out0;
wire v$EQ20_6667_out0;
wire v$EQ20_6668_out0;
wire v$EQ20_6669_out0;
wire v$EQ21_2017_out0;
wire v$EQ21_2018_out0;
wire v$EQ21_2019_out0;
wire v$EQ21_2020_out0;
wire v$EQ22_1599_out0;
wire v$EQ22_1600_out0;
wire v$EQ22_1601_out0;
wire v$EQ22_1602_out0;
wire v$EQ23_1913_out0;
wire v$EQ23_1914_out0;
wire v$EQ23_1915_out0;
wire v$EQ23_1916_out0;
wire v$EQ24_1445_out0;
wire v$EQ24_1446_out0;
wire v$EQ24_1447_out0;
wire v$EQ24_1448_out0;
wire v$EQ2_11025_out0;
wire v$EQ2_11026_out0;
wire v$EQ2_11320_out0;
wire v$EQ2_11321_out0;
wire v$EQ2_11498_out0;
wire v$EQ2_11499_out0;
wire v$EQ2_11951_out0;
wire v$EQ2_11952_out0;
wire v$EQ2_13294_out0;
wire v$EQ2_13295_out0;
wire v$EQ2_1923_out0;
wire v$EQ2_1924_out0;
wire v$EQ2_2910_out0;
wire v$EQ2_2911_out0;
wire v$EQ2_5448_out0;
wire v$EQ2_5449_out0;
wire v$EQ2_7104_out0;
wire v$EQ2_7105_out0;
wire v$EQ2_7440_out0;
wire v$EQ2_7441_out0;
wire v$EQ2_8518_out0;
wire v$EQ2_8519_out0;
wire v$EQ2_9180_out0;
wire v$EQ2_9181_out0;
wire v$EQ2_9605_out0;
wire v$EQ2_9606_out0;
wire v$EQ2_9607_out0;
wire v$EQ2_9608_out0;
wire v$EQ2_9691_out0;
wire v$EQ2_9692_out0;
wire v$EQ3_10598_out0;
wire v$EQ3_10599_out0;
wire v$EQ3_10785_out0;
wire v$EQ3_10786_out0;
wire v$EQ3_11624_out0;
wire v$EQ3_11625_out0;
wire v$EQ3_12697_out0;
wire v$EQ3_12698_out0;
wire v$EQ3_1515_out0;
wire v$EQ3_1516_out0;
wire v$EQ3_2888_out0;
wire v$EQ3_2889_out0;
wire v$EQ3_3683_out0;
wire v$EQ3_3684_out0;
wire v$EQ3_3768_out0;
wire v$EQ3_3769_out0;
wire v$EQ3_4843_out0;
wire v$EQ3_4844_out0;
wire v$EQ3_5414_out0;
wire v$EQ3_5415_out0;
wire v$EQ3_7532_out0;
wire v$EQ3_7533_out0;
wire v$EQ3_7911_out0;
wire v$EQ3_7912_out0;
wire v$EQ3_9316_out0;
wire v$EQ3_9317_out0;
wire v$EQ3_9693_out0;
wire v$EQ3_9694_out0;
wire v$EQ3_991_out0;
wire v$EQ3_992_out0;
wire v$EQ3_993_out0;
wire v$EQ3_994_out0;
wire v$EQ4_11584_out0;
wire v$EQ4_11585_out0;
wire v$EQ4_11654_out0;
wire v$EQ4_11655_out0;
wire v$EQ4_11767_out0;
wire v$EQ4_11768_out0;
wire v$EQ4_13241_out0;
wire v$EQ4_13242_out0;
wire v$EQ4_13243_out0;
wire v$EQ4_13244_out0;
wire v$EQ4_1519_out0;
wire v$EQ4_1520_out0;
wire v$EQ4_1767_out0;
wire v$EQ4_1768_out0;
wire v$EQ4_3659_out0;
wire v$EQ4_3660_out0;
wire v$EQ4_6379_out0;
wire v$EQ4_6380_out0;
wire v$EQ4_6581_out0;
wire v$EQ4_6582_out0;
wire v$EQ4_8382_out0;
wire v$EQ4_8383_out0;
wire v$EQ5_1062_out0;
wire v$EQ5_1063_out0;
wire v$EQ5_1729_out0;
wire v$EQ5_1730_out0;
wire v$EQ5_2013_out0;
wire v$EQ5_2014_out0;
wire v$EQ5_2015_out0;
wire v$EQ5_2016_out0;
wire v$EQ5_2252_out0;
wire v$EQ5_2253_out0;
wire v$EQ5_3256_out0;
wire v$EQ5_3257_out0;
wire v$EQ5_6345_out0;
wire v$EQ5_6346_out0;
wire v$EQ5_6738_out0;
wire v$EQ5_6739_out0;
wire v$EQ5_733_out0;
wire v$EQ5_734_out0;
wire v$EQ5_9756_out0;
wire v$EQ5_9757_out0;
wire v$EQ6_11090_out0;
wire v$EQ6_11091_out0;
wire v$EQ6_11337_out0;
wire v$EQ6_11338_out0;
wire v$EQ6_11402_out0;
wire v$EQ6_11403_out0;
wire v$EQ6_2668_out0;
wire v$EQ6_2669_out0;
wire v$EQ6_3671_out0;
wire v$EQ6_3672_out0;
wire v$EQ6_3673_out0;
wire v$EQ6_3674_out0;
wire v$EQ6_4423_out0;
wire v$EQ6_4424_out0;
wire v$EQ6_773_out0;
wire v$EQ6_774_out0;
wire v$EQ7_11947_out0;
wire v$EQ7_11948_out0;
wire v$EQ7_13267_out0;
wire v$EQ7_13268_out0;
wire v$EQ7_201_out0;
wire v$EQ7_202_out0;
wire v$EQ7_2208_out0;
wire v$EQ7_2209_out0;
wire v$EQ7_2788_out0;
wire v$EQ7_2789_out0;
wire v$EQ7_2790_out0;
wire v$EQ7_2791_out0;
wire v$EQ8_217_out0;
wire v$EQ8_218_out0;
wire v$EQ8_9715_out0;
wire v$EQ8_9716_out0;
wire v$EQ8_9797_out0;
wire v$EQ8_9798_out0;
wire v$EQ8_9799_out0;
wire v$EQ8_9800_out0;
wire v$EQ9_12558_out0;
wire v$EQ9_12559_out0;
wire v$EQ9_12993_out0;
wire v$EQ9_12994_out0;
wire v$EQ9_5486_out0;
wire v$EQ9_5487_out0;
wire v$EQ9_9300_out0;
wire v$EQ9_9301_out0;
wire v$EQ9_9302_out0;
wire v$EQ9_9303_out0;
wire v$EQUAL_11046_out0;
wire v$EQUAL_11047_out0;
wire v$EQUAL_7464_out0;
wire v$EQUAL_7465_out0;
wire v$EQ_2185_out0;
wire v$EQ_2186_out0;
wire v$EQ_2421_out0;
wire v$EQ_2422_out0;
wire v$EQ_2994_out0;
wire v$EQ_2995_out0;
wire v$EQ_360_out0;
wire v$EQ_361_out0;
wire v$EQ_4165_out0;
wire v$EQ_4166_out0;
wire v$EQ_8992_out0;
wire v$EQ_8993_out0;
wire v$EQ_9954_out0;
wire v$EQ_9955_out0;
wire v$ERR_8428_out0;
wire v$ERR_8429_out0;
wire v$EVENPARITY_9157_out0;
wire v$EVENPARITY_9158_out0;
wire v$EXEC1$FPU_9221_out0;
wire v$EXEC1$FPU_9222_out0;
wire v$EXEC1$VIEW$MULTIPLIER_11514_out0;
wire v$EXEC1$VIEW$MULTIPLIER_11515_out0;
wire v$EXEC1_12950_out0;
wire v$EXEC1_12951_out0;
wire v$EXEC1_13169_out0;
wire v$EXEC1_13170_out0;
wire v$EXEC1_13347_out0;
wire v$EXEC1_13348_out0;
wire v$EXEC1_2564_out0;
wire v$EXEC1_2565_out0;
wire v$EXEC1_5456_out0;
wire v$EXEC1_5457_out0;
wire v$EXEC1_5458_out0;
wire v$EXEC1_5459_out0;
wire v$EXEC1_5460_out0;
wire v$EXEC1_5461_out0;
wire v$EXEC1_5462_out0;
wire v$EXEC1_5463_out0;
wire v$EXEC1_5464_out0;
wire v$EXEC1_5465_out0;
wire v$EXEC1_5466_out0;
wire v$EXEC1_5467_out0;
wire v$EXEC1_5468_out0;
wire v$EXEC1_5469_out0;
wire v$EXEC1_5470_out0;
wire v$EXEC1_5471_out0;
wire v$EXEC1_5472_out0;
wire v$EXEC1_5473_out0;
wire v$EXEC1_5474_out0;
wire v$EXEC1_5475_out0;
wire v$EXEC1_5476_out0;
wire v$EXEC1_5477_out0;
wire v$EXEC1_6827_out0;
wire v$EXEC1_6828_out0;
wire v$EXEC2_1091_out0;
wire v$EXEC2_1092_out0;
wire v$EXEC2_11098_out0;
wire v$EXEC2_11099_out0;
wire v$EXEC2_11473_out0;
wire v$EXEC2_11474_out0;
wire v$EXEC2_12457_out0;
wire v$EXEC2_12458_out0;
wire v$EXEC2_2720_out0;
wire v$EXEC2_2721_out0;
wire v$EXEC2_3042_out0;
wire v$EXEC2_3043_out0;
wire v$EXEC2_358_out0;
wire v$EXEC2_359_out0;
wire v$EXEC2_461_out0;
wire v$EXEC2_462_out0;
wire v$EXEC2_5520_out0;
wire v$EXEC2_5521_out0;
wire v$EXEC2_5557_out0;
wire v$EXEC2_5558_out0;
wire v$EXEC2_6435_out0;
wire v$EXEC2_6436_out0;
wire v$EXEC2_6611_out0;
wire v$EXEC2_6612_out0;
wire v$EXEC2_701_out0;
wire v$EXEC2_702_out0;
wire v$EXP$SAME_11626_out0;
wire v$EXP$SAME_11627_out0;
wire v$EXP$SAME_1875_out0;
wire v$EXP$SAME_1876_out0;
wire v$EXP$SAME_408_out0;
wire v$EXP$SAME_409_out0;
wire v$EXTHALT_12666_out0;
wire v$EXTHALT_12667_out0;
wire v$EXTHALT_4456_out0;
wire v$EXTHALT_4457_out0;
wire v$E_12165_out0;
wire v$E_12166_out0;
wire v$Error_2475_out0;
wire v$Error_2476_out0;
wire v$F0_11052_out0;
wire v$F0_11053_out0;
wire v$F1_2195_out0;
wire v$F1_2196_out0;
wire v$F2_7871_out0;
wire v$F2_7872_out0;
wire v$F3_5730_out0;
wire v$F3_5731_out0;
wire v$FPU$LOAD$B_7556_out0;
wire v$FPU$LOAD$B_7557_out0;
wire v$FPU$LOAD$STORE_7238_out0;
wire v$FPU$LOAD$STORE_7239_out0;
wire v$F_1111_out0;
wire v$F_1112_out0;
wire v$G10_10226_out0;
wire v$G10_10227_out0;
wire v$G10_11273_out0;
wire v$G10_11274_out0;
wire v$G10_11275_out0;
wire v$G10_11276_out0;
wire v$G10_1141_out0;
wire v$G10_1142_out0;
wire v$G10_11578_out0;
wire v$G10_11579_out0;
wire v$G10_12927_out0;
wire v$G10_12928_out0;
wire v$G10_13153_out0;
wire v$G10_13154_out0;
wire v$G10_1683_out0;
wire v$G10_1684_out0;
wire v$G10_2511_out0;
wire v$G10_2512_out0;
wire v$G10_4679_out0;
wire v$G10_4680_out0;
wire v$G10_471_out0;
wire v$G10_472_out0;
wire v$G10_605_out0;
wire v$G10_606_out0;
wire v$G10_607_out0;
wire v$G10_608_out0;
wire v$G10_609_out0;
wire v$G10_610_out0;
wire v$G10_611_out0;
wire v$G10_612_out0;
wire v$G10_613_out0;
wire v$G10_614_out0;
wire v$G10_615_out0;
wire v$G10_616_out0;
wire v$G10_617_out0;
wire v$G10_618_out0;
wire v$G10_619_out0;
wire v$G10_620_out0;
wire v$G10_621_out0;
wire v$G10_622_out0;
wire v$G10_623_out0;
wire v$G10_624_out0;
wire v$G10_625_out0;
wire v$G10_626_out0;
wire v$G10_627_out0;
wire v$G10_628_out0;
wire v$G10_629_out0;
wire v$G10_630_out0;
wire v$G10_631_out0;
wire v$G10_632_out0;
wire v$G10_633_out0;
wire v$G10_634_out0;
wire v$G10_635_out0;
wire v$G10_636_out0;
wire v$G10_637_out0;
wire v$G10_638_out0;
wire v$G10_639_out0;
wire v$G10_640_out0;
wire v$G10_641_out0;
wire v$G10_642_out0;
wire v$G10_643_out0;
wire v$G10_644_out0;
wire v$G10_645_out0;
wire v$G10_646_out0;
wire v$G10_647_out0;
wire v$G10_648_out0;
wire v$G10_649_out0;
wire v$G10_650_out0;
wire v$G10_651_out0;
wire v$G10_652_out0;
wire v$G10_653_out0;
wire v$G10_654_out0;
wire v$G10_655_out0;
wire v$G10_656_out0;
wire v$G10_657_out0;
wire v$G10_658_out0;
wire v$G10_659_out0;
wire v$G10_660_out0;
wire v$G10_661_out0;
wire v$G10_662_out0;
wire v$G10_663_out0;
wire v$G10_664_out0;
wire v$G10_6837_out0;
wire v$G10_6838_out0;
wire v$G10_8887_out0;
wire v$G10_8888_out0;
wire v$G10_9949_out0;
wire v$G10_9950_out0;
wire v$G10_9966_out0;
wire v$G10_9967_out0;
wire v$G11_10906_out0;
wire v$G11_10907_out0;
wire v$G11_10908_out0;
wire v$G11_10909_out0;
wire v$G11_10910_out0;
wire v$G11_10911_out0;
wire v$G11_10912_out0;
wire v$G11_10913_out0;
wire v$G11_10914_out0;
wire v$G11_10915_out0;
wire v$G11_10916_out0;
wire v$G11_10917_out0;
wire v$G11_10918_out0;
wire v$G11_10919_out0;
wire v$G11_10920_out0;
wire v$G11_10921_out0;
wire v$G11_10922_out0;
wire v$G11_10923_out0;
wire v$G11_10924_out0;
wire v$G11_10925_out0;
wire v$G11_10926_out0;
wire v$G11_10927_out0;
wire v$G11_10928_out0;
wire v$G11_10929_out0;
wire v$G11_1211_out0;
wire v$G11_1212_out0;
wire v$G11_12785_out0;
wire v$G11_12786_out0;
wire v$G11_1739_out0;
wire v$G11_1740_out0;
wire v$G11_1773_out0;
wire v$G11_1774_out0;
wire v$G11_1955_out0;
wire v$G11_1956_out0;
wire v$G11_3264_out0;
wire v$G11_3265_out0;
wire v$G11_5694_out0;
wire v$G11_5695_out0;
wire v$G11_5718_out0;
wire v$G11_5719_out0;
wire v$G11_5747_out0;
wire v$G11_5748_out0;
wire v$G11_6081_out0;
wire v$G11_6082_out0;
wire v$G11_6083_out0;
wire v$G11_6084_out0;
wire v$G11_6085_out0;
wire v$G11_6086_out0;
wire v$G11_6087_out0;
wire v$G11_6088_out0;
wire v$G11_6089_out0;
wire v$G11_6090_out0;
wire v$G11_6091_out0;
wire v$G11_6092_out0;
wire v$G11_6093_out0;
wire v$G11_6094_out0;
wire v$G11_6095_out0;
wire v$G11_6096_out0;
wire v$G11_6097_out0;
wire v$G11_6098_out0;
wire v$G11_6099_out0;
wire v$G11_6100_out0;
wire v$G11_6101_out0;
wire v$G11_6102_out0;
wire v$G11_6103_out0;
wire v$G11_6104_out0;
wire v$G11_6105_out0;
wire v$G11_6106_out0;
wire v$G11_6107_out0;
wire v$G11_6108_out0;
wire v$G11_6109_out0;
wire v$G11_6110_out0;
wire v$G11_6111_out0;
wire v$G11_6112_out0;
wire v$G11_6113_out0;
wire v$G11_6114_out0;
wire v$G11_6115_out0;
wire v$G11_6116_out0;
wire v$G11_6117_out0;
wire v$G11_6118_out0;
wire v$G11_6119_out0;
wire v$G11_6120_out0;
wire v$G11_6121_out0;
wire v$G11_6122_out0;
wire v$G11_6123_out0;
wire v$G11_6124_out0;
wire v$G11_6125_out0;
wire v$G11_6126_out0;
wire v$G11_6127_out0;
wire v$G11_6128_out0;
wire v$G11_6129_out0;
wire v$G11_6130_out0;
wire v$G11_6131_out0;
wire v$G11_6132_out0;
wire v$G11_6133_out0;
wire v$G11_6134_out0;
wire v$G11_6135_out0;
wire v$G11_6136_out0;
wire v$G11_6137_out0;
wire v$G11_6138_out0;
wire v$G11_6139_out0;
wire v$G11_6140_out0;
wire v$G11_6564_out0;
wire v$G11_6565_out0;
wire v$G11_7645_out0;
wire v$G11_7646_out0;
wire v$G11_823_out0;
wire v$G11_824_out0;
wire v$G11_8976_out0;
wire v$G11_8977_out0;
wire v$G11_9962_out0;
wire v$G11_9963_out0;
wire v$G12_10062_out0;
wire v$G12_10063_out0;
wire v$G12_11404_out0;
wire v$G12_11405_out0;
wire v$G12_1148_out0;
wire v$G12_1149_out0;
wire v$G12_11546_out0;
wire v$G12_11547_out0;
wire v$G12_11548_out0;
wire v$G12_11549_out0;
wire v$G12_11550_out0;
wire v$G12_11551_out0;
wire v$G12_11552_out0;
wire v$G12_11553_out0;
wire v$G12_11554_out0;
wire v$G12_11555_out0;
wire v$G12_11556_out0;
wire v$G12_11557_out0;
wire v$G12_11558_out0;
wire v$G12_11559_out0;
wire v$G12_11560_out0;
wire v$G12_11561_out0;
wire v$G12_11562_out0;
wire v$G12_11563_out0;
wire v$G12_11564_out0;
wire v$G12_11565_out0;
wire v$G12_11566_out0;
wire v$G12_11567_out0;
wire v$G12_11568_out0;
wire v$G12_11569_out0;
wire v$G12_2328_out0;
wire v$G12_2329_out0;
wire v$G12_3238_out0;
wire v$G12_3239_out0;
wire v$G12_4181_out0;
wire v$G12_4182_out0;
wire v$G12_6662_out0;
wire v$G12_6663_out0;
wire v$G12_7686_out0;
wire v$G12_7687_out0;
wire v$G12_7750_out0;
wire v$G12_7751_out0;
wire v$G12_9318_out0;
wire v$G12_9319_out0;
wire v$G12_995_out0;
wire v$G12_996_out0;
wire v$G13_10192_out0;
wire v$G13_10193_out0;
wire v$G13_10418_out0;
wire v$G13_10419_out0;
wire v$G13_11612_out0;
wire v$G13_11613_out0;
wire v$G13_186_out0;
wire v$G13_187_out0;
wire v$G13_3006_out0;
wire v$G13_3007_out0;
wire v$G13_3054_out0;
wire v$G13_3055_out0;
wire v$G13_3056_out0;
wire v$G13_3057_out0;
wire v$G13_3058_out0;
wire v$G13_3059_out0;
wire v$G13_3060_out0;
wire v$G13_3061_out0;
wire v$G13_3062_out0;
wire v$G13_3063_out0;
wire v$G13_3064_out0;
wire v$G13_3065_out0;
wire v$G13_3066_out0;
wire v$G13_3067_out0;
wire v$G13_3068_out0;
wire v$G13_3069_out0;
wire v$G13_3070_out0;
wire v$G13_3071_out0;
wire v$G13_3072_out0;
wire v$G13_3073_out0;
wire v$G13_3074_out0;
wire v$G13_3075_out0;
wire v$G13_3076_out0;
wire v$G13_3077_out0;
wire v$G13_5410_out0;
wire v$G13_5411_out0;
wire v$G13_6807_out0;
wire v$G13_6808_out0;
wire v$G13_7935_out0;
wire v$G13_7936_out0;
wire v$G13_883_out0;
wire v$G13_884_out0;
wire v$G13_9010_out0;
wire v$G13_9011_out0;
wire v$G14_10042_out0;
wire v$G14_10043_out0;
wire v$G14_10607_out0;
wire v$G14_10608_out0;
wire v$G14_11038_out0;
wire v$G14_11039_out0;
wire v$G14_12092_out0;
wire v$G14_12093_out0;
wire v$G14_13117_out0;
wire v$G14_13118_out0;
wire v$G14_3504_out0;
wire v$G14_3505_out0;
wire v$G14_3629_out0;
wire v$G14_3630_out0;
wire v$G14_4141_out0;
wire v$G14_4142_out0;
wire v$G14_4440_out0;
wire v$G14_4441_out0;
wire v$G14_7830_out0;
wire v$G14_7831_out0;
wire v$G14_8284_out0;
wire v$G14_8285_out0;
wire v$G14_8286_out0;
wire v$G14_8287_out0;
wire v$G14_867_out0;
wire v$G14_868_out0;
wire v$G15_1030_out0;
wire v$G15_1031_out0;
wire v$G15_1205_out0;
wire v$G15_1206_out0;
wire v$G15_12619_out0;
wire v$G15_12620_out0;
wire v$G15_13187_out0;
wire v$G15_13188_out0;
wire v$G15_1579_out0;
wire v$G15_1580_out0;
wire v$G15_2890_out0;
wire v$G15_2891_out0;
wire v$G15_3722_out0;
wire v$G15_3723_out0;
wire v$G15_8965_out0;
wire v$G15_8966_out0;
wire v$G15_8990_out0;
wire v$G15_8991_out0;
wire v$G15_9165_out0;
wire v$G15_9166_out0;
wire v$G15_9195_out0;
wire v$G15_9196_out0;
wire v$G15_9197_out0;
wire v$G15_9198_out0;
wire v$G15_9199_out0;
wire v$G15_9200_out0;
wire v$G15_9201_out0;
wire v$G15_9202_out0;
wire v$G15_9203_out0;
wire v$G15_9204_out0;
wire v$G15_9205_out0;
wire v$G15_9206_out0;
wire v$G15_9207_out0;
wire v$G15_9208_out0;
wire v$G15_9209_out0;
wire v$G15_9210_out0;
wire v$G15_9211_out0;
wire v$G15_9212_out0;
wire v$G15_9213_out0;
wire v$G15_9214_out0;
wire v$G15_9215_out0;
wire v$G15_9216_out0;
wire v$G15_9217_out0;
wire v$G15_9218_out0;
wire v$G15_9960_out0;
wire v$G15_9961_out0;
wire v$G16_11911_out0;
wire v$G16_11912_out0;
wire v$G16_11913_out0;
wire v$G16_11914_out0;
wire v$G16_11915_out0;
wire v$G16_11916_out0;
wire v$G16_11917_out0;
wire v$G16_11918_out0;
wire v$G16_11919_out0;
wire v$G16_11920_out0;
wire v$G16_11921_out0;
wire v$G16_11922_out0;
wire v$G16_11923_out0;
wire v$G16_11924_out0;
wire v$G16_11925_out0;
wire v$G16_11926_out0;
wire v$G16_11927_out0;
wire v$G16_11928_out0;
wire v$G16_11929_out0;
wire v$G16_11930_out0;
wire v$G16_11931_out0;
wire v$G16_11932_out0;
wire v$G16_11933_out0;
wire v$G16_11934_out0;
wire v$G16_12037_out0;
wire v$G16_12038_out0;
wire v$G16_12044_out0;
wire v$G16_12045_out0;
wire v$G16_13408_out0;
wire v$G16_13409_out0;
wire v$G16_1783_out0;
wire v$G16_1784_out0;
wire v$G16_2222_out0;
wire v$G16_2223_out0;
wire v$G16_2547_out0;
wire v$G16_2548_out0;
wire v$G16_3103_out0;
wire v$G16_3104_out0;
wire v$G16_4405_out0;
wire v$G16_4406_out0;
wire v$G16_4419_out0;
wire v$G16_4420_out0;
wire v$G16_544_out0;
wire v$G16_545_out0;
wire v$G16_7742_out0;
wire v$G16_7743_out0;
wire v$G17_10145_out0;
wire v$G17_10146_out0;
wire v$G17_291_out0;
wire v$G17_292_out0;
wire v$G17_3706_out0;
wire v$G17_3707_out0;
wire v$G17_3720_out0;
wire v$G17_3721_out0;
wire v$G17_3764_out0;
wire v$G17_3765_out0;
wire v$G17_5670_out0;
wire v$G17_5671_out0;
wire v$G17_5672_out0;
wire v$G17_5673_out0;
wire v$G17_5674_out0;
wire v$G17_5675_out0;
wire v$G17_5676_out0;
wire v$G17_5677_out0;
wire v$G17_5678_out0;
wire v$G17_5679_out0;
wire v$G17_5680_out0;
wire v$G17_5681_out0;
wire v$G17_5682_out0;
wire v$G17_5683_out0;
wire v$G17_5684_out0;
wire v$G17_5685_out0;
wire v$G17_5686_out0;
wire v$G17_5687_out0;
wire v$G17_5688_out0;
wire v$G17_5689_out0;
wire v$G17_5690_out0;
wire v$G17_5691_out0;
wire v$G17_5692_out0;
wire v$G17_5693_out0;
wire v$G17_6070_out0;
wire v$G17_6071_out0;
wire v$G17_6145_out0;
wire v$G17_6146_out0;
wire v$G17_7508_out0;
wire v$G17_7509_out0;
wire v$G17_7915_out0;
wire v$G17_7916_out0;
wire v$G17_9354_out0;
wire v$G17_9355_out0;
wire v$G18_12843_out0;
wire v$G18_12844_out0;
wire v$G18_1749_out0;
wire v$G18_1750_out0;
wire v$G18_2105_out0;
wire v$G18_2106_out0;
wire v$G18_3366_out0;
wire v$G18_3367_out0;
wire v$G18_3368_out0;
wire v$G18_3369_out0;
wire v$G18_3370_out0;
wire v$G18_3371_out0;
wire v$G18_3372_out0;
wire v$G18_3373_out0;
wire v$G18_3374_out0;
wire v$G18_3375_out0;
wire v$G18_3376_out0;
wire v$G18_3377_out0;
wire v$G18_3378_out0;
wire v$G18_3379_out0;
wire v$G18_3380_out0;
wire v$G18_3381_out0;
wire v$G18_3382_out0;
wire v$G18_3383_out0;
wire v$G18_3384_out0;
wire v$G18_3385_out0;
wire v$G18_3386_out0;
wire v$G18_3387_out0;
wire v$G18_3388_out0;
wire v$G18_3389_out0;
wire v$G18_5076_out0;
wire v$G18_5077_out0;
wire v$G18_5876_out0;
wire v$G18_5877_out0;
wire v$G18_6825_out0;
wire v$G18_6826_out0;
wire v$G18_7271_out0;
wire v$G18_7272_out0;
wire v$G18_9091_out0;
wire v$G18_9092_out0;
wire v$G18_9163_out0;
wire v$G18_9164_out0;
wire v$G19_11088_out0;
wire v$G19_11089_out0;
wire v$G19_11146_out0;
wire v$G19_11147_out0;
wire v$G19_11223_out0;
wire v$G19_11224_out0;
wire v$G19_11762_out0;
wire v$G19_11763_out0;
wire v$G19_1347_out0;
wire v$G19_1348_out0;
wire v$G19_1593_out0;
wire v$G19_1594_out0;
wire v$G19_272_out0;
wire v$G19_273_out0;
wire v$G19_5745_out0;
wire v$G19_5746_out0;
wire v$G19_6817_out0;
wire v$G19_6818_out0;
wire v$G19_6819_out0;
wire v$G19_6820_out0;
wire v$G19_9396_out0;
wire v$G19_9397_out0;
wire v$G1_10445_out0;
wire v$G1_10446_out0;
wire v$G1_10609_out0;
wire v$G1_10610_out0;
wire v$G1_1066_out0;
wire v$G1_1067_out0;
wire v$G1_10855_out0;
wire v$G1_10856_out0;
wire v$G1_11011_out0;
wire v$G1_11012_out0;
wire v$G1_11209_out0;
wire v$G1_11210_out0;
wire v$G1_11211_out0;
wire v$G1_11212_out0;
wire v$G1_11213_out0;
wire v$G1_11214_out0;
wire v$G1_11215_out0;
wire v$G1_11216_out0;
wire v$G1_11306_out0;
wire v$G1_11307_out0;
wire v$G1_11308_out0;
wire v$G1_11309_out0;
wire v$G1_11310_out0;
wire v$G1_11311_out0;
wire v$G1_11312_out0;
wire v$G1_11313_out0;
wire v$G1_11314_out0;
wire v$G1_11315_out0;
wire v$G1_11316_out0;
wire v$G1_11317_out0;
wire v$G1_11506_out0;
wire v$G1_11507_out0;
wire v$G1_11574_out0;
wire v$G1_11575_out0;
wire v$G1_12074_out0;
wire v$G1_12075_out0;
wire v$G1_12250_out0;
wire v$G1_12251_out0;
wire v$G1_12252_out0;
wire v$G1_12253_out0;
wire v$G1_12670_out0;
wire v$G1_12671_out0;
wire v$G1_13283_out0;
wire v$G1_13284_out0;
wire v$G1_160_out0;
wire v$G1_161_out0;
wire v$G1_2894_out0;
wire v$G1_2895_out0;
wire v$G1_30_out0;
wire v$G1_31_out0;
wire v$G1_3667_out0;
wire v$G1_3668_out0;
wire v$G1_4832_out0;
wire v$G1_4833_out0;
wire v$G1_483_out0;
wire v$G1_484_out0;
wire v$G1_4923_out0;
wire v$G1_4924_out0;
wire v$G1_4931_out0;
wire v$G1_511_out0;
wire v$G1_512_out0;
wire v$G1_6037_out0;
wire v$G1_6038_out0;
wire v$G1_6039_out0;
wire v$G1_6040_out0;
wire v$G1_6387_out0;
wire v$G1_6388_out0;
wire v$G1_6389_out0;
wire v$G1_6390_out0;
wire v$G1_6391_out0;
wire v$G1_6392_out0;
wire v$G1_6393_out0;
wire v$G1_6394_out0;
wire v$G1_6877_out0;
wire v$G1_6878_out0;
wire v$G1_7899_out0;
wire v$G1_7900_out0;
wire v$G1_794_out0;
wire v$G1_795_out0;
wire v$G1_8621_out0;
wire v$G1_8622_out0;
wire v$G1_8623_out0;
wire v$G1_8760_out0;
wire v$G1_8761_out0;
wire v$G1_8792_out0;
wire v$G1_8793_out0;
wire v$G1_8794_out0;
wire v$G1_8795_out0;
wire v$G1_9116_out0;
wire v$G1_9117_out0;
wire v$G1_9792_out0;
wire v$G1_9855_out0;
wire v$G1_9856_out0;
wire v$G1_9970_out0;
wire v$G1_9971_out0;
wire v$G1_9972_out0;
wire v$G1_9973_out0;
wire v$G1_9974_out0;
wire v$G1_9975_out0;
wire v$G20_11140_out0;
wire v$G20_11141_out0;
wire v$G20_12991_out0;
wire v$G20_12992_out0;
wire v$G20_1501_out0;
wire v$G20_1502_out0;
wire v$G20_3698_out0;
wire v$G20_3699_out0;
wire v$G20_4995_out0;
wire v$G20_4996_out0;
wire v$G20_6619_out0;
wire v$G20_6620_out0;
wire v$G20_6621_out0;
wire v$G20_6622_out0;
wire v$G20_6623_out0;
wire v$G20_6624_out0;
wire v$G20_6625_out0;
wire v$G20_6626_out0;
wire v$G20_6627_out0;
wire v$G20_6628_out0;
wire v$G20_6629_out0;
wire v$G20_6630_out0;
wire v$G20_6631_out0;
wire v$G20_6632_out0;
wire v$G20_6633_out0;
wire v$G20_6634_out0;
wire v$G20_6635_out0;
wire v$G20_6636_out0;
wire v$G20_6637_out0;
wire v$G20_6638_out0;
wire v$G20_6639_out0;
wire v$G20_6640_out0;
wire v$G20_6641_out0;
wire v$G20_6642_out0;
wire v$G20_7530_out0;
wire v$G20_7531_out0;
wire v$G20_7982_out0;
wire v$G20_7983_out0;
wire v$G20_8064_out0;
wire v$G20_8065_out0;
wire v$G20_8393_out0;
wire v$G20_8394_out0;
wire v$G21_10066_out0;
wire v$G21_10067_out0;
wire v$G21_10619_out0;
wire v$G21_10620_out0;
wire v$G21_11040_out0;
wire v$G21_11041_out0;
wire v$G21_12498_out0;
wire v$G21_12499_out0;
wire v$G21_13310_out0;
wire v$G21_13311_out0;
wire v$G21_2224_out0;
wire v$G21_2225_out0;
wire v$G21_2226_out0;
wire v$G21_2227_out0;
wire v$G21_2228_out0;
wire v$G21_2229_out0;
wire v$G21_2230_out0;
wire v$G21_2231_out0;
wire v$G21_2232_out0;
wire v$G21_2233_out0;
wire v$G21_2234_out0;
wire v$G21_2235_out0;
wire v$G21_2236_out0;
wire v$G21_2237_out0;
wire v$G21_2238_out0;
wire v$G21_2239_out0;
wire v$G21_2240_out0;
wire v$G21_2241_out0;
wire v$G21_2242_out0;
wire v$G21_2243_out0;
wire v$G21_2244_out0;
wire v$G21_2245_out0;
wire v$G21_2246_out0;
wire v$G21_2247_out0;
wire v$G21_4790_out0;
wire v$G21_4791_out0;
wire v$G21_5060_out0;
wire v$G21_5061_out0;
wire v$G21_7669_out0;
wire v$G21_7670_out0;
wire v$G21_9642_out0;
wire v$G21_9643_out0;
wire v$G22_10639_out0;
wire v$G22_10640_out0;
wire v$G22_10900_out0;
wire v$G22_10901_out0;
wire v$G22_11070_out0;
wire v$G22_11071_out0;
wire v$G22_2984_out0;
wire v$G22_2985_out0;
wire v$G22_3274_out0;
wire v$G22_3275_out0;
wire v$G22_3708_out0;
wire v$G22_3709_out0;
wire v$G22_4865_out0;
wire v$G22_4866_out0;
wire v$G22_8901_out0;
wire v$G22_8902_out0;
wire v$G22_8903_out0;
wire v$G22_8904_out0;
wire v$G22_8905_out0;
wire v$G22_8906_out0;
wire v$G22_8907_out0;
wire v$G22_8908_out0;
wire v$G22_8909_out0;
wire v$G22_8910_out0;
wire v$G22_8911_out0;
wire v$G22_8912_out0;
wire v$G22_8913_out0;
wire v$G22_8914_out0;
wire v$G22_8915_out0;
wire v$G22_8916_out0;
wire v$G22_8917_out0;
wire v$G22_8918_out0;
wire v$G22_8919_out0;
wire v$G22_8920_out0;
wire v$G22_8921_out0;
wire v$G22_8922_out0;
wire v$G22_8923_out0;
wire v$G22_8924_out0;
wire v$G23_11817_out0;
wire v$G23_11818_out0;
wire v$G23_1199_out0;
wire v$G23_1200_out0;
wire v$G23_12511_out0;
wire v$G23_12512_out0;
wire v$G23_13291_out0;
wire v$G23_13292_out0;
wire v$G23_3040_out0;
wire v$G23_3041_out0;
wire v$G23_4753_out0;
wire v$G23_4754_out0;
wire v$G23_6381_out0;
wire v$G23_6382_out0;
wire v$G23_6562_out0;
wire v$G23_6563_out0;
wire v$G23_7948_out0;
wire v$G23_7949_out0;
wire v$G23_7950_out0;
wire v$G23_7951_out0;
wire v$G23_7952_out0;
wire v$G23_7953_out0;
wire v$G23_7954_out0;
wire v$G23_7955_out0;
wire v$G23_7956_out0;
wire v$G23_7957_out0;
wire v$G23_7958_out0;
wire v$G23_7959_out0;
wire v$G23_7960_out0;
wire v$G23_7961_out0;
wire v$G23_7962_out0;
wire v$G23_7963_out0;
wire v$G23_7964_out0;
wire v$G23_7965_out0;
wire v$G23_7966_out0;
wire v$G23_7967_out0;
wire v$G23_7968_out0;
wire v$G23_7969_out0;
wire v$G23_7970_out0;
wire v$G23_7971_out0;
wire v$G23_9472_out0;
wire v$G23_9473_out0;
wire v$G24_10947_out0;
wire v$G24_10948_out0;
wire v$G24_10949_out0;
wire v$G24_10950_out0;
wire v$G24_10951_out0;
wire v$G24_10952_out0;
wire v$G24_10953_out0;
wire v$G24_10954_out0;
wire v$G24_10955_out0;
wire v$G24_10956_out0;
wire v$G24_10957_out0;
wire v$G24_10958_out0;
wire v$G24_10959_out0;
wire v$G24_10960_out0;
wire v$G24_10961_out0;
wire v$G24_10962_out0;
wire v$G24_10963_out0;
wire v$G24_10964_out0;
wire v$G24_10965_out0;
wire v$G24_10966_out0;
wire v$G24_10967_out0;
wire v$G24_10968_out0;
wire v$G24_10969_out0;
wire v$G24_10970_out0;
wire v$G24_12076_out0;
wire v$G24_12077_out0;
wire v$G24_12707_out0;
wire v$G24_12708_out0;
wire v$G24_13080_out0;
wire v$G24_13081_out0;
wire v$G24_2107_out0;
wire v$G24_2108_out0;
wire v$G24_386_out0;
wire v$G24_387_out0;
wire v$G24_5412_out0;
wire v$G24_5413_out0;
wire v$G24_6574_out0;
wire v$G24_6575_out0;
wire v$G24_6893_out0;
wire v$G24_6894_out0;
wire v$G24_7868_out0;
wire v$G24_7869_out0;
wire v$G24_9384_out0;
wire v$G24_9385_out0;
wire v$G25_10025_out0;
wire v$G25_10026_out0;
wire v$G25_11283_out0;
wire v$G25_11284_out0;
wire v$G25_12841_out0;
wire v$G25_12842_out0;
wire v$G25_1387_out0;
wire v$G25_1388_out0;
wire v$G25_2250_out0;
wire v$G25_2251_out0;
wire v$G25_540_out0;
wire v$G25_541_out0;
wire v$G25_7203_out0;
wire v$G25_7204_out0;
wire v$G25_7205_out0;
wire v$G25_7206_out0;
wire v$G25_7207_out0;
wire v$G25_7208_out0;
wire v$G25_7209_out0;
wire v$G25_7210_out0;
wire v$G25_7211_out0;
wire v$G25_7212_out0;
wire v$G25_7213_out0;
wire v$G25_7214_out0;
wire v$G25_7215_out0;
wire v$G25_7216_out0;
wire v$G25_7217_out0;
wire v$G25_7218_out0;
wire v$G25_7219_out0;
wire v$G25_7220_out0;
wire v$G25_7221_out0;
wire v$G25_7222_out0;
wire v$G25_7223_out0;
wire v$G25_7224_out0;
wire v$G25_7225_out0;
wire v$G25_7226_out0;
wire v$G25_8408_out0;
wire v$G25_8409_out0;
wire v$G25_8634_out0;
wire v$G25_8635_out0;
wire v$G25_9422_out0;
wire v$G25_9423_out0;
wire v$G25_9956_out0;
wire v$G25_9957_out0;
wire v$G26_10232_out0;
wire v$G26_10233_out0;
wire v$G26_11199_out0;
wire v$G26_11200_out0;
wire v$G26_11205_out0;
wire v$G26_11206_out0;
wire v$G26_2796_out0;
wire v$G26_2797_out0;
wire v$G26_6879_out0;
wire v$G26_6880_out0;
wire v$G26_7414_out0;
wire v$G26_7415_out0;
wire v$G26_7416_out0;
wire v$G26_7417_out0;
wire v$G26_8296_out0;
wire v$G26_8297_out0;
wire v$G26_8786_out0;
wire v$G26_8787_out0;
wire v$G26_9193_out0;
wire v$G26_9194_out0;
wire v$G27_11608_out0;
wire v$G27_11609_out0;
wire v$G27_13157_out0;
wire v$G27_13158_out0;
wire v$G27_1425_out0;
wire v$G27_1426_out0;
wire v$G27_225_out0;
wire v$G27_226_out0;
wire v$G27_3185_out0;
wire v$G27_3186_out0;
wire v$G27_3187_out0;
wire v$G27_3188_out0;
wire v$G27_3189_out0;
wire v$G27_3190_out0;
wire v$G27_3191_out0;
wire v$G27_3192_out0;
wire v$G27_3193_out0;
wire v$G27_3194_out0;
wire v$G27_3195_out0;
wire v$G27_3196_out0;
wire v$G27_3197_out0;
wire v$G27_3198_out0;
wire v$G27_3199_out0;
wire v$G27_3200_out0;
wire v$G27_3201_out0;
wire v$G27_3202_out0;
wire v$G27_3203_out0;
wire v$G27_3204_out0;
wire v$G27_3205_out0;
wire v$G27_3206_out0;
wire v$G27_3207_out0;
wire v$G27_3208_out0;
wire v$G27_6811_out0;
wire v$G27_6812_out0;
wire v$G27_7526_out0;
wire v$G27_7527_out0;
wire v$G27_7528_out0;
wire v$G27_7529_out0;
wire v$G28_10029_out0;
wire v$G28_10030_out0;
wire v$G28_10676_out0;
wire v$G28_10677_out0;
wire v$G28_10902_out0;
wire v$G28_10903_out0;
wire v$G28_13203_out0;
wire v$G28_13204_out0;
wire v$G28_1895_out0;
wire v$G28_1896_out0;
wire v$G28_2473_out0;
wire v$G28_2474_out0;
wire v$G28_7110_out0;
wire v$G28_7111_out0;
wire v$G28_7730_out0;
wire v$G28_7731_out0;
wire v$G28_8638_out0;
wire v$G28_8639_out0;
wire v$G28_8640_out0;
wire v$G28_8641_out0;
wire v$G28_8642_out0;
wire v$G28_8643_out0;
wire v$G28_8644_out0;
wire v$G28_8645_out0;
wire v$G28_8646_out0;
wire v$G28_8647_out0;
wire v$G28_8648_out0;
wire v$G28_8649_out0;
wire v$G28_8650_out0;
wire v$G28_8651_out0;
wire v$G28_8652_out0;
wire v$G28_8653_out0;
wire v$G28_8654_out0;
wire v$G28_8655_out0;
wire v$G28_8656_out0;
wire v$G28_8657_out0;
wire v$G28_8658_out0;
wire v$G28_8659_out0;
wire v$G28_8660_out0;
wire v$G28_8661_out0;
wire v$G29_11007_out0;
wire v$G29_11008_out0;
wire v$G29_2332_out0;
wire v$G29_2333_out0;
wire v$G29_3728_out0;
wire v$G29_3729_out0;
wire v$G29_390_out0;
wire v$G29_391_out0;
wire v$G29_5042_out0;
wire v$G29_5043_out0;
wire v$G29_5378_out0;
wire v$G29_5379_out0;
wire v$G29_6859_out0;
wire v$G29_6860_out0;
wire v$G29_6861_out0;
wire v$G29_6862_out0;
wire v$G29_9392_out0;
wire v$G29_9393_out0;
wire v$G2_10344_out0;
wire v$G2_10345_out0;
wire v$G2_10346_out0;
wire v$G2_10347_out0;
wire v$G2_10348_out0;
wire v$G2_10349_out0;
wire v$G2_10350_out0;
wire v$G2_10351_out0;
wire v$G2_10352_out0;
wire v$G2_10353_out0;
wire v$G2_10354_out0;
wire v$G2_10355_out0;
wire v$G2_1044_out0;
wire v$G2_1045_out0;
wire v$G2_10819_out0;
wire v$G2_10820_out0;
wire v$G2_10999_out0;
wire v$G2_11000_out0;
wire v$G2_11082_out0;
wire v$G2_11083_out0;
wire v$G2_11580_out0;
wire v$G2_11581_out0;
wire v$G2_12108_out0;
wire v$G2_12109_out0;
wire v$G2_12220_out0;
wire v$G2_12221_out0;
wire v$G2_12222_out0;
wire v$G2_12223_out0;
wire v$G2_12224_out0;
wire v$G2_12225_out0;
wire v$G2_12226_out0;
wire v$G2_12227_out0;
wire v$G2_12489_out0;
wire v$G2_12490_out0;
wire v$G2_12962_out0;
wire v$G2_12963_out0;
wire v$G2_12964_out0;
wire v$G2_12965_out0;
wire v$G2_13111_out0;
wire v$G2_13112_out0;
wire v$G2_13322_out0;
wire v$G2_13323_out0;
wire v$G2_1355_out0;
wire v$G2_1356_out0;
wire v$G2_2437_out0;
wire v$G2_2438_out0;
wire v$G2_2792_out0;
wire v$G2_2793_out0;
wire v$G2_3435_out0;
wire v$G2_3436_out0;
wire v$G2_3619_out0;
wire v$G2_3620_out0;
wire v$G2_3675_out0;
wire v$G2_3676_out0;
wire v$G2_5108_out0;
wire v$G2_5115_out0;
wire v$G2_5116_out0;
wire v$G2_5117_out0;
wire v$G2_529_out0;
wire v$G2_530_out0;
wire v$G2_5310_out0;
wire v$G2_5311_out0;
wire v$G2_5639_out0;
wire v$G2_5802_out0;
wire v$G2_5803_out0;
wire v$G2_62_out0;
wire v$G2_6316_out0;
wire v$G2_6317_out0;
wire v$G2_63_out0;
wire v$G2_6949_out0;
wire v$G2_6950_out0;
wire v$G2_6951_out0;
wire v$G2_6952_out0;
wire v$G2_7517_out0;
wire v$G2_7692_out0;
wire v$G2_7693_out0;
wire v$G2_7694_out0;
wire v$G2_7695_out0;
wire v$G2_8548_out0;
wire v$G2_8549_out0;
wire v$G2_8550_out0;
wire v$G2_8551_out0;
wire v$G2_8552_out0;
wire v$G2_8553_out0;
wire v$G2_8554_out0;
wire v$G2_8555_out0;
wire v$G2_9239_out0;
wire v$G2_9240_out0;
wire v$G2_9887_out0;
wire v$G2_9888_out0;
wire v$G30_11118_out0;
wire v$G30_11119_out0;
wire v$G30_13247_out0;
wire v$G30_13248_out0;
wire v$G30_1389_out0;
wire v$G30_1390_out0;
wire v$G30_3316_out0;
wire v$G30_3317_out0;
wire v$G30_897_out0;
wire v$G30_898_out0;
wire v$G30_948_out0;
wire v$G30_949_out0;
wire v$G30_950_out0;
wire v$G30_951_out0;
wire v$G30_952_out0;
wire v$G30_953_out0;
wire v$G30_954_out0;
wire v$G30_955_out0;
wire v$G30_956_out0;
wire v$G30_957_out0;
wire v$G30_958_out0;
wire v$G30_959_out0;
wire v$G30_960_out0;
wire v$G30_961_out0;
wire v$G30_962_out0;
wire v$G30_963_out0;
wire v$G30_964_out0;
wire v$G30_965_out0;
wire v$G30_966_out0;
wire v$G30_967_out0;
wire v$G30_968_out0;
wire v$G30_969_out0;
wire v$G30_970_out0;
wire v$G30_971_out0;
wire v$G31_10787_out0;
wire v$G31_10788_out0;
wire v$G31_10789_out0;
wire v$G31_10790_out0;
wire v$G31_10791_out0;
wire v$G31_10792_out0;
wire v$G31_10793_out0;
wire v$G31_10794_out0;
wire v$G31_10795_out0;
wire v$G31_10796_out0;
wire v$G31_10797_out0;
wire v$G31_10798_out0;
wire v$G31_10799_out0;
wire v$G31_10800_out0;
wire v$G31_10801_out0;
wire v$G31_10802_out0;
wire v$G31_10803_out0;
wire v$G31_10804_out0;
wire v$G31_10805_out0;
wire v$G31_10806_out0;
wire v$G31_10807_out0;
wire v$G31_10808_out0;
wire v$G31_10809_out0;
wire v$G31_10810_out0;
wire v$G31_13271_out0;
wire v$G31_13272_out0;
wire v$G31_6588_out0;
wire v$G31_6589_out0;
wire v$G31_7100_out0;
wire v$G31_7101_out0;
wire v$G31_997_out0;
wire v$G31_998_out0;
wire v$G32_1001_out0;
wire v$G32_1002_out0;
wire v$G32_11448_out0;
wire v$G32_11449_out0;
wire v$G32_11512_out0;
wire v$G32_11513_out0;
wire v$G32_321_out0;
wire v$G32_322_out0;
wire v$G32_323_out0;
wire v$G32_324_out0;
wire v$G32_325_out0;
wire v$G32_326_out0;
wire v$G32_327_out0;
wire v$G32_328_out0;
wire v$G32_329_out0;
wire v$G32_330_out0;
wire v$G32_331_out0;
wire v$G32_332_out0;
wire v$G32_333_out0;
wire v$G32_334_out0;
wire v$G32_335_out0;
wire v$G32_336_out0;
wire v$G32_337_out0;
wire v$G32_338_out0;
wire v$G32_339_out0;
wire v$G32_340_out0;
wire v$G32_341_out0;
wire v$G32_342_out0;
wire v$G32_343_out0;
wire v$G32_344_out0;
wire v$G32_6353_out0;
wire v$G32_6354_out0;
wire v$G32_7679_out0;
wire v$G32_7680_out0;
wire v$G33_3506_out0;
wire v$G33_3507_out0;
wire v$G33_502_out0;
wire v$G33_503_out0;
wire v$G33_7075_out0;
wire v$G33_7076_out0;
wire v$G33_8722_out0;
wire v$G33_8723_out0;
wire v$G33_8724_out0;
wire v$G33_8725_out0;
wire v$G33_8726_out0;
wire v$G33_8727_out0;
wire v$G33_8728_out0;
wire v$G33_8729_out0;
wire v$G33_8730_out0;
wire v$G33_8731_out0;
wire v$G33_8732_out0;
wire v$G33_8733_out0;
wire v$G33_8734_out0;
wire v$G33_8735_out0;
wire v$G33_8736_out0;
wire v$G33_8737_out0;
wire v$G33_8738_out0;
wire v$G33_8739_out0;
wire v$G33_8740_out0;
wire v$G33_8741_out0;
wire v$G33_8742_out0;
wire v$G33_8743_out0;
wire v$G33_8744_out0;
wire v$G33_8745_out0;
wire v$G34_12121_out0;
wire v$G34_12122_out0;
wire v$G34_12123_out0;
wire v$G34_12124_out0;
wire v$G34_12125_out0;
wire v$G34_12126_out0;
wire v$G34_12127_out0;
wire v$G34_12128_out0;
wire v$G34_12129_out0;
wire v$G34_12130_out0;
wire v$G34_12131_out0;
wire v$G34_12132_out0;
wire v$G34_12133_out0;
wire v$G34_12134_out0;
wire v$G34_12135_out0;
wire v$G34_12136_out0;
wire v$G34_12137_out0;
wire v$G34_12138_out0;
wire v$G34_12139_out0;
wire v$G34_12140_out0;
wire v$G34_12141_out0;
wire v$G34_12142_out0;
wire v$G34_12143_out0;
wire v$G34_12144_out0;
wire v$G34_3310_out0;
wire v$G34_3311_out0;
wire v$G34_777_out0;
wire v$G34_778_out0;
wire v$G35_2986_out0;
wire v$G35_2987_out0;
wire v$G35_445_out0;
wire v$G35_446_out0;
wire v$G35_6881_out0;
wire v$G35_6882_out0;
wire v$G35_8276_out0;
wire v$G35_8277_out0;
wire v$G35_9911_out0;
wire v$G35_9912_out0;
wire v$G35_9913_out0;
wire v$G35_9914_out0;
wire v$G35_9915_out0;
wire v$G35_9916_out0;
wire v$G35_9917_out0;
wire v$G35_9918_out0;
wire v$G35_9919_out0;
wire v$G35_9920_out0;
wire v$G35_9921_out0;
wire v$G35_9922_out0;
wire v$G35_9923_out0;
wire v$G35_9924_out0;
wire v$G35_9925_out0;
wire v$G35_9926_out0;
wire v$G35_9927_out0;
wire v$G35_9928_out0;
wire v$G35_9929_out0;
wire v$G35_9930_out0;
wire v$G35_9931_out0;
wire v$G35_9932_out0;
wire v$G35_9933_out0;
wire v$G35_9934_out0;
wire v$G36_11766_out0;
wire v$G36_12163_out0;
wire v$G36_12164_out0;
wire v$G36_3923_out0;
wire v$G36_3924_out0;
wire v$G36_3925_out0;
wire v$G36_3926_out0;
wire v$G36_3927_out0;
wire v$G36_3928_out0;
wire v$G36_3929_out0;
wire v$G36_3930_out0;
wire v$G36_3931_out0;
wire v$G36_3932_out0;
wire v$G36_3933_out0;
wire v$G36_3934_out0;
wire v$G36_3935_out0;
wire v$G36_3936_out0;
wire v$G36_3937_out0;
wire v$G36_3938_out0;
wire v$G36_3939_out0;
wire v$G36_3940_out0;
wire v$G36_3941_out0;
wire v$G36_3942_out0;
wire v$G36_3943_out0;
wire v$G36_3944_out0;
wire v$G36_3945_out0;
wire v$G36_3946_out0;
wire v$G36_7154_out0;
wire v$G36_7155_out0;
wire v$G36_9492_out0;
wire v$G36_9493_out0;
wire v$G37_13137_out0;
wire v$G37_13138_out0;
wire v$G37_394_out0;
wire v$G37_395_out0;
wire v$G37_585_out0;
wire v$G37_586_out0;
wire v$G37_743_out0;
wire v$G37_744_out0;
wire v$G37_745_out0;
wire v$G37_746_out0;
wire v$G38_4889_out0;
wire v$G38_4890_out0;
wire v$G38_4891_out0;
wire v$G38_4892_out0;
wire v$G38_4893_out0;
wire v$G38_4894_out0;
wire v$G38_4895_out0;
wire v$G38_4896_out0;
wire v$G38_4897_out0;
wire v$G38_4898_out0;
wire v$G38_4899_out0;
wire v$G38_4900_out0;
wire v$G38_4901_out0;
wire v$G38_4902_out0;
wire v$G38_4903_out0;
wire v$G38_4904_out0;
wire v$G38_4905_out0;
wire v$G38_4906_out0;
wire v$G38_4907_out0;
wire v$G38_4908_out0;
wire v$G38_4909_out0;
wire v$G38_4910_out0;
wire v$G38_4911_out0;
wire v$G38_4912_out0;
wire v$G38_6823_out0;
wire v$G38_6824_out0;
wire v$G39_11939_out0;
wire v$G39_11940_out0;
wire v$G39_12167_out0;
wire v$G39_12168_out0;
wire v$G39_12169_out0;
wire v$G39_12170_out0;
wire v$G39_4047_out0;
wire v$G39_4048_out0;
wire v$G3_0_out0;
wire v$G3_11055_out0;
wire v$G3_11056_out0;
wire v$G3_11192_out0;
wire v$G3_11193_out0;
wire v$G3_11270_out0;
wire v$G3_12256_out0;
wire v$G3_12257_out0;
wire v$G3_12513_out0;
wire v$G3_12514_out0;
wire v$G3_12515_out0;
wire v$G3_13101_out0;
wire v$G3_13102_out0;
wire v$G3_1369_out0;
wire v$G3_1370_out0;
wire v$G3_1507_out0;
wire v$G3_1508_out0;
wire v$G3_1509_out0;
wire v$G3_1510_out0;
wire v$G3_1511_out0;
wire v$G3_1512_out0;
wire v$G3_1513_out0;
wire v$G3_1514_out0;
wire v$G3_1573_out0;
wire v$G3_1574_out0;
wire v$G3_1738_out0;
wire v$G3_1_out0;
wire v$G3_22_out0;
wire v$G3_23_out0;
wire v$G3_2658_out0;
wire v$G3_2659_out0;
wire v$G3_2662_out0;
wire v$G3_2663_out0;
wire v$G3_2802_out0;
wire v$G3_2803_out0;
wire v$G3_3149_out0;
wire v$G3_3150_out0;
wire v$G3_3394_out0;
wire v$G3_5062_out0;
wire v$G3_5063_out0;
wire v$G3_5064_out0;
wire v$G3_5065_out0;
wire v$G3_5080_out0;
wire v$G3_5081_out0;
wire v$G3_5136_out0;
wire v$G3_5137_out0;
wire v$G3_5549_out0;
wire v$G3_5550_out0;
wire v$G3_6059_out0;
wire v$G3_6060_out0;
wire v$G3_6061_out0;
wire v$G3_6062_out0;
wire v$G3_6063_out0;
wire v$G3_6064_out0;
wire v$G3_6065_out0;
wire v$G3_6066_out0;
wire v$G3_6067_out0;
wire v$G3_6068_out0;
wire v$G3_6377_out0;
wire v$G3_6378_out0;
wire v$G3_6429_out0;
wire v$G3_6430_out0;
wire v$G3_6660_out0;
wire v$G3_6661_out0;
wire v$G3_6809_out0;
wire v$G3_6810_out0;
wire v$G3_7242_out0;
wire v$G3_7243_out0;
wire v$G3_8305_out0;
wire v$G3_8306_out0;
wire v$G3_8307_out0;
wire v$G3_8308_out0;
wire v$G3_8309_out0;
wire v$G3_8310_out0;
wire v$G3_8311_out0;
wire v$G3_8312_out0;
wire v$G3_8313_out0;
wire v$G3_8314_out0;
wire v$G3_8315_out0;
wire v$G3_8316_out0;
wire v$G3_8317_out0;
wire v$G3_8318_out0;
wire v$G3_8319_out0;
wire v$G3_8320_out0;
wire v$G3_8321_out0;
wire v$G3_8322_out0;
wire v$G3_8323_out0;
wire v$G3_8324_out0;
wire v$G3_8325_out0;
wire v$G3_8326_out0;
wire v$G3_8327_out0;
wire v$G3_8328_out0;
wire v$G3_8329_out0;
wire v$G3_8330_out0;
wire v$G3_8331_out0;
wire v$G3_8332_out0;
wire v$G3_8333_out0;
wire v$G3_8334_out0;
wire v$G3_8335_out0;
wire v$G3_8336_out0;
wire v$G3_8337_out0;
wire v$G3_8338_out0;
wire v$G3_8339_out0;
wire v$G3_8340_out0;
wire v$G3_8341_out0;
wire v$G3_8342_out0;
wire v$G3_8343_out0;
wire v$G3_8344_out0;
wire v$G3_8345_out0;
wire v$G3_8346_out0;
wire v$G3_8347_out0;
wire v$G3_8348_out0;
wire v$G3_8349_out0;
wire v$G3_8350_out0;
wire v$G3_8351_out0;
wire v$G3_8352_out0;
wire v$G3_8353_out0;
wire v$G3_8354_out0;
wire v$G3_8355_out0;
wire v$G3_8356_out0;
wire v$G3_8357_out0;
wire v$G3_8358_out0;
wire v$G3_8359_out0;
wire v$G3_8360_out0;
wire v$G3_8361_out0;
wire v$G3_8362_out0;
wire v$G3_8363_out0;
wire v$G3_8364_out0;
wire v$G3_8587_out0;
wire v$G3_8588_out0;
wire v$G3_8684_out0;
wire v$G3_8685_out0;
wire v$G3_8686_out0;
wire v$G3_8687_out0;
wire v$G3_9569_out0;
wire v$G3_9570_out0;
wire v$G40_10438_out0;
wire v$G40_10439_out0;
wire v$G40_8934_out0;
wire v$G40_8935_out0;
wire v$G40_8936_out0;
wire v$G40_8937_out0;
wire v$G40_8938_out0;
wire v$G40_8939_out0;
wire v$G40_8940_out0;
wire v$G40_8941_out0;
wire v$G40_8942_out0;
wire v$G40_8943_out0;
wire v$G40_8944_out0;
wire v$G40_8945_out0;
wire v$G40_8946_out0;
wire v$G40_8947_out0;
wire v$G40_8948_out0;
wire v$G40_8949_out0;
wire v$G40_8950_out0;
wire v$G40_8951_out0;
wire v$G40_8952_out0;
wire v$G40_8953_out0;
wire v$G40_8954_out0;
wire v$G40_8955_out0;
wire v$G40_8956_out0;
wire v$G40_8957_out0;
wire v$G40_9224_out0;
wire v$G40_9225_out0;
wire v$G41_13147_out0;
wire v$G41_13148_out0;
wire v$G41_7156_out0;
wire v$G41_7157_out0;
wire v$G41_7158_out0;
wire v$G41_7159_out0;
wire v$G41_7160_out0;
wire v$G41_7161_out0;
wire v$G41_7162_out0;
wire v$G41_7163_out0;
wire v$G41_7164_out0;
wire v$G41_7165_out0;
wire v$G41_7166_out0;
wire v$G41_7167_out0;
wire v$G41_7168_out0;
wire v$G41_7169_out0;
wire v$G41_7170_out0;
wire v$G41_7171_out0;
wire v$G41_7172_out0;
wire v$G41_7173_out0;
wire v$G41_7174_out0;
wire v$G41_7175_out0;
wire v$G41_7176_out0;
wire v$G41_7177_out0;
wire v$G41_7178_out0;
wire v$G41_7179_out0;
wire v$G42_13143_out0;
wire v$G42_13144_out0;
wire v$G42_6544_out0;
wire v$G42_6545_out0;
wire v$G43_319_out0;
wire v$G43_320_out0;
wire v$G43_4800_out0;
wire v$G43_4801_out0;
wire v$G44_5734_out0;
wire v$G45_10651_out0;
wire v$G45_11949_out0;
wire v$G45_11950_out0;
wire v$G46_11285_out0;
wire v$G46_11286_out0;
wire v$G46_7181_out0;
wire v$G46_7182_out0;
wire v$G47_3665_out0;
wire v$G47_3666_out0;
wire v$G47_753_out0;
wire v$G47_754_out0;
wire v$G48_1203_out0;
wire v$G48_1204_out0;
wire v$G48_13173_out0;
wire v$G48_13174_out0;
wire v$G48_3270_out0;
wire v$G48_3271_out0;
wire v$G49_3615_out0;
wire v$G49_3616_out0;
wire v$G49_6992_out0;
wire v$G49_6993_out0;
wire v$G49_7290_out0;
wire v$G49_7291_out0;
wire v$G4_10044_out0;
wire v$G4_10045_out0;
wire v$G4_10436_out0;
wire v$G4_10437_out0;
wire v$G4_10637_out0;
wire v$G4_10638_out0;
wire v$G4_10750_out0;
wire v$G4_10751_out0;
wire v$G4_10821_out0;
wire v$G4_10822_out0;
wire v$G4_11042_out0;
wire v$G4_11043_out0;
wire v$G4_12318_out0;
wire v$G4_12319_out0;
wire v$G4_12320_out0;
wire v$G4_12321_out0;
wire v$G4_12322_out0;
wire v$G4_12323_out0;
wire v$G4_12324_out0;
wire v$G4_12325_out0;
wire v$G4_12326_out0;
wire v$G4_12327_out0;
wire v$G4_12328_out0;
wire v$G4_12329_out0;
wire v$G4_12330_out0;
wire v$G4_12331_out0;
wire v$G4_12332_out0;
wire v$G4_12333_out0;
wire v$G4_12334_out0;
wire v$G4_12335_out0;
wire v$G4_12336_out0;
wire v$G4_12337_out0;
wire v$G4_12338_out0;
wire v$G4_12339_out0;
wire v$G4_12340_out0;
wire v$G4_12341_out0;
wire v$G4_12342_out0;
wire v$G4_12343_out0;
wire v$G4_12344_out0;
wire v$G4_12345_out0;
wire v$G4_12346_out0;
wire v$G4_12347_out0;
wire v$G4_12348_out0;
wire v$G4_12349_out0;
wire v$G4_12350_out0;
wire v$G4_12351_out0;
wire v$G4_12352_out0;
wire v$G4_12353_out0;
wire v$G4_12354_out0;
wire v$G4_12355_out0;
wire v$G4_12356_out0;
wire v$G4_12357_out0;
wire v$G4_12358_out0;
wire v$G4_12359_out0;
wire v$G4_12360_out0;
wire v$G4_12361_out0;
wire v$G4_12362_out0;
wire v$G4_12363_out0;
wire v$G4_12364_out0;
wire v$G4_12365_out0;
wire v$G4_12366_out0;
wire v$G4_12367_out0;
wire v$G4_12368_out0;
wire v$G4_12369_out0;
wire v$G4_12370_out0;
wire v$G4_12371_out0;
wire v$G4_12372_out0;
wire v$G4_12373_out0;
wire v$G4_12374_out0;
wire v$G4_12375_out0;
wire v$G4_12376_out0;
wire v$G4_12377_out0;
wire v$G4_12393_out0;
wire v$G4_12394_out0;
wire v$G4_12987_out0;
wire v$G4_12988_out0;
wire v$G4_1665_out0;
wire v$G4_1666_out0;
wire v$G4_2746_out0;
wire v$G4_2747_out0;
wire v$G4_2748_out0;
wire v$G4_2749_out0;
wire v$G4_2750_out0;
wire v$G4_2751_out0;
wire v$G4_2752_out0;
wire v$G4_2753_out0;
wire v$G4_3292_out0;
wire v$G4_3293_out0;
wire v$G4_4055_out0;
wire v$G4_4056_out0;
wire v$G4_4057_out0;
wire v$G4_4058_out0;
wire v$G4_4059_out0;
wire v$G4_4060_out0;
wire v$G4_4061_out0;
wire v$G4_4062_out0;
wire v$G4_4063_out0;
wire v$G4_4064_out0;
wire v$G4_4065_out0;
wire v$G4_4066_out0;
wire v$G4_4429_out0;
wire v$G4_5100_out0;
wire v$G4_5101_out0;
wire v$G4_5283_out0;
wire v$G4_5284_out0;
wire v$G4_559_out0;
wire v$G4_560_out0;
wire v$G4_7633_out0;
wire v$G4_7634_out0;
wire v$G4_7635_out0;
wire v$G4_7636_out0;
wire v$G4_7637_out0;
wire v$G4_7638_out0;
wire v$G4_7639_out0;
wire v$G4_7640_out0;
wire v$G4_7641_out0;
wire v$G4_7642_out0;
wire v$G4_7665_out0;
wire v$G4_7666_out0;
wire v$G4_7760_out0;
wire v$G4_7761_out0;
wire v$G4_8791_out0;
wire v$G4_9398_out0;
wire v$G4_9399_out0;
wire v$G4_9611_out0;
wire v$G4_9612_out0;
wire v$G4_9889_out0;
wire v$G4_9890_out0;
wire v$G50_11471_out0;
wire v$G50_11472_out0;
wire v$G50_12147_out0;
wire v$G50_12148_out0;
wire v$G50_8804_out0;
wire v$G50_8805_out0;
wire v$G50_8876_out0;
wire v$G51_13389_out0;
wire v$G51_1633_out0;
wire v$G51_1634_out0;
wire v$G51_2159_out0;
wire v$G51_2160_out0;
wire v$G51_9413_out0;
wire v$G51_9414_out0;
wire v$G52_11142_out0;
wire v$G52_11143_out0;
wire v$G52_1732_out0;
wire v$G52_1733_out0;
wire v$G52_5403_out0;
wire v$G53_11048_out0;
wire v$G53_11049_out0;
wire v$G53_12287_out0;
wire v$G53_8369_out0;
wire v$G53_8370_out0;
wire v$G54_1052_out0;
wire v$G54_1053_out0;
wire v$G54_5642_out0;
wire v$G54_5643_out0;
wire v$G54_8868_out0;
wire v$G54_9597_out0;
wire v$G54_9598_out0;
wire v$G55_11730_out0;
wire v$G55_11731_out0;
wire v$G55_12935_out0;
wire v$G55_12936_out0;
wire v$G55_3437_out0;
wire v$G55_3438_out0;
wire v$G55_9243_out0;
wire v$G56_12500_out0;
wire v$G56_1877_out0;
wire v$G56_1878_out0;
wire v$G56_372_out0;
wire v$G56_373_out0;
wire v$G57_12731_out0;
wire v$G57_6225_out0;
wire v$G57_6226_out0;
wire v$G57_7492_out0;
wire v$G57_7493_out0;
wire v$G57_9018_out0;
wire v$G57_9019_out0;
wire v$G58_1431_out0;
wire v$G58_1432_out0;
wire v$G58_162_out0;
wire v$G58_163_out0;
wire v$G58_4796_out0;
wire v$G58_4797_out0;
wire v$G59_10432_out0;
wire v$G59_10433_out0;
wire v$G59_1484_out0;
wire v$G59_2552_out0;
wire v$G59_2553_out0;
wire v$G5_10018_out0;
wire v$G5_10019_out0;
wire v$G5_10022_out0;
wire v$G5_10023_out0;
wire v$G5_10553_out0;
wire v$G5_10554_out0;
wire v$G5_11019_out0;
wire v$G5_11020_out0;
wire v$G5_11287_out0;
wire v$G5_11288_out0;
wire v$G5_11318_out0;
wire v$G5_11319_out0;
wire v$G5_1162_out0;
wire v$G5_11636_out0;
wire v$G5_11637_out0;
wire v$G5_1163_out0;
wire v$G5_12296_out0;
wire v$G5_12297_out0;
wire v$G5_12298_out0;
wire v$G5_12299_out0;
wire v$G5_12300_out0;
wire v$G5_12301_out0;
wire v$G5_12302_out0;
wire v$G5_12303_out0;
wire v$G5_12304_out0;
wire v$G5_12305_out0;
wire v$G5_12306_out0;
wire v$G5_12307_out0;
wire v$G5_12662_out0;
wire v$G5_12663_out0;
wire v$G5_1570_out0;
wire v$G5_3817_out0;
wire v$G5_3846_out0;
wire v$G5_3847_out0;
wire v$G5_3848_out0;
wire v$G5_3849_out0;
wire v$G5_3850_out0;
wire v$G5_3851_out0;
wire v$G5_3852_out0;
wire v$G5_3853_out0;
wire v$G5_3854_out0;
wire v$G5_3855_out0;
wire v$G5_3856_out0;
wire v$G5_3857_out0;
wire v$G5_3858_out0;
wire v$G5_3859_out0;
wire v$G5_3860_out0;
wire v$G5_3861_out0;
wire v$G5_3862_out0;
wire v$G5_3863_out0;
wire v$G5_3864_out0;
wire v$G5_3865_out0;
wire v$G5_3866_out0;
wire v$G5_3867_out0;
wire v$G5_3868_out0;
wire v$G5_3869_out0;
wire v$G5_3870_out0;
wire v$G5_3871_out0;
wire v$G5_3872_out0;
wire v$G5_3873_out0;
wire v$G5_3874_out0;
wire v$G5_3875_out0;
wire v$G5_3876_out0;
wire v$G5_3877_out0;
wire v$G5_3878_out0;
wire v$G5_3879_out0;
wire v$G5_3880_out0;
wire v$G5_3881_out0;
wire v$G5_3882_out0;
wire v$G5_3883_out0;
wire v$G5_3884_out0;
wire v$G5_3885_out0;
wire v$G5_3886_out0;
wire v$G5_3887_out0;
wire v$G5_3888_out0;
wire v$G5_3889_out0;
wire v$G5_3890_out0;
wire v$G5_3891_out0;
wire v$G5_3892_out0;
wire v$G5_3893_out0;
wire v$G5_3894_out0;
wire v$G5_3895_out0;
wire v$G5_3896_out0;
wire v$G5_3897_out0;
wire v$G5_3898_out0;
wire v$G5_3899_out0;
wire v$G5_3900_out0;
wire v$G5_3901_out0;
wire v$G5_3902_out0;
wire v$G5_3903_out0;
wire v$G5_3904_out0;
wire v$G5_3905_out0;
wire v$G5_4215_out0;
wire v$G5_4216_out0;
wire v$G5_423_out0;
wire v$G5_424_out0;
wire v$G5_425_out0;
wire v$G5_426_out0;
wire v$G5_427_out0;
wire v$G5_428_out0;
wire v$G5_429_out0;
wire v$G5_430_out0;
wire v$G5_431_out0;
wire v$G5_432_out0;
wire v$G5_4704_out0;
wire v$G5_4705_out0;
wire v$G5_4706_out0;
wire v$G5_4707_out0;
wire v$G5_4708_out0;
wire v$G5_4709_out0;
wire v$G5_4710_out0;
wire v$G5_4711_out0;
wire v$G5_4712_out0;
wire v$G5_4713_out0;
wire v$G5_4714_out0;
wire v$G5_4715_out0;
wire v$G5_4716_out0;
wire v$G5_4717_out0;
wire v$G5_4718_out0;
wire v$G5_4719_out0;
wire v$G5_4720_out0;
wire v$G5_4721_out0;
wire v$G5_4722_out0;
wire v$G5_4723_out0;
wire v$G5_4724_out0;
wire v$G5_4725_out0;
wire v$G5_4726_out0;
wire v$G5_4727_out0;
wire v$G5_5122_out0;
wire v$G5_5123_out0;
wire v$G5_5904_out0;
wire v$G5_5905_out0;
wire v$G5_7012_out0;
wire v$G5_7013_out0;
wire v$G5_8400_out0;
wire v$G5_8401_out0;
wire v$G5_9119_out0;
wire v$G5_9120_out0;
wire v$G60_13385_out0;
wire v$G60_13386_out0;
wire v$G60_6463_out0;
wire v$G60_6464_out0;
wire v$G61_11531_out0;
wire v$G61_11532_out0;
wire v$G61_5755_out0;
wire v$G61_5756_out0;
wire v$G61_7438_out0;
wire v$G61_7439_out0;
wire v$G62_10313_out0;
wire v$G62_10314_out0;
wire v$G62_7570_out0;
wire v$G62_7571_out0;
wire v$G62_7744_out0;
wire v$G63_11847_out0;
wire v$G63_11848_out0;
wire v$G63_6734_out0;
wire v$G63_6735_out0;
wire v$G63_9223_out0;
wire v$G64_10577_out0;
wire v$G64_10578_out0;
wire v$G64_4407_out0;
wire v$G64_4408_out0;
wire v$G64_4444_out0;
wire v$G64_5316_out0;
wire v$G64_5317_out0;
wire v$G65_12942_out0;
wire v$G65_12943_out0;
wire v$G65_1383_out0;
wire v$G65_1384_out0;
wire v$G65_6054_out0;
wire v$G65_9509_out0;
wire v$G65_9510_out0;
wire v$G66_10587_out0;
wire v$G66_10588_out0;
wire v$G66_11892_out0;
wire v$G66_11893_out0;
wire v$G66_5924_out0;
wire v$G66_5925_out0;
wire v$G66_6177_out0;
wire v$G67_7297_out0;
wire v$G67_7298_out0;
wire v$G67_9285_out0;
wire v$G67_9496_out0;
wire v$G67_9497_out0;
wire v$G68_10170_out0;
wire v$G68_10489_out0;
wire v$G68_10490_out0;
wire v$G68_12849_out0;
wire v$G68_12850_out0;
wire v$G69_11035_out0;
wire v$G69_489_out0;
wire v$G69_490_out0;
wire v$G69_5702_out0;
wire v$G69_5703_out0;
wire v$G6_10833_out0;
wire v$G6_10834_out0;
wire v$G6_10835_out0;
wire v$G6_10836_out0;
wire v$G6_10837_out0;
wire v$G6_10838_out0;
wire v$G6_10839_out0;
wire v$G6_10840_out0;
wire v$G6_10841_out0;
wire v$G6_10842_out0;
wire v$G6_10843_out0;
wire v$G6_10844_out0;
wire v$G6_10845_out0;
wire v$G6_10846_out0;
wire v$G6_10847_out0;
wire v$G6_10848_out0;
wire v$G6_10849_out0;
wire v$G6_10850_out0;
wire v$G6_10851_out0;
wire v$G6_10852_out0;
wire v$G6_10853_out0;
wire v$G6_10854_out0;
wire v$G6_1174_out0;
wire v$G6_1175_out0;
wire v$G6_11846_out0;
wire v$G6_12207_out0;
wire v$G6_1891_out0;
wire v$G6_1892_out0;
wire v$G6_2050_out0;
wire v$G6_2051_out0;
wire v$G6_2205_out0;
wire v$G6_2256_out0;
wire v$G6_2257_out0;
wire v$G6_2258_out0;
wire v$G6_2259_out0;
wire v$G6_2260_out0;
wire v$G6_2261_out0;
wire v$G6_2262_out0;
wire v$G6_2263_out0;
wire v$G6_2264_out0;
wire v$G6_2265_out0;
wire v$G6_2266_out0;
wire v$G6_2267_out0;
wire v$G6_2268_out0;
wire v$G6_2269_out0;
wire v$G6_2270_out0;
wire v$G6_2271_out0;
wire v$G6_2272_out0;
wire v$G6_2273_out0;
wire v$G6_2274_out0;
wire v$G6_2275_out0;
wire v$G6_2276_out0;
wire v$G6_2277_out0;
wire v$G6_2278_out0;
wire v$G6_2279_out0;
wire v$G6_2280_out0;
wire v$G6_2281_out0;
wire v$G6_2282_out0;
wire v$G6_2283_out0;
wire v$G6_2284_out0;
wire v$G6_2285_out0;
wire v$G6_2286_out0;
wire v$G6_2287_out0;
wire v$G6_2288_out0;
wire v$G6_2289_out0;
wire v$G6_2290_out0;
wire v$G6_2291_out0;
wire v$G6_2292_out0;
wire v$G6_2293_out0;
wire v$G6_2294_out0;
wire v$G6_2295_out0;
wire v$G6_2296_out0;
wire v$G6_2297_out0;
wire v$G6_2298_out0;
wire v$G6_2299_out0;
wire v$G6_2300_out0;
wire v$G6_2301_out0;
wire v$G6_2302_out0;
wire v$G6_2303_out0;
wire v$G6_2304_out0;
wire v$G6_2305_out0;
wire v$G6_2306_out0;
wire v$G6_2307_out0;
wire v$G6_2308_out0;
wire v$G6_2309_out0;
wire v$G6_2310_out0;
wire v$G6_2311_out0;
wire v$G6_2312_out0;
wire v$G6_2313_out0;
wire v$G6_2314_out0;
wire v$G6_2315_out0;
wire v$G6_231_out0;
wire v$G6_232_out0;
wire v$G6_3710_out0;
wire v$G6_3711_out0;
wire v$G6_382_out0;
wire v$G6_383_out0;
wire v$G6_3951_out0;
wire v$G6_3952_out0;
wire v$G6_4177_out0;
wire v$G6_4178_out0;
wire v$G6_4183_out0;
wire v$G6_4184_out0;
wire v$G6_4185_out0;
wire v$G6_4186_out0;
wire v$G6_4187_out0;
wire v$G6_4188_out0;
wire v$G6_4189_out0;
wire v$G6_4190_out0;
wire v$G6_4191_out0;
wire v$G6_4192_out0;
wire v$G6_4193_out0;
wire v$G6_4194_out0;
wire v$G6_4195_out0;
wire v$G6_4196_out0;
wire v$G6_4197_out0;
wire v$G6_4198_out0;
wire v$G6_4554_out0;
wire v$G6_4555_out0;
wire v$G6_4556_out0;
wire v$G6_4557_out0;
wire v$G6_4558_out0;
wire v$G6_4559_out0;
wire v$G6_4560_out0;
wire v$G6_4561_out0;
wire v$G6_4562_out0;
wire v$G6_4563_out0;
wire v$G6_4564_out0;
wire v$G6_4565_out0;
wire v$G6_4566_out0;
wire v$G6_4567_out0;
wire v$G6_4568_out0;
wire v$G6_4569_out0;
wire v$G6_4570_out0;
wire v$G6_4571_out0;
wire v$G6_4572_out0;
wire v$G6_4573_out0;
wire v$G6_4574_out0;
wire v$G6_4575_out0;
wire v$G6_4576_out0;
wire v$G6_4577_out0;
wire v$G6_5056_out0;
wire v$G6_5057_out0;
wire v$G6_5440_out0;
wire v$G6_5441_out0;
wire v$G6_6314_out0;
wire v$G6_6315_out0;
wire v$G6_7724_out0;
wire v$G6_7725_out0;
wire v$G6_7901_out0;
wire v$G6_7902_out0;
wire v$G6_8632_out0;
wire v$G6_8633_out0;
wire v$G6_9184_out0;
wire v$G6_9185_out0;
wire v$G70_6845_out0;
wire v$G70_6846_out0;
wire v$G70_9421_out0;
wire v$G71_10591_out0;
wire v$G71_10592_out0;
wire v$G72_3918_out0;
wire v$G74_10988_out0;
wire v$G77_12941_out0;
wire v$G78_4825_out0;
wire v$G79_8390_out0;
wire v$G7_10034_out0;
wire v$G7_10035_out0;
wire v$G7_1007_out0;
wire v$G7_1008_out0;
wire v$G7_10153_out0;
wire v$G7_1164_out0;
wire v$G7_1165_out0;
wire v$G7_1166_out0;
wire v$G7_1167_out0;
wire v$G7_12491_out0;
wire v$G7_12865_out0;
wire v$G7_12866_out0;
wire v$G7_12867_out0;
wire v$G7_12868_out0;
wire v$G7_12869_out0;
wire v$G7_12870_out0;
wire v$G7_12871_out0;
wire v$G7_12872_out0;
wire v$G7_12873_out0;
wire v$G7_12874_out0;
wire v$G7_12875_out0;
wire v$G7_12876_out0;
wire v$G7_12877_out0;
wire v$G7_12878_out0;
wire v$G7_12879_out0;
wire v$G7_12880_out0;
wire v$G7_12881_out0;
wire v$G7_12882_out0;
wire v$G7_12883_out0;
wire v$G7_12884_out0;
wire v$G7_12885_out0;
wire v$G7_12886_out0;
wire v$G7_12887_out0;
wire v$G7_12888_out0;
wire v$G7_12889_out0;
wire v$G7_12890_out0;
wire v$G7_12891_out0;
wire v$G7_12892_out0;
wire v$G7_12893_out0;
wire v$G7_12894_out0;
wire v$G7_12895_out0;
wire v$G7_12896_out0;
wire v$G7_12897_out0;
wire v$G7_12898_out0;
wire v$G7_12899_out0;
wire v$G7_12900_out0;
wire v$G7_12901_out0;
wire v$G7_12902_out0;
wire v$G7_12903_out0;
wire v$G7_12904_out0;
wire v$G7_12905_out0;
wire v$G7_12906_out0;
wire v$G7_12907_out0;
wire v$G7_12908_out0;
wire v$G7_12909_out0;
wire v$G7_12910_out0;
wire v$G7_12911_out0;
wire v$G7_12912_out0;
wire v$G7_12913_out0;
wire v$G7_12914_out0;
wire v$G7_12915_out0;
wire v$G7_12916_out0;
wire v$G7_12917_out0;
wire v$G7_12918_out0;
wire v$G7_12919_out0;
wire v$G7_12920_out0;
wire v$G7_12921_out0;
wire v$G7_12922_out0;
wire v$G7_12923_out0;
wire v$G7_12924_out0;
wire v$G7_13277_out0;
wire v$G7_13278_out0;
wire v$G7_1889_out0;
wire v$G7_1890_out0;
wire v$G7_5269_out0;
wire v$G7_5270_out0;
wire v$G7_5374_out0;
wire v$G7_5375_out0;
wire v$G7_6593_out0;
wire v$G7_6594_out0;
wire v$G7_6595_out0;
wire v$G7_6596_out0;
wire v$G7_6597_out0;
wire v$G7_6598_out0;
wire v$G7_6599_out0;
wire v$G7_6600_out0;
wire v$G7_6601_out0;
wire v$G7_6602_out0;
wire v$G7_6603_out0;
wire v$G7_6604_out0;
wire v$G7_6605_out0;
wire v$G7_6606_out0;
wire v$G7_6607_out0;
wire v$G7_6608_out0;
wire v$G7_6617_out0;
wire v$G7_6658_out0;
wire v$G7_6659_out0;
wire v$G7_7231_out0;
wire v$G7_7232_out0;
wire v$G7_727_out0;
wire v$G7_728_out0;
wire v$G7_7596_out0;
wire v$G7_7597_out0;
wire v$G7_7976_out0;
wire v$G7_7977_out0;
wire v$G7_8288_out0;
wire v$G7_8289_out0;
wire v$G7_9002_out0;
wire v$G7_9003_out0;
wire v$G7_9129_out0;
wire v$G7_9130_out0;
wire v$G7_9511_out0;
wire v$G7_9512_out0;
wire v$G7_9513_out0;
wire v$G7_9514_out0;
wire v$G7_9515_out0;
wire v$G7_9516_out0;
wire v$G7_9517_out0;
wire v$G7_9518_out0;
wire v$G7_9519_out0;
wire v$G7_9520_out0;
wire v$G7_9521_out0;
wire v$G7_9522_out0;
wire v$G7_9703_out0;
wire v$G7_9704_out0;
wire v$G83_357_out0;
wire v$G84_504_out0;
wire v$G85_4217_out0;
wire v$G86_9099_out0;
wire v$G87_3518_out0;
wire v$G88_4994_out0;
wire v$G89_12562_out0;
wire v$G8_1036_out0;
wire v$G8_1037_out0;
wire v$G8_1038_out0;
wire v$G8_1039_out0;
wire v$G8_1040_out0;
wire v$G8_1041_out0;
wire v$G8_1042_out0;
wire v$G8_1043_out0;
wire v$G8_10770_out0;
wire v$G8_10771_out0;
wire v$G8_10979_out0;
wire v$G8_1170_out0;
wire v$G8_1171_out0;
wire v$G8_1189_out0;
wire v$G8_1190_out0;
wire v$G8_12674_out0;
wire v$G8_12675_out0;
wire v$G8_13406_out0;
wire v$G8_13407_out0;
wire v$G8_1349_out0;
wire v$G8_1350_out0;
wire v$G8_211_out0;
wire v$G8_212_out0;
wire v$G8_2439_out0;
wire v$G8_2440_out0;
wire v$G8_2441_out0;
wire v$G8_2442_out0;
wire v$G8_2443_out0;
wire v$G8_2444_out0;
wire v$G8_2445_out0;
wire v$G8_2446_out0;
wire v$G8_2447_out0;
wire v$G8_2448_out0;
wire v$G8_2449_out0;
wire v$G8_2450_out0;
wire v$G8_2451_out0;
wire v$G8_2452_out0;
wire v$G8_2453_out0;
wire v$G8_2454_out0;
wire v$G8_2455_out0;
wire v$G8_2456_out0;
wire v$G8_2457_out0;
wire v$G8_2458_out0;
wire v$G8_2459_out0;
wire v$G8_2460_out0;
wire v$G8_2461_out0;
wire v$G8_2462_out0;
wire v$G8_3224_out0;
wire v$G8_3225_out0;
wire v$G8_4049_out0;
wire v$G8_4050_out0;
wire v$G8_4071_out0;
wire v$G8_4072_out0;
wire v$G8_509_out0;
wire v$G8_510_out0;
wire v$G8_6322_out0;
wire v$G8_6323_out0;
wire v$G8_6485_out0;
wire v$G8_6486_out0;
wire v$G8_7301_out0;
wire v$G8_7302_out0;
wire v$G8_7762_out0;
wire v$G8_7763_out0;
wire v$G8_7764_out0;
wire v$G8_7765_out0;
wire v$G8_7766_out0;
wire v$G8_7767_out0;
wire v$G8_7768_out0;
wire v$G8_7769_out0;
wire v$G8_7770_out0;
wire v$G8_7771_out0;
wire v$G8_7772_out0;
wire v$G8_7773_out0;
wire v$G8_7774_out0;
wire v$G8_7775_out0;
wire v$G8_7776_out0;
wire v$G8_7777_out0;
wire v$G8_7778_out0;
wire v$G8_7779_out0;
wire v$G8_7780_out0;
wire v$G8_7781_out0;
wire v$G8_7782_out0;
wire v$G8_7783_out0;
wire v$G8_7784_out0;
wire v$G8_7785_out0;
wire v$G8_7786_out0;
wire v$G8_7787_out0;
wire v$G8_7788_out0;
wire v$G8_7789_out0;
wire v$G8_7790_out0;
wire v$G8_7791_out0;
wire v$G8_7792_out0;
wire v$G8_7793_out0;
wire v$G8_7794_out0;
wire v$G8_7795_out0;
wire v$G8_7796_out0;
wire v$G8_7797_out0;
wire v$G8_7798_out0;
wire v$G8_7799_out0;
wire v$G8_7800_out0;
wire v$G8_7801_out0;
wire v$G8_7802_out0;
wire v$G8_7803_out0;
wire v$G8_7804_out0;
wire v$G8_7805_out0;
wire v$G8_7806_out0;
wire v$G8_7807_out0;
wire v$G8_7808_out0;
wire v$G8_7809_out0;
wire v$G8_7810_out0;
wire v$G8_7811_out0;
wire v$G8_7812_out0;
wire v$G8_7813_out0;
wire v$G8_7814_out0;
wire v$G8_7815_out0;
wire v$G8_7816_out0;
wire v$G8_7817_out0;
wire v$G8_7818_out0;
wire v$G8_7819_out0;
wire v$G8_7820_out0;
wire v$G8_7821_out0;
wire v$G8_8068_out0;
wire v$G8_8069_out0;
wire v$G8_8123_out0;
wire v$G8_8124_out0;
wire v$G8_8973_out0;
wire v$G8_8974_out0;
wire v$G8_9652_out0;
wire v$G8_9653_out0;
wire v$G8_9654_out0;
wire v$G8_9655_out0;
wire v$G8_9656_out0;
wire v$G8_9657_out0;
wire v$G8_9658_out0;
wire v$G8_9659_out0;
wire v$G8_9660_out0;
wire v$G8_9661_out0;
wire v$G8_9662_out0;
wire v$G8_9663_out0;
wire v$G90_5561_out0;
wire v$G9_10434_out0;
wire v$G9_10435_out0;
wire v$G9_10503_out0;
wire v$G9_10504_out0;
wire v$G9_10505_out0;
wire v$G9_10506_out0;
wire v$G9_10507_out0;
wire v$G9_10508_out0;
wire v$G9_10509_out0;
wire v$G9_10510_out0;
wire v$G9_10511_out0;
wire v$G9_10512_out0;
wire v$G9_10513_out0;
wire v$G9_10514_out0;
wire v$G9_10515_out0;
wire v$G9_10516_out0;
wire v$G9_10517_out0;
wire v$G9_10518_out0;
wire v$G9_10813_out0;
wire v$G9_10814_out0;
wire v$G9_10859_out0;
wire v$G9_10860_out0;
wire v$G9_11217_out0;
wire v$G9_11218_out0;
wire v$G9_11572_out0;
wire v$G9_11573_out0;
wire v$G9_11973_out0;
wire v$G9_11974_out0;
wire v$G9_12027_out0;
wire v$G9_12028_out0;
wire v$G9_12066_out0;
wire v$G9_12067_out0;
wire v$G9_12395_out0;
wire v$G9_12396_out0;
wire v$G9_12397_out0;
wire v$G9_12398_out0;
wire v$G9_12399_out0;
wire v$G9_12400_out0;
wire v$G9_12401_out0;
wire v$G9_12402_out0;
wire v$G9_12403_out0;
wire v$G9_12404_out0;
wire v$G9_12405_out0;
wire v$G9_12406_out0;
wire v$G9_12407_out0;
wire v$G9_12408_out0;
wire v$G9_12409_out0;
wire v$G9_12410_out0;
wire v$G9_12411_out0;
wire v$G9_12412_out0;
wire v$G9_12413_out0;
wire v$G9_12414_out0;
wire v$G9_12415_out0;
wire v$G9_12416_out0;
wire v$G9_12417_out0;
wire v$G9_12418_out0;
wire v$G9_12419_out0;
wire v$G9_12420_out0;
wire v$G9_12421_out0;
wire v$G9_12422_out0;
wire v$G9_12423_out0;
wire v$G9_12424_out0;
wire v$G9_12425_out0;
wire v$G9_12426_out0;
wire v$G9_12427_out0;
wire v$G9_12428_out0;
wire v$G9_12429_out0;
wire v$G9_12430_out0;
wire v$G9_12431_out0;
wire v$G9_12432_out0;
wire v$G9_12433_out0;
wire v$G9_12434_out0;
wire v$G9_12435_out0;
wire v$G9_12436_out0;
wire v$G9_12437_out0;
wire v$G9_12438_out0;
wire v$G9_12439_out0;
wire v$G9_12440_out0;
wire v$G9_12441_out0;
wire v$G9_12442_out0;
wire v$G9_12443_out0;
wire v$G9_12444_out0;
wire v$G9_12445_out0;
wire v$G9_12446_out0;
wire v$G9_12447_out0;
wire v$G9_12448_out0;
wire v$G9_12449_out0;
wire v$G9_12450_out0;
wire v$G9_12451_out0;
wire v$G9_12452_out0;
wire v$G9_12453_out0;
wire v$G9_12454_out0;
wire v$G9_12526_out0;
wire v$G9_12527_out0;
wire v$G9_1435_out0;
wire v$G9_1436_out0;
wire v$G9_2141_out0;
wire v$G9_2142_out0;
wire v$G9_3818_out0;
wire v$G9_3819_out0;
wire v$G9_4233_out0;
wire v$G9_4234_out0;
wire v$G9_4349_out0;
wire v$G9_4350_out0;
wire v$G9_473_out0;
wire v$G9_474_out0;
wire v$G9_5922_out0;
wire v$G9_5923_out0;
wire v$G9_9012_out0;
wire v$G9_9013_out0;
wire v$HALT$PREV$PREV$PREV_5277_out0;
wire v$HALT$PREV$PREV$PREV_5278_out0;
wire v$HALT$PREV$PREV_12829_out0;
wire v$HALT$PREV$PREV_12830_out0;
wire v$HALT$PREV_6935_out0;
wire v$HALT$PREV_6936_out0;
wire v$HALT0_290_out0;
wire v$HALT0_3824_out0;
wire v$HALT0_7510_out0;
wire v$HALT0_9525_out0;
wire v$HALT1_13013_out0;
wire v$HALT1_1859_out0;
wire v$HALT1_2849_out0;
wire v$HALT1_4838_out0;
wire v$HALTED_7627_out0;
wire v$HALTED_7628_out0;
wire v$HALTSEL_10098_out0;
wire v$HALTVALID_5289_out0;
wire v$HALTVALID_8869_out0;
wire v$HALT_11481_out0;
wire v$HALT_12505_out0;
wire v$HALT_12506_out0;
wire v$HALT_1675_out0;
wire v$HALT_1676_out0;
wire v$HALT_5113_out0;
wire v$HALT_5114_out0;
wire v$HALT_531_out0;
wire v$HALT_8544_out0;
wire v$HALT_8545_out0;
wire v$HIGHER$OUT_2537_out0;
wire v$HIGHER$OUT_2538_out0;
wire v$HIGHER$OUT_2539_out0;
wire v$HIGHER$OUT_2540_out0;
wire v$HIGHER$OUT_2541_out0;
wire v$HIGHER$OUT_2542_out0;
wire v$HIGHER$OUT_2543_out0;
wire v$HIGHER$OUT_2544_out0;
wire v$HIGHER$OUT_5318_out0;
wire v$HIGHER$OUT_5319_out0;
wire v$HIGHER$OUT_5320_out0;
wire v$HIGHER$OUT_5321_out0;
wire v$HIGHER$SAME_10331_out0;
wire v$HIGHER$SAME_10332_out0;
wire v$HIGHER$SAME_10333_out0;
wire v$HIGHER$SAME_10334_out0;
wire v$HIGHER$SAME_10335_out0;
wire v$HIGHER$SAME_10336_out0;
wire v$HIGHER$SAME_10337_out0;
wire v$HIGHER$SAME_10338_out0;
wire v$HIGHER$SAME_6366_out0;
wire v$HIGHER$SAME_6367_out0;
wire v$HIGHER$SAME_6368_out0;
wire v$HIGHER$SAME_6369_out0;
wire v$I0EN_5551_out0;
wire v$I0EN_5552_out0;
wire v$I0P_1365_out0;
wire v$I0P_1366_out0;
wire v$I0P_3002_out0;
wire v$I0P_3003_out0;
wire v$I0P_6869_out0;
wire v$I0P_6870_out0;
wire v$I0REGISTERWRITE_2048_out0;
wire v$I0REGISTERWRITE_2049_out0;
wire v$I0_13167_out0;
wire v$I0_13168_out0;
wire v$I1EN_13089_out0;
wire v$I1EN_13090_out0;
wire v$I1P_10166_out0;
wire v$I1P_10167_out0;
wire v$I1P_1427_out0;
wire v$I1P_1428_out0;
wire v$I1P_4447_out0;
wire v$I1P_4448_out0;
wire v$I1REGISTERWRITE_1698_out0;
wire v$I1REGISTERWRITE_1699_out0;
wire v$I1_3282_out0;
wire v$I1_3283_out0;
wire v$I2EN_10989_out0;
wire v$I2EN_10990_out0;
wire v$I2P_1179_out0;
wire v$I2P_1180_out0;
wire v$I2P_4445_out0;
wire v$I2P_4446_out0;
wire v$I2P_5068_out0;
wire v$I2P_5069_out0;
wire v$I2REGISTERWRITE_7720_out0;
wire v$I2REGISTERWRITE_7721_out0;
wire v$I2_9881_out0;
wire v$I2_9882_out0;
wire v$I3EN_12565_out0;
wire v$I3EN_12566_out0;
wire v$I3P_6221_out0;
wire v$I3P_6222_out0;
wire v$I3P_7124_out0;
wire v$I3P_7125_out0;
wire v$I3P_9176_out0;
wire v$I3P_9177_out0;
wire v$I3REGISTERWRITE_521_out0;
wire v$I3REGISTERWRITE_522_out0;
wire v$I3_3228_out0;
wire v$I3_3229_out0;
wire v$IGNORE_11642_out0;
wire v$IGNORE_11643_out0;
wire v$IGNORE_3653_out0;
wire v$IGNORE_3654_out0;
wire v$IGNORE_5757_out0;
wire v$IGNORE_7524_out0;
wire v$IGNORE_7525_out0;
wire v$INCOMINGINTERRUPT_1054_out0;
wire v$INCOMINGINTERRUPT_1055_out0;
wire v$ININTERRUPT_433_out0;
wire v$ININTERRUPT_434_out0;
wire v$ININT_10758_out0;
wire v$ININT_10759_out0;
wire v$INITIAL$FETCH$OCCURRED_759_out0;
wire v$INITIAL$FETCH$OCCURRED_760_out0;
wire v$INIT_7077_out0;
wire v$INIT_7078_out0;
wire v$INT2_7675_out0;
wire v$INT2_7676_out0;
wire v$INT3_12861_out0;
wire v$INT3_12862_out0;
wire v$INT3_9426_out0;
wire v$INT3_9427_out0;
wire v$INTCAPTURE0_9104_out0;
wire v$INTCAPTURE0_9105_out0;
wire v$INTCLEAR_5308_out0;
wire v$INTCLEAR_5309_out0;
wire v$INTCLR_194_out0;
wire v$INTCLR_195_out0;
wire v$INTCOUNT_5050_out0;
wire v$INTCOUNT_5051_out0;
wire v$INTDISABLE_1581_out0;
wire v$INTDISABLE_1582_out0;
wire v$INTDISABLE_3392_out0;
wire v$INTDISABLE_3393_out0;
wire v$INTENABLE_12210_out0;
wire v$INTENABLE_12211_out0;
wire v$INTENABLE_1705_out0;
wire v$INTENABLE_1706_out0;
wire v$INTERRUPT0_7520_out0;
wire v$INTERRUPT0_7521_out0;
wire v$INTERRUPT0_979_out0;
wire v$INTERRUPT0_980_out0;
wire v$INTERRUPT1_12516_out0;
wire v$INTERRUPT1_12517_out0;
wire v$INTERRUPT1_5758_out0;
wire v$INTERRUPT1_5759_out0;
wire v$INTERRUPT2_2562_out0;
wire v$INTERRUPT2_2563_out0;
wire v$INTERRUPT2_857_out0;
wire v$INTERRUPT2_858_out0;
wire v$INTERRUPT3_1583_out0;
wire v$INTERRUPT3_1584_out0;
wire v$INTERRUPT3_2210_out0;
wire v$INTERRUPT3_2211_out0;
wire v$INTERRUPTOVERFLOW_10426_out0;
wire v$INTERRUPTOVERFLOW_10427_out0;
wire v$INTERRUPTOVERFLOW_1160_out0;
wire v$INTERRUPTOVERFLOW_1161_out0;
wire v$INTERRUPTSENABLED_6576_out0;
wire v$INTERRUPTSENABLED_6577_out0;
wire v$INTOVERFLOW_11219_out0;
wire v$INTOVERFLOW_11220_out0;
wire v$IR1$15_3786_out0;
wire v$IR1$15_3787_out0;
wire v$IR1$C$L_6754_out0;
wire v$IR1$C$L_6755_out0;
wire v$IR1$IS$FPU$ARITHMETIC_595_out0;
wire v$IR1$IS$FPU$ARITHMETIC_596_out0;
wire v$IR1$IS$LDST_8802_out0;
wire v$IR1$IS$LDST_8803_out0;
wire v$IR1$IS$STORE_3101_out0;
wire v$IR1$IS$STORE_3102_out0;
wire v$IR1$LS_11519_out0;
wire v$IR1$LS_11520_out0;
wire v$IR1$L_3512_out0;
wire v$IR1$L_3513_out0;
wire v$IR1$P_2407_out0;
wire v$IR1$P_2408_out0;
wire v$IR1$S$WB_264_out0;
wire v$IR1$S$WB_265_out0;
wire v$IR1$S_5370_out0;
wire v$IR1$S_5371_out0;
wire v$IR1$U_10127_out0;
wire v$IR1$U_10128_out0;
wire v$IR1$VALID$VIEWER_817_out0;
wire v$IR1$VALID$VIEWER_818_out0;
wire v$IR1$VALID_12593_out0;
wire v$IR1$VALID_12594_out0;
wire v$IR1$VALID_13109_out0;
wire v$IR1$VALID_13110_out0;
wire v$IR1$VALID_2556_out0;
wire v$IR1$VALID_2557_out0;
wire v$IR1$VALID_3778_out0;
wire v$IR1$VALID_3779_out0;
wire v$IR1$VALID_58_out0;
wire v$IR1$VALID_59_out0;
wire v$IR1$VALID_6451_out0;
wire v$IR1$VALID_6452_out0;
wire v$IR1$VALID_9411_out0;
wire v$IR1$VALID_9412_out0;
wire v$IR1$W_11628_out0;
wire v$IR1$W_11629_out0;
wire v$IR15_7010_out0;
wire v$IR15_7011_out0;
wire v$IR15_7240_out0;
wire v$IR15_7241_out0;
wire v$IR2$15_5012_out0;
wire v$IR2$15_5013_out0;
wire v$IR2$FPU$32BIT_7600_out0;
wire v$IR2$FPU$32BIT_7601_out0;
wire v$IR2$FPU$LOADA_10585_out0;
wire v$IR2$FPU$LOADA_10586_out0;
wire v$IR2$FPU$LOAD_2912_out0;
wire v$IR2$FPU$LOAD_2913_out0;
wire v$IR2$FPU$L_7070_out0;
wire v$IR2$FPU$L_7071_out0;
wire v$IR2$IS$FPU_1696_out0;
wire v$IR2$IS$FPU_1697_out0;
wire v$IR2$IS$FPU_4798_out0;
wire v$IR2$IS$FPU_4799_out0;
wire v$IR2$IS$FPU_7643_out0;
wire v$IR2$IS$FPU_7644_out0;
wire v$IR2$IS$LDST_3050_out0;
wire v$IR2$IS$LDST_3051_out0;
wire v$IR2$LS_11050_out0;
wire v$IR2$LS_11051_out0;
wire v$IR2$L_8105_out0;
wire v$IR2$L_8106_out0;
wire v$IR2$P_12145_out0;
wire v$IR2$P_12146_out0;
wire v$IR2$REG$IMMEDIATE_4213_out0;
wire v$IR2$REG$IMMEDIATE_4214_out0;
wire v$IR2$S$WB_12240_out0;
wire v$IR2$S$WB_12241_out0;
wire v$IR2$S_463_out0;
wire v$IR2$S_464_out0;
wire v$IR2$U_3921_out0;
wire v$IR2$U_3922_out0;
wire v$IR2$VALID$AND$NOT$FLOAD_3272_out0;
wire v$IR2$VALID$AND$NOT$FLOAD_3273_out0;
wire v$IR2$VALID$AND$NOT$FLOAD_4883_out0;
wire v$IR2$VALID$AND$NOT$FLOAD_4884_out0;
wire v$IR2$VALID$VIEWER_3820_out0;
wire v$IR2$VALID$VIEWER_3821_out0;
wire v$IR2$VALID_10171_out0;
wire v$IR2$VALID_10172_out0;
wire v$IR2$VALID_11092_out0;
wire v$IR2$VALID_11093_out0;
wire v$IR2$VALID_13383_out0;
wire v$IR2$VALID_13384_out0;
wire v$IR2$VALID_2898_out0;
wire v$IR2$VALID_2899_out0;
wire v$IR2$VALID_4452_out0;
wire v$IR2$VALID_4453_out0;
wire v$IR2$VALID_5003_out0;
wire v$IR2$VALID_5004_out0;
wire v$IR2$VALID_6998_out0;
wire v$IR2$VALID_6999_out0;
wire v$IR2$VALID_7594_out0;
wire v$IR2$VALID_7595_out0;
wire v$IR2$VALID_8838_out0;
wire v$IR2$VALID_8839_out0;
wire v$IR2$W_10422_out0;
wire v$IR2$W_10423_out0;
wire v$IS$32$BITS_12390_out0;
wire v$IS$32$BITS_12391_out0;
wire v$IS$32$BITS_2837_out0;
wire v$IS$32$BITS_2838_out0;
wire v$IS$32$BITS_527_out0;
wire v$IS$32$BITS_528_out0;
wire v$IS$32$BITS_9430_out0;
wire v$IS$32$BITS_9431_out0;
wire v$IS$32$BIT_7152_out0;
wire v$IS$32$BIT_7153_out0;
wire v$IS$32$BIT_7259_out0;
wire v$IS$32$BIT_7260_out0;
wire v$IS$A$LARGER_10027_out0;
wire v$IS$A$LARGER_10028_out0;
wire v$IS$A$LARGER_11176_out0;
wire v$IS$A$LARGER_11177_out0;
wire v$IS$A$LARGER_11880_out0;
wire v$IS$A$LARGER_11881_out0;
wire v$IS$A$LARGER_4806_out0;
wire v$IS$A$LARGER_4807_out0;
wire v$IS$A$LARGER_6990_out0;
wire v$IS$A$LARGER_6991_out0;
wire v$IS$FPU$HAZARD_278_out0;
wire v$IS$FPU$HAZARD_279_out0;
wire v$IS$IR1$FMUL_10613_out0;
wire v$IS$IR1$FMUL_10614_out0;
wire v$IS$IR1$FMUL_1725_out0;
wire v$IS$IR1$FMUL_1726_out0;
wire v$IS$IR2$DATA$PROCESSING_6664_out0;
wire v$IS$IR2$DATA$PROCESSING_6665_out0;
wire v$IS$SUB$MANTISA$ADDER_1897_out0;
wire v$IS$SUB$MANTISA$ADDER_1898_out0;
wire v$IS$SUB$VIEW_197_out0;
wire v$IS$SUB$VIEW_198_out0;
wire v$IS$SUB_10742_out0;
wire v$IS$SUB_10743_out0;
wire v$IS$SUB_3087_out0;
wire v$IS$SUB_3088_out0;
wire v$IS$SUB_8690_out0;
wire v$IS$SUB_8691_out0;
wire v$IS$SUM$0_10892_out0;
wire v$IS$SUM$0_10893_out0;
wire v$IS$SUM$0_10944_out0;
wire v$IS$SUM$0_10945_out0;
wire v$IS$SUM$0_402_out0;
wire v$IS$SUM$0_403_out0;
wire v$ISINTERRUPTED_7651_out0;
wire v$ISINTERRUPTED_7652_out0;
wire v$ISINTERRUPTED_7745_out0;
wire v$ISINTERRUPTED_7746_out0;
wire v$ISMOV_2786_out0;
wire v$ISMOV_2787_out0;
wire v$ISMOV_4660_out0;
wire v$ISMOV_4661_out0;
wire v$ISMOV_6007_out0;
wire v$ISMOV_6008_out0;
wire v$ISMOV_8272_out0;
wire v$ISMOV_8273_out0;
wire v$JEQ_12805_out0;
wire v$JEQ_12806_out0;
wire v$JEQ_869_out0;
wire v$JEQ_870_out0;
wire v$JLO_10309_out0;
wire v$JLO_10310_out0;
wire v$JLO_5611_out0;
wire v$JLO_5612_out0;
wire v$JLS_1096_out0;
wire v$JLS_1097_out0;
wire v$JLS_11527_out0;
wire v$JLS_11528_out0;
wire v$JMI_72_out0;
wire v$JMI_73_out0;
wire v$JMI_8762_out0;
wire v$JMI_8763_out0;
wire v$JMP_2998_out0;
wire v$JMP_2999_out0;
wire v$JMP_861_out0;
wire v$JMP_862_out0;
wire v$LASTQ_7873_out0;
wire v$LASTQ_7874_out0;
wire v$LASTQ_7875_out0;
wire v$LASTQ_7876_out0;
wire v$LASTQ_7877_out0;
wire v$LASTQ_7878_out0;
wire v$LASTQ_7879_out0;
wire v$LASTQ_7880_out0;
wire v$LASTQ_7881_out0;
wire v$LASTQ_7882_out0;
wire v$LASTQ_7883_out0;
wire v$LASTQ_7884_out0;
wire v$LASTQ_7885_out0;
wire v$LASTQ_7886_out0;
wire v$LASTQ_7887_out0;
wire v$LASTQ_7888_out0;
wire v$LASTQ_7889_out0;
wire v$LASTQ_7890_out0;
wire v$LASTQ_7891_out0;
wire v$LASTQ_7892_out0;
wire v$LASTQ_7893_out0;
wire v$LASTQ_7894_out0;
wire v$LDMAINPC_9191_out0;
wire v$LDMAINPC_9192_out0;
wire v$LDMAIN_1919_out0;
wire v$LDMAIN_1920_out0;
wire v$LDMAIN_9330_out0;
wire v$LDMAIN_9331_out0;
wire v$LDSTRAMMUX_11304_out0;
wire v$LDSTRAMMUX_11305_out0;
wire v$LEFT$SHIFT_6043_out0;
wire v$LEFT$SHIFT_6044_out0;
wire v$LEFT$SHIFT_6045_out0;
wire v$LEFT$SHIFT_6046_out0;
wire v$LEFT$SHIFT_6047_out0;
wire v$LEFT$SHIFT_6048_out0;
wire v$LEFT$SHIFT_6049_out0;
wire v$LEFT$SHIFT_6050_out0;
wire v$LEFT$SHIFT_8476_out0;
wire v$LEFT$SHIFT_8477_out0;
wire v$LEFT$SHIFT_8478_out0;
wire v$LEFT$SHIFT_8479_out0;
wire v$LEFT$SHIFT_8480_out0;
wire v$LEFT$SHIFT_8481_out0;
wire v$LEFT$SHIFT_8482_out0;
wire v$LEFT$SHIFT_8483_out0;
wire v$LEFT$SHIT_1795_out0;
wire v$LEFT$SHIT_1796_out0;
wire v$LEFT$SHIT_1797_out0;
wire v$LEFT$SHIT_1798_out0;
wire v$LEFT$SHIT_1799_out0;
wire v$LEFT$SHIT_1800_out0;
wire v$LEFT$SHIT_1801_out0;
wire v$LEFT$SHIT_1802_out0;
wire v$LEFT$SHIT_1803_out0;
wire v$LEFT$SHIT_1804_out0;
wire v$LEFT$SHIT_1805_out0;
wire v$LEFT$SHIT_1806_out0;
wire v$LEFT$SHIT_1807_out0;
wire v$LEFT$SHIT_1808_out0;
wire v$LEFT$SHIT_1809_out0;
wire v$LEFT$SHIT_1810_out0;
wire v$LEFT$SHIT_1811_out0;
wire v$LEFT$SHIT_1812_out0;
wire v$LEFT$SHIT_1813_out0;
wire v$LEFT$SHIT_1814_out0;
wire v$LEFT$SHIT_1815_out0;
wire v$LEFT$SHIT_1816_out0;
wire v$LEFT$SHIT_1817_out0;
wire v$LEFT$SHIT_1818_out0;
wire v$LEFT$SHIT_1819_out0;
wire v$LEFT$SHIT_1820_out0;
wire v$LEFT$SHIT_1821_out0;
wire v$LEFT$SHIT_1822_out0;
wire v$LEFT$SHIT_1823_out0;
wire v$LEFT$SHIT_1824_out0;
wire v$LEFT$SHIT_1825_out0;
wire v$LEFT$SHIT_1826_out0;
wire v$LEFT$SHIT_1827_out0;
wire v$LEFT$SHIT_1828_out0;
wire v$LEFT$SHIT_1829_out0;
wire v$LEFT$SHIT_1830_out0;
wire v$LEFT$SHIT_1831_out0;
wire v$LEFT$SHIT_1832_out0;
wire v$LEFT$SHIT_1833_out0;
wire v$LEFT$SHIT_1834_out0;
wire v$LEFT$SHIT_1835_out0;
wire v$LEFT$SHIT_1836_out0;
wire v$LEFT$SHIT_1837_out0;
wire v$LEFT$SHIT_1838_out0;
wire v$LEFT$SHIT_1839_out0;
wire v$LEFT$SHIT_1840_out0;
wire v$LEFT$SHIT_1841_out0;
wire v$LEFT$SHIT_1842_out0;
wire v$LEFT$SHIT_1843_out0;
wire v$LEFT$SHIT_1844_out0;
wire v$LEFT$SHIT_1845_out0;
wire v$LEFT$SHIT_1846_out0;
wire v$LEFT$SHIT_1847_out0;
wire v$LEFT$SHIT_1848_out0;
wire v$LEFT$SHIT_1849_out0;
wire v$LEFT$SHIT_1850_out0;
wire v$LEFT$SHIT_1851_out0;
wire v$LEFT$SHIT_1852_out0;
wire v$LEFT$SHIT_1853_out0;
wire v$LEFT$SHIT_1854_out0;
wire v$LEFT$SHIT_1855_out0;
wire v$LEFT$SHIT_1856_out0;
wire v$LEFT$SHIT_1857_out0;
wire v$LEFT$SHIT_1858_out0;
wire v$LOADA_3453_out0;
wire v$LOADA_3454_out0;
wire v$LOADA_3519_out0;
wire v$LOADA_3520_out0;
wire v$LOAD_4208_out0;
wire v$LOAD_4209_out0;
wire v$LOAD_7522_out0;
wire v$LOAD_7523_out0;
wire v$LOWER$OUT_2902_out0;
wire v$LOWER$OUT_2903_out0;
wire v$LOWER$OUT_2904_out0;
wire v$LOWER$OUT_2905_out0;
wire v$LOWER$OUT_2906_out0;
wire v$LOWER$OUT_2907_out0;
wire v$LOWER$OUT_2908_out0;
wire v$LOWER$OUT_2909_out0;
wire v$LOWER$OUT_4434_out0;
wire v$LOWER$OUT_4435_out0;
wire v$LOWER$OUT_4436_out0;
wire v$LOWER$OUT_4437_out0;
wire v$LOWER$PART_4327_out0;
wire v$LOWER$PART_4328_out0;
wire v$LOWER$PART_4329_out0;
wire v$LOWER$PART_4330_out0;
wire v$LOWER$SAME_2501_out0;
wire v$LOWER$SAME_2502_out0;
wire v$LOWER$SAME_2503_out0;
wire v$LOWER$SAME_2504_out0;
wire v$LOWER$SAME_6757_out0;
wire v$LOWER$SAME_6758_out0;
wire v$LOWER$SAME_6759_out0;
wire v$LOWER$SAME_6760_out0;
wire v$LOWER$SAME_6761_out0;
wire v$LOWER$SAME_6762_out0;
wire v$LOWER$SAME_6763_out0;
wire v$LOWER$SAME_6764_out0;
wire v$LSB_5342_out0;
wire v$LSB_5343_out0;
wire v$MANTISA$SAME_1363_out0;
wire v$MANTISA$SAME_1364_out0;
wire v$MEMHALT_12595_out0;
wire v$MEMHALT_12596_out0;
wire v$MI$LDST_12071_out0;
wire v$MI$LDST_12072_out0;
wire v$MI_1351_out0;
wire v$MI_1352_out0;
wire v$MI_4239_out0;
wire v$MI_4240_out0;
wire v$MI_5906_out0;
wire v$MI_5907_out0;
wire v$MI_7673_out0;
wire v$MI_7674_out0;
wire v$MI_7903_out0;
wire v$MI_7904_out0;
wire v$MI_8107_out0;
wire v$MI_8108_out0;
wire v$MI_9752_out0;
wire v$MI_9753_out0;
wire v$MODEEN_10428_out0;
wire v$MODEEN_10429_out0;
wire v$MODEEN_3782_out0;
wire v$MODEEN_3783_out0;
wire v$MODEWRITE_10070_out0;
wire v$MODEWRITE_10071_out0;
wire v$MULTIPLYING$BIT_1607_out0;
wire v$MULTIPLYING$BIT_1608_out0;
wire v$MULTIPLYING$BIT_1609_out0;
wire v$MULTIPLYING$BIT_1610_out0;
wire v$MULTIPLYING$BIT_1611_out0;
wire v$MULTIPLYING$BIT_1612_out0;
wire v$MULTIPLYING$BIT_1613_out0;
wire v$MULTIPLYING$BIT_1614_out0;
wire v$MULTIPLYING$BIT_1615_out0;
wire v$MULTIPLYING$BIT_1616_out0;
wire v$MULTIPLYING$BIT_1617_out0;
wire v$MULTIPLYING$BIT_1618_out0;
wire v$MULTIPLYING$BIT_1619_out0;
wire v$MULTIPLYING$BIT_1620_out0;
wire v$MULTIPLYING$BIT_1621_out0;
wire v$MULTIPLYING$BIT_1622_out0;
wire v$MULTIPLYING$BIT_1623_out0;
wire v$MULTIPLYING$BIT_1624_out0;
wire v$MULTIPLYING$BIT_1625_out0;
wire v$MULTIPLYING$BIT_1626_out0;
wire v$MULTIPLYING$BIT_1627_out0;
wire v$MULTIPLYING$BIT_1628_out0;
wire v$MULTIPLYING$BIT_1629_out0;
wire v$MULTIPLYING$BIT_1630_out0;
wire v$MUL_12088_out0;
wire v$MUL_12089_out0;
wire v$MUX10_10936_out0;
wire v$MUX10_10937_out0;
wire v$MUX10_10938_out0;
wire v$MUX10_10939_out0;
wire v$MUX10_11502_out0;
wire v$MUX10_11503_out0;
wire v$MUX11_12709_out0;
wire v$MUX11_12710_out0;
wire v$MUX11_12711_out0;
wire v$MUX11_12712_out0;
wire v$MUX11_487_out0;
wire v$MUX11_488_out0;
wire v$MUX12_12609_out0;
wire v$MUX12_12610_out0;
wire v$MUX12_12611_out0;
wire v$MUX12_12612_out0;
wire v$MUX13_9228_out0;
wire v$MUX13_9229_out0;
wire v$MUX13_9230_out0;
wire v$MUX13_9231_out0;
wire v$MUX14_1723_out0;
wire v$MUX14_1724_out0;
wire v$MUX14_3312_out0;
wire v$MUX14_3313_out0;
wire v$MUX14_3314_out0;
wire v$MUX14_3315_out0;
wire v$MUX15_547_out0;
wire v$MUX15_548_out0;
wire v$MUX15_549_out0;
wire v$MUX15_550_out0;
wire v$MUX16_11809_out0;
wire v$MUX16_11810_out0;
wire v$MUX16_11811_out0;
wire v$MUX16_11812_out0;
wire v$MUX17_11616_out0;
wire v$MUX17_11617_out0;
wire v$MUX17_11618_out0;
wire v$MUX17_11619_out0;
wire v$MUX18_3258_out0;
wire v$MUX18_3259_out0;
wire v$MUX18_3260_out0;
wire v$MUX18_3261_out0;
wire v$MUX19_4393_out0;
wire v$MUX19_4394_out0;
wire v$MUX19_4395_out0;
wire v$MUX19_4396_out0;
wire v$MUX1_12005_out0;
wire v$MUX1_12006_out0;
wire v$MUX1_12007_out0;
wire v$MUX1_12008_out0;
wire v$MUX1_12009_out0;
wire v$MUX1_12010_out0;
wire v$MUX1_12011_out0;
wire v$MUX1_12012_out0;
wire v$MUX1_12013_out0;
wire v$MUX1_12014_out0;
wire v$MUX1_12015_out0;
wire v$MUX1_12016_out0;
wire v$MUX1_12017_out0;
wire v$MUX1_12018_out0;
wire v$MUX1_12019_out0;
wire v$MUX1_12020_out0;
wire v$MUX1_12021_out0;
wire v$MUX1_12022_out0;
wire v$MUX1_12023_out0;
wire v$MUX1_12024_out0;
wire v$MUX1_12025_out0;
wire v$MUX1_12026_out0;
wire v$MUX1_1489_out0;
wire v$MUX1_1490_out0;
wire v$MUX1_1491_out0;
wire v$MUX1_1492_out0;
wire v$MUX1_1493_out0;
wire v$MUX1_1494_out0;
wire v$MUX1_1495_out0;
wire v$MUX1_1496_out0;
wire v$MUX1_1497_out0;
wire v$MUX1_1498_out0;
wire v$MUX1_1499_out0;
wire v$MUX1_1500_out0;
wire v$MUX1_1635_out0;
wire v$MUX1_1636_out0;
wire v$MUX1_1637_out0;
wire v$MUX1_1638_out0;
wire v$MUX1_3405_out0;
wire v$MUX1_3406_out0;
wire v$MUX1_345_out0;
wire v$MUX1_346_out0;
wire v$MUX1_5175_out0;
wire v$MUX1_5176_out0;
wire v$MUX20_7410_out0;
wire v$MUX20_7411_out0;
wire v$MUX20_7412_out0;
wire v$MUX20_7413_out0;
wire v$MUX21_3294_out0;
wire v$MUX21_3295_out0;
wire v$MUX21_3296_out0;
wire v$MUX21_3297_out0;
wire v$MUX22_11542_out0;
wire v$MUX22_11543_out0;
wire v$MUX22_11544_out0;
wire v$MUX22_11545_out0;
wire v$MUX23_11379_out0;
wire v$MUX23_11380_out0;
wire v$MUX23_11381_out0;
wire v$MUX23_11382_out0;
wire v$MUX24_12821_out0;
wire v$MUX24_12822_out0;
wire v$MUX24_12823_out0;
wire v$MUX24_12824_out0;
wire v$MUX25_5870_out0;
wire v$MUX25_5871_out0;
wire v$MUX25_5872_out0;
wire v$MUX25_5873_out0;
wire v$MUX2_3252_out0;
wire v$MUX2_3253_out0;
wire v$MUX2_4675_out0;
wire v$MUX2_4676_out0;
wire v$MUX2_8006_out0;
wire v$MUX2_8007_out0;
wire v$MUX2_8870_out0;
wire v$MUX2_8871_out0;
wire v$MUX2_9170_out0;
wire v$MUX2_9171_out0;
wire v$MUX2_9172_out0;
wire v$MUX2_9173_out0;
wire v$MUX2_9342_out0;
wire v$MUX2_9343_out0;
wire v$MUX2_9344_out0;
wire v$MUX2_9345_out0;
wire v$MUX2_9346_out0;
wire v$MUX2_9347_out0;
wire v$MUX2_9348_out0;
wire v$MUX2_9349_out0;
wire v$MUX2_9350_out0;
wire v$MUX2_9351_out0;
wire v$MUX2_9352_out0;
wire v$MUX2_9353_out0;
wire v$MUX3_12536_out0;
wire v$MUX3_12537_out0;
wire v$MUX3_4145_out0;
wire v$MUX3_4146_out0;
wire v$MUX3_5138_out0;
wire v$MUX3_5139_out0;
wire v$MUX3_5140_out0;
wire v$MUX3_5141_out0;
wire v$MUX3_665_out0;
wire v$MUX3_666_out0;
wire v$MUX3_6670_out0;
wire v$MUX3_6671_out0;
wire v$MUX3_6672_out0;
wire v$MUX3_6673_out0;
wire v$MUX3_6674_out0;
wire v$MUX3_6675_out0;
wire v$MUX3_6676_out0;
wire v$MUX3_6677_out0;
wire v$MUX3_6678_out0;
wire v$MUX3_6679_out0;
wire v$MUX3_6680_out0;
wire v$MUX3_6681_out0;
wire v$MUX4_10904_out0;
wire v$MUX4_10905_out0;
wire v$MUX4_11896_out0;
wire v$MUX4_11897_out0;
wire v$MUX4_11898_out0;
wire v$MUX4_11899_out0;
wire v$MUX4_11900_out0;
wire v$MUX4_11901_out0;
wire v$MUX4_11902_out0;
wire v$MUX4_11903_out0;
wire v$MUX4_11904_out0;
wire v$MUX4_11905_out0;
wire v$MUX4_11906_out0;
wire v$MUX4_11907_out0;
wire v$MUX4_12118_out0;
wire v$MUX4_12119_out0;
wire v$MUX4_5324_out0;
wire v$MUX4_5325_out0;
wire v$MUX4_5326_out0;
wire v$MUX4_5327_out0;
wire v$MUX4_7488_out0;
wire v$MUX4_7489_out0;
wire v$MUX4_8278_out0;
wire v$MUX4_8279_out0;
wire v$MUX5_10781_out0;
wire v$MUX5_10782_out0;
wire v$MUX5_12110_out0;
wire v$MUX5_12111_out0;
wire v$MUX5_13207_out0;
wire v$MUX5_13208_out0;
wire v$MUX5_4698_out0;
wire v$MUX5_4699_out0;
wire v$MUX5_4700_out0;
wire v$MUX5_4701_out0;
wire v$MUX5_6500_out0;
wire v$MUX5_6501_out0;
wire v$MUX5_6502_out0;
wire v$MUX5_6503_out0;
wire v$MUX5_6504_out0;
wire v$MUX5_6505_out0;
wire v$MUX5_6506_out0;
wire v$MUX5_6507_out0;
wire v$MUX5_6508_out0;
wire v$MUX5_6509_out0;
wire v$MUX5_6510_out0;
wire v$MUX5_6511_out0;
wire v$MUX5_7647_out0;
wire v$MUX5_7648_out0;
wire v$MUX6_11420_out0;
wire v$MUX6_11421_out0;
wire v$MUX6_11422_out0;
wire v$MUX6_11423_out0;
wire v$MUX6_6364_out0;
wire v$MUX6_6365_out0;
wire v$MUX6_6937_out0;
wire v$MUX6_6938_out0;
wire v$MUX6_6939_out0;
wire v$MUX6_6940_out0;
wire v$MUX6_6941_out0;
wire v$MUX6_6942_out0;
wire v$MUX6_6943_out0;
wire v$MUX6_6944_out0;
wire v$MUX6_6945_out0;
wire v$MUX6_6946_out0;
wire v$MUX6_6947_out0;
wire v$MUX6_6948_out0;
wire v$MUX6_9127_out0;
wire v$MUX6_9128_out0;
wire v$MUX6_9277_out0;
wire v$MUX6_9278_out0;
wire v$MUX7_12679_out0;
wire v$MUX7_12680_out0;
wire v$MUX7_12681_out0;
wire v$MUX7_12682_out0;
wire v$MUX7_12683_out0;
wire v$MUX7_12684_out0;
wire v$MUX7_12685_out0;
wire v$MUX7_12686_out0;
wire v$MUX7_12687_out0;
wire v$MUX7_12688_out0;
wire v$MUX7_12689_out0;
wire v$MUX7_12690_out0;
wire v$MUX7_496_out0;
wire v$MUX7_497_out0;
wire v$MUX7_498_out0;
wire v$MUX7_499_out0;
wire v$MUX7_6471_out0;
wire v$MUX7_6472_out0;
wire v$MUX7_7229_out0;
wire v$MUX7_7230_out0;
wire v$MUX8$OUT_8994_out0;
wire v$MUX8$OUT_8995_out0;
wire v$MUX8_1711_out0;
wire v$MUX8_1712_out0;
wire v$MUX8_1713_out0;
wire v$MUX8_1714_out0;
wire v$MUX8_2316_out0;
wire v$MUX8_2317_out0;
wire v$MUX8_2318_out0;
wire v$MUX8_2319_out0;
wire v$MUX8_2320_out0;
wire v$MUX8_2321_out0;
wire v$MUX8_2322_out0;
wire v$MUX8_2323_out0;
wire v$MUX8_2324_out0;
wire v$MUX8_2325_out0;
wire v$MUX8_2326_out0;
wire v$MUX8_2327_out0;
wire v$MUX8_3004_out0;
wire v$MUX8_3005_out0;
wire v$MUX8_725_out0;
wire v$MUX8_726_out0;
wire v$MUX9_5726_out0;
wire v$MUX9_5727_out0;
wire v$MUX9_5728_out0;
wire v$MUX9_5729_out0;
wire v$ModeRegAdd_2724_out0;
wire v$ModeRegAdd_2725_out0;
wire v$ModeWrite_3091_out0;
wire v$ModeWrite_3092_out0;
wire v$NEED$SHIFT$OP1_3226_out0;
wire v$NEED$SHIFT$OP1_3227_out0;
wire v$NEWINTERRUPT_3080_out0;
wire v$NEWINTERRUPT_3081_out0;
wire v$NEWINTERRUPT_3679_out0;
wire v$NEWINTERRUPT_3680_out0;
wire v$NEWINTERRUPT_4784_out0;
wire v$NEWINTERRUPT_4785_out0;
wire v$NEWINT_12597_out0;
wire v$NEWINT_12598_out0;
wire v$NEXTINTERRUPT_11825_out0;
wire v$NEXTINTERRUPT_11826_out0;
wire v$NEXTINTERRUPT_13115_out0;
wire v$NEXTINTERRUPT_13116_out0;
wire v$NEXTINTERRUPT_13199_out0;
wire v$NEXTINTERRUPT_13200_out0;
wire v$NEXTINTERRUPT_8406_out0;
wire v$NEXTINTERRUPT_8407_out0;
wire v$NEXTINT_4763_out0;
wire v$NEXTINT_4764_out0;
wire v$NEXTSTATE_9107_out0;
wire v$NEXTSTATE_9108_out0;
wire v$NEXTSTATE_9109_out0;
wire v$NE_2135_out0;
wire v$NE_2136_out0;
wire v$NF_9947_out0;
wire v$NF_9948_out0;
wire v$NOT$USED$CARRY_13402_out0;
wire v$NOT$USED$CARRY_13403_out0;
wire v$NOT$USED$CARRY_13404_out0;
wire v$NOT$USED$CARRY_13405_out0;
wire v$NOT$USED1_9760_out0;
wire v$NOT$USED1_9761_out0;
wire v$NOT$USED1_9762_out0;
wire v$NOT$USED1_9763_out0;
wire v$NOT$USED1_9764_out0;
wire v$NOT$USED1_9765_out0;
wire v$NOT$USED1_9766_out0;
wire v$NOT$USED1_9767_out0;
wire v$NOT$USED_11148_out0;
wire v$NOT$USED_11149_out0;
wire v$NOT$USED_11150_out0;
wire v$NOT$USED_11151_out0;
wire v$NOT$USED_1667_out0;
wire v$NOT$USED_1668_out0;
wire v$NOT$USED_3696_out0;
wire v$NOT$USED_3697_out0;
wire v$NP_4857_out0;
wire v$NP_4858_out0;
wire v$NQ0_10672_out0;
wire v$NQ0_10673_out0;
wire v$NQ0_10890_out0;
wire v$NQ0_10891_out0;
wire v$NQ0_5322_out0;
wire v$NQ0_5323_out0;
wire v$NQ1_11780_out0;
wire v$NQ1_11781_out0;
wire v$NQ1_219_out0;
wire v$NQ1_220_out0;
wire v$NQ1_7276_out0;
wire v$NQ1_7277_out0;
wire v$NQ2_11764_out0;
wire v$NQ2_11765_out0;
wire v$NQ2_13211_out0;
wire v$NQ2_13212_out0;
wire v$NQ2_1741_out0;
wire v$NQ2_1742_out0;
wire v$NQ3_1759_out0;
wire v$NQ3_1760_out0;
wire v$NQ3_721_out0;
wire v$NQ3_722_out0;
wire v$NR_11728_out0;
wire v$NR_11729_out0;
wire v$NS_12937_out0;
wire v$NS_12938_out0;
wire v$ODDPARITY_11132_out0;
wire v$ODDPARITY_11133_out0;
wire v$OFF_2756_out0;
wire v$OFF_2757_out0;
wire v$OUTPUT_13145_out0;
wire v$OUTPUT_6891_out0;
wire v$OUTPUT_6892_out0;
wire v$OUT_2549_out0;
wire v$OUT_2550_out0;
wire v$OUT_2622_out0;
wire v$OUT_2623_out0;
wire v$OUT_2624_out0;
wire v$OUT_2625_out0;
wire v$OUT_2626_out0;
wire v$OUT_2627_out0;
wire v$OUT_2628_out0;
wire v$OUT_2629_out0;
wire v$OUT_2630_out0;
wire v$OUT_2631_out0;
wire v$OUT_2632_out0;
wire v$OUT_2633_out0;
wire v$OUT_2634_out0;
wire v$OUT_2635_out0;
wire v$OUT_2636_out0;
wire v$OUT_2637_out0;
wire v$OUT_2638_out0;
wire v$OUT_2639_out0;
wire v$OUT_2640_out0;
wire v$OUT_2641_out0;
wire v$OUT_2642_out0;
wire v$OUT_2643_out0;
wire v$OUT_2644_out0;
wire v$OUT_2645_out0;
wire v$OUT_2646_out0;
wire v$OUT_2647_out0;
wire v$OUT_2648_out0;
wire v$OUT_2649_out0;
wire v$OUT_2650_out0;
wire v$OUT_2651_out0;
wire v$OUT_2652_out0;
wire v$OUT_2653_out0;
wire v$OUT_6185_out0;
wire v$OUT_6186_out0;
wire v$OUT_6187_out0;
wire v$OUT_6188_out0;
wire v$OUT_6467_out0;
wire v$OUT_6468_out0;
wire v$OUT_6469_out0;
wire v$OUT_6470_out0;
wire v$OUT_9286_out0;
wire v$OUT_9287_out0;
wire v$OUT_9288_out0;
wire v$OUT_9289_out0;
wire v$OUT_9290_out0;
wire v$OUT_9291_out0;
wire v$OUT_9292_out0;
wire v$OUT_9293_out0;
wire v$OVERFLOW_10307_out0;
wire v$OVERFLOW_10308_out0;
wire v$OVERFLOW_13127_out0;
wire v$OVERFLOW_13128_out0;
wire v$OVERFLOW_13177_out0;
wire v$OVERFLOW_13178_out0;
wire v$OVERFLOW_2338_out0;
wire v$OVERFLOW_2339_out0;
wire v$OVERFLOW_355_out0;
wire v$OVERFLOW_356_out0;
wire v$OddParity_7008_out0;
wire v$OddParity_7009_out0;
wire v$PARITY_7858_out0;
wire v$PARITY_7859_out0;
wire v$PCHALTVIEWER_947_out0;
wire v$PCHALT_11644_out0;
wire v$PCHALT_8399_out0;
wire v$PHALT0$PREV_5150_out0;
wire v$PHALT0_7479_out0;
wire v$PHALT1$PREV_4956_out0;
wire v$PHALT1_6182_out0;
wire v$PHALTVIEWER_1551_out0;
wire v$PHALT_10440_out0;
wire v$PHALT_12284_out0;
wire v$PHALT_834_out0;
wire v$PIPELINE$RESTART_13261_out0;
wire v$PIPELINE$RESTART_13262_out0;
wire v$PIPELINE$RESTART_4073_out0;
wire v$PIPELINE$RESTART_4074_out0;
wire v$PIPELINEHALT_10164_out0;
wire v$PIPELINEHALT_10165_out0;
wire v$PIPELINERESTART_1353_out0;
wire v$PIPELINERESTART_1354_out0;
wire v$P_5784_out0;
wire v$P_5785_out0;
wire v$ParityCheck_11289_out0;
wire v$ParityCheck_11290_out0;
wire v$ParityEN_11013_out0;
wire v$ParityEN_11014_out0;
wire v$Q0P_11821_out0;
wire v$Q0P_11822_out0;
wire v$Q0P_7944_out0;
wire v$Q0P_7945_out0;
wire v$Q0_13018_out0;
wire v$Q0_13019_out0;
wire v$Q0_74_out0;
wire v$Q0_75_out0;
wire v$Q0_9249_out0;
wire v$Q0_9250_out0;
wire v$Q1P_3774_out0;
wire v$Q1P_3775_out0;
wire v$Q1P_7261_out0;
wire v$Q1P_7262_out0;
wire v$Q1_3089_out0;
wire v$Q1_3090_out0;
wire v$Q1_7197_out0;
wire v$Q1_7198_out0;
wire v$Q1_9713_out0;
wire v$Q1_9714_out0;
wire v$Q2P_2850_out0;
wire v$Q2P_2851_out0;
wire v$Q2P_4041_out0;
wire v$Q2P_4042_out0;
wire v$Q2_12285_out0;
wire v$Q2_12286_out0;
wire v$Q2_1883_out0;
wire v$Q2_1884_out0;
wire v$Q2_3703_out0;
wire v$Q2_3704_out0;
wire v$Q3P_7500_out0;
wire v$Q3P_7501_out0;
wire v$Q3P_9332_out0;
wire v$Q3P_9333_out0;
wire v$Q3_12999_out0;
wire v$Q3_13000_out0;
wire v$Q3_13107_out0;
wire v$Q3_13108_out0;
wire v$Q_9528_out0;
wire v$Q_9529_out0;
wire v$Q_9530_out0;
wire v$Q_9531_out0;
wire v$Q_9532_out0;
wire v$Q_9533_out0;
wire v$Q_9534_out0;
wire v$Q_9535_out0;
wire v$Q_9536_out0;
wire v$Q_9537_out0;
wire v$Q_9538_out0;
wire v$Q_9539_out0;
wire v$Q_9540_out0;
wire v$Q_9541_out0;
wire v$Q_9542_out0;
wire v$Q_9543_out0;
wire v$Q_9544_out0;
wire v$Q_9545_out0;
wire v$Q_9546_out0;
wire v$Q_9547_out0;
wire v$Q_9548_out0;
wire v$Q_9549_out0;
wire v$R0_10497_out0;
wire v$R0_10498_out0;
wire v$R0_1143_out0;
wire v$R0_4666_out0;
wire v$R1_10327_out0;
wire v$R1_10328_out0;
wire v$R1_12676_out0;
wire v$R1_7681_out0;
wire v$R2_2554_out0;
wire v$R2_2555_out0;
wire v$R3_10621_out0;
wire v$R3_10622_out0;
wire v$RAMWEN0_11645_out0;
wire v$RAMWEN1_7089_out0;
wire v$RAMWENVIEWER_12120_out0;
wire v$RAMWEN_10932_out0;
wire v$RAMWEN_10933_out0;
wire v$RAMWEN_12732_out0;
wire v$RAMWEN_5302_out0;
wire v$RAMWEN_5303_out0;
wire v$READ$REQUEST0_13146_out0;
wire v$READ$REQUEST0_7434_out0;
wire v$READ$REQUEST1_11877_out0;
wire v$READ$REQUEST1_4462_out0;
wire v$READ$REQUEST_11632_out0;
wire v$READ$REQUEST_11633_out0;
wire v$READ$REQUEST_5332_out0;
wire v$READ$REQUEST_5333_out0;
wire v$READ$REQUEST_9841_out0;
wire v$READ$REQUEST_9842_out0;
wire v$RECIEVEDPARITY_4231_out0;
wire v$RECIEVEDPARITY_4232_out0;
wire v$RR0VIEWER_10024_out0;
wire v$RR0_5596_out0;
wire v$RR1REGoutVIEWER_4979_out0;
wire v$RR1VIEWER_10343_out0;
wire v$RR1_1093_out0;
wire v$RXBIT_6165_out0;
wire v$RXBIT_6166_out0;
wire v$RXCLK_11062_out0;
wire v$RXCLK_11063_out0;
wire v$RXCLK_507_out0;
wire v$RXCLK_508_out0;
wire v$RXDISABLE_5404_out0;
wire v$RXDISABLE_5405_out0;
wire v$RXENABLE_2429_out0;
wire v$RXENABLE_2430_out0;
wire v$RXErrorSet_2187_out0;
wire v$RXErrorSet_2188_out0;
wire v$RXFLAG_10319_out0;
wire v$RXFLAG_10320_out0;
wire v$RXFLAG_7909_out0;
wire v$RXFLAG_7910_out0;
wire v$RXFlagSet_6347_out0;
wire v$RXFlagSet_6348_out0;
wire v$RXINTERRUPT_10185_out0;
wire v$RXINTERRUPT_10186_out0;
wire v$RXINTERRUPT_10643_out0;
wire v$RXINTERRUPT_10644_out0;
wire v$RXINT_8180_out0;
wire v$RXINT_8181_out0;
wire v$RXREAD_10641_out0;
wire v$RXREAD_10642_out0;
wire v$RXREAD_11072_out0;
wire v$RXREAD_11073_out0;
wire v$RXRead_11475_out0;
wire v$RXRead_11476_out0;
wire v$RXRegAdd_8613_out0;
wire v$RXRegAdd_8614_out0;
wire v$RXReset_11610_out0;
wire v$RXReset_11611_out0;
wire v$RXSET_10048_out0;
wire v$RXSET_10049_out0;
wire v$RXSHIFT_388_out0;
wire v$RXSHIFT_389_out0;
wire v$RX_1727_out0;
wire v$RX_1728_out0;
wire v$RX_3217_out0;
wire v$RX_3218_out0;
wire v$RX_40_out0;
wire v$RX_41_out0;
wire v$RX_4204_out0;
wire v$RX_4205_out0;
wire v$RX_4652_out0;
wire v$RX_4653_out0;
wire v$RXflag_11059_out0;
wire v$RXflag_11060_out0;
wire v$RXlast_8470_out0;
wire v$RXlast_8471_out0;
wire v$RXoverflow_6516_out0;
wire v$RXoverflow_6517_out0;
wire v$RXreset_3961_out0;
wire v$RXreset_3962_out0;
wire v$RXset_3477_out0;
wire v$RXset_3478_out0;
wire v$RXset_891_out0;
wire v$RXset_892_out0;
wire v$R_11791_out0;
wire v$R_13032_out0;
wire v$R_13033_out0;
wire v$R_13034_out0;
wire v$R_13035_out0;
wire v$R_13036_out0;
wire v$R_13037_out0;
wire v$R_13038_out0;
wire v$R_13039_out0;
wire v$R_13040_out0;
wire v$R_13041_out0;
wire v$R_13042_out0;
wire v$R_13043_out0;
wire v$R_13044_out0;
wire v$R_13045_out0;
wire v$R_13046_out0;
wire v$R_13047_out0;
wire v$R_13048_out0;
wire v$R_13049_out0;
wire v$R_13050_out0;
wire v$R_13051_out0;
wire v$R_13052_out0;
wire v$R_13053_out0;
wire v$R_6019_out0;
wire v$R_6020_out0;
wire v$R_719_out0;
wire v$R_720_out0;
wire v$R_789_out0;
wire v$R_790_out0;
wire v$R_791_out0;
wire v$RceivedParity_13191_out0;
wire v$RceivedParity_13192_out0;
wire v$RecievedParity_6514_out0;
wire v$RecievedParity_6515_out0;
wire v$SAME$H_451_out0;
wire v$SAME$H_452_out0;
wire v$SAME$H_6167_out0;
wire v$SAME$H_6168_out0;
wire v$SAME$L_11525_out0;
wire v$SAME$L_11526_out0;
wire v$SAME$L_6459_out0;
wire v$SAME$L_6460_out0;
wire v$SAME_13064_out0;
wire v$SAME_13065_out0;
wire v$SAME_13066_out0;
wire v$SAME_13067_out0;
wire v$SAME_13068_out0;
wire v$SAME_13069_out0;
wire v$SAME_13070_out0;
wire v$SAME_13071_out0;
wire v$SAME_13351_out0;
wire v$SAME_13352_out0;
wire v$SAME_13353_out0;
wire v$SAME_13354_out0;
wire v$SAME_13355_out0;
wire v$SAME_13356_out0;
wire v$SAME_13357_out0;
wire v$SAME_13358_out0;
wire v$SAME_13359_out0;
wire v$SAME_13360_out0;
wire v$SAME_13361_out0;
wire v$SAME_13362_out0;
wire v$SAME_13363_out0;
wire v$SAME_13364_out0;
wire v$SAME_13365_out0;
wire v$SAME_13366_out0;
wire v$SAME_13367_out0;
wire v$SAME_13368_out0;
wire v$SAME_13369_out0;
wire v$SAME_13370_out0;
wire v$SAME_13371_out0;
wire v$SAME_13372_out0;
wire v$SAME_13373_out0;
wire v$SAME_13374_out0;
wire v$SAME_13375_out0;
wire v$SAME_13376_out0;
wire v$SAME_13377_out0;
wire v$SAME_13378_out0;
wire v$SAME_13379_out0;
wire v$SAME_13380_out0;
wire v$SAME_13381_out0;
wire v$SAME_13382_out0;
wire v$SAME_4265_out0;
wire v$SAME_4266_out0;
wire v$SAME_6171_out0;
wire v$SAME_6172_out0;
wire v$SAME_6173_out0;
wire v$SAME_6174_out0;
wire v$SEL10_2841_out0;
wire v$SEL10_2842_out0;
wire v$SEL10_4877_out0;
wire v$SEL10_4878_out0;
wire v$SEL10_6487_out0;
wire v$SEL10_6488_out0;
wire v$SEL10_6489_out0;
wire v$SEL10_6490_out0;
wire v$SEL10_8248_out0;
wire v$SEL10_8249_out0;
wire v$SEL10_8250_out0;
wire v$SEL10_8251_out0;
wire v$SEL10_8252_out0;
wire v$SEL10_8253_out0;
wire v$SEL10_8254_out0;
wire v$SEL10_8255_out0;
wire v$SEL10_8256_out0;
wire v$SEL10_8257_out0;
wire v$SEL10_8258_out0;
wire v$SEL10_8259_out0;
wire v$SEL10_8260_out0;
wire v$SEL10_8261_out0;
wire v$SEL10_8262_out0;
wire v$SEL10_8263_out0;
wire v$SEL10_8264_out0;
wire v$SEL10_8265_out0;
wire v$SEL10_8266_out0;
wire v$SEL10_8267_out0;
wire v$SEL10_8268_out0;
wire v$SEL10_8269_out0;
wire v$SEL10_8270_out0;
wire v$SEL10_8271_out0;
wire v$SEL10_989_out0;
wire v$SEL10_990_out0;
wire v$SEL11_10831_out0;
wire v$SEL11_10832_out0;
wire v$SEL11_11105_out0;
wire v$SEL11_11106_out0;
wire v$SEL11_4834_out0;
wire v$SEL11_4835_out0;
wire v$SEL11_4836_out0;
wire v$SEL11_4837_out0;
wire v$SEL11_5832_out0;
wire v$SEL11_5833_out0;
wire v$SEL11_729_out0;
wire v$SEL11_730_out0;
wire v$SEL11_7974_out0;
wire v$SEL11_7975_out0;
wire v$SEL12_581_out0;
wire v$SEL12_582_out0;
wire v$SEL12_741_out0;
wire v$SEL12_742_out0;
wire v$SEL12_9362_out0;
wire v$SEL12_9363_out0;
wire v$SEL12_9364_out0;
wire v$SEL12_9365_out0;
wire v$SEL13_12388_out0;
wire v$SEL13_12389_out0;
wire v$SEL13_2590_out0;
wire v$SEL13_2591_out0;
wire v$SEL13_4694_out0;
wire v$SEL13_4695_out0;
wire v$SEL13_4696_out0;
wire v$SEL13_4697_out0;
wire v$SEL14_11462_out0;
wire v$SEL14_11463_out0;
wire v$SEL14_11464_out0;
wire v$SEL14_11465_out0;
wire v$SEL14_3219_out0;
wire v$SEL14_3220_out0;
wire v$SEL15_3278_out0;
wire v$SEL15_3279_out0;
wire v$SEL15_3280_out0;
wire v$SEL15_3281_out0;
wire v$SEL15_6433_out0;
wire v$SEL15_6434_out0;
wire v$SEL15_9174_out0;
wire v$SEL15_9175_out0;
wire v$SEL16_11943_out0;
wire v$SEL16_11944_out0;
wire v$SEL16_11945_out0;
wire v$SEL16_11946_out0;
wire v$SEL17_11249_out0;
wire v$SEL17_11250_out0;
wire v$SEL17_11251_out0;
wire v$SEL17_11252_out0;
wire v$SEL18_7420_out0;
wire v$SEL18_7421_out0;
wire v$SEL18_7422_out0;
wire v$SEL18_7423_out0;
wire v$SEL19_8464_out0;
wire v$SEL19_8465_out0;
wire v$SEL19_8466_out0;
wire v$SEL19_8467_out0;
wire v$SEL1_1191_out0;
wire v$SEL1_1192_out0;
wire v$SEL1_1193_out0;
wire v$SEL1_1194_out0;
wire v$SEL1_1195_out0;
wire v$SEL1_1196_out0;
wire v$SEL1_1197_out0;
wire v$SEL1_1198_out0;
wire v$SEL1_12809_out0;
wire v$SEL1_12810_out0;
wire v$SEL1_12811_out0;
wire v$SEL1_12812_out0;
wire v$SEL1_2216_out0;
wire v$SEL1_2217_out0;
wire v$SEL1_2433_out0;
wire v$SEL1_2434_out0;
wire v$SEL1_4765_out0;
wire v$SEL1_4817_out0;
wire v$SEL1_4818_out0;
wire v$SEL1_4819_out0;
wire v$SEL1_4820_out0;
wire v$SEL1_7324_out0;
wire v$SEL1_7325_out0;
wire v$SEL1_7326_out0;
wire v$SEL1_7327_out0;
wire v$SEL1_7328_out0;
wire v$SEL1_7329_out0;
wire v$SEL1_7330_out0;
wire v$SEL1_7331_out0;
wire v$SEL1_7332_out0;
wire v$SEL1_7333_out0;
wire v$SEL1_7334_out0;
wire v$SEL1_7335_out0;
wire v$SEL1_7336_out0;
wire v$SEL1_7337_out0;
wire v$SEL1_7338_out0;
wire v$SEL1_7339_out0;
wire v$SEL1_7340_out0;
wire v$SEL1_7341_out0;
wire v$SEL1_7342_out0;
wire v$SEL1_7343_out0;
wire v$SEL1_7344_out0;
wire v$SEL1_7345_out0;
wire v$SEL1_7346_out0;
wire v$SEL1_7347_out0;
wire v$SEL1_8929_out0;
wire v$SEL1_8930_out0;
wire v$SEL1_8931_out0;
wire v$SEL1_8932_out0;
wire v$SEL1_9025_out0;
wire v$SEL1_9026_out0;
wire v$SEL1_9027_out0;
wire v$SEL1_9028_out0;
wire v$SEL1_9029_out0;
wire v$SEL1_9030_out0;
wire v$SEL1_9031_out0;
wire v$SEL1_9032_out0;
wire v$SEL1_9033_out0;
wire v$SEL1_9034_out0;
wire v$SEL1_9035_out0;
wire v$SEL1_9036_out0;
wire v$SEL1_9037_out0;
wire v$SEL1_9038_out0;
wire v$SEL1_9039_out0;
wire v$SEL1_9040_out0;
wire v$SEL1_9041_out0;
wire v$SEL1_9042_out0;
wire v$SEL1_9043_out0;
wire v$SEL1_9044_out0;
wire v$SEL1_9045_out0;
wire v$SEL1_9046_out0;
wire v$SEL1_9047_out0;
wire v$SEL1_9048_out0;
wire v$SEL1_9049_out0;
wire v$SEL1_9050_out0;
wire v$SEL1_9051_out0;
wire v$SEL1_9052_out0;
wire v$SEL1_9053_out0;
wire v$SEL1_9054_out0;
wire v$SEL1_9055_out0;
wire v$SEL1_9056_out0;
wire v$SEL1_9057_out0;
wire v$SEL1_9058_out0;
wire v$SEL1_9059_out0;
wire v$SEL1_9060_out0;
wire v$SEL1_9061_out0;
wire v$SEL1_9062_out0;
wire v$SEL1_9063_out0;
wire v$SEL1_9064_out0;
wire v$SEL1_9065_out0;
wire v$SEL1_9066_out0;
wire v$SEL1_9067_out0;
wire v$SEL1_9068_out0;
wire v$SEL1_9069_out0;
wire v$SEL1_9070_out0;
wire v$SEL1_9071_out0;
wire v$SEL1_9072_out0;
wire v$SEL1_9073_out0;
wire v$SEL1_9074_out0;
wire v$SEL1_9075_out0;
wire v$SEL1_9076_out0;
wire v$SEL1_9077_out0;
wire v$SEL1_9078_out0;
wire v$SEL1_9079_out0;
wire v$SEL1_9080_out0;
wire v$SEL1_9081_out0;
wire v$SEL1_9082_out0;
wire v$SEL1_9083_out0;
wire v$SEL1_9084_out0;
wire v$SEL20_5666_out0;
wire v$SEL20_5667_out0;
wire v$SEL20_5668_out0;
wire v$SEL20_5669_out0;
wire v$SEL21_7286_out0;
wire v$SEL21_7287_out0;
wire v$SEL21_7288_out0;
wire v$SEL21_7289_out0;
wire v$SEL22_4990_out0;
wire v$SEL22_4991_out0;
wire v$SEL22_4992_out0;
wire v$SEL22_4993_out0;
wire v$SEL23_5155_out0;
wire v$SEL23_5156_out0;
wire v$SEL23_5157_out0;
wire v$SEL23_5158_out0;
wire v$SEL24_11975_out0;
wire v$SEL24_11976_out0;
wire v$SEL24_11977_out0;
wire v$SEL24_11978_out0;
wire v$SEL27_11434_out0;
wire v$SEL27_11435_out0;
wire v$SEL27_11436_out0;
wire v$SEL27_11437_out0;
wire v$SEL28_4925_out0;
wire v$SEL28_4926_out0;
wire v$SEL28_4927_out0;
wire v$SEL28_4928_out0;
wire v$SEL29_11666_out0;
wire v$SEL29_11667_out0;
wire v$SEL29_11668_out0;
wire v$SEL29_11669_out0;
wire v$SEL2_11054_out0;
wire v$SEL2_11672_out0;
wire v$SEL2_11673_out0;
wire v$SEL2_11674_out0;
wire v$SEL2_11675_out0;
wire v$SEL2_11676_out0;
wire v$SEL2_11677_out0;
wire v$SEL2_11678_out0;
wire v$SEL2_11679_out0;
wire v$SEL2_11680_out0;
wire v$SEL2_11681_out0;
wire v$SEL2_11682_out0;
wire v$SEL2_11683_out0;
wire v$SEL2_11684_out0;
wire v$SEL2_11685_out0;
wire v$SEL2_11686_out0;
wire v$SEL2_11687_out0;
wire v$SEL2_11688_out0;
wire v$SEL2_11689_out0;
wire v$SEL2_11690_out0;
wire v$SEL2_11691_out0;
wire v$SEL2_11692_out0;
wire v$SEL2_11693_out0;
wire v$SEL2_11694_out0;
wire v$SEL2_11695_out0;
wire v$SEL2_13056_out0;
wire v$SEL2_13057_out0;
wire v$SEL2_13058_out0;
wire v$SEL2_13059_out0;
wire v$SEL2_13060_out0;
wire v$SEL2_13061_out0;
wire v$SEL2_13062_out0;
wire v$SEL2_13063_out0;
wire v$SEL2_13163_out0;
wire v$SEL2_13164_out0;
wire v$SEL2_13165_out0;
wire v$SEL2_13166_out0;
wire v$SEL2_2427_out0;
wire v$SEL2_2428_out0;
wire v$SEL2_5201_out0;
wire v$SEL2_5202_out0;
wire v$SEL2_5203_out0;
wire v$SEL2_5204_out0;
wire v$SEL2_5205_out0;
wire v$SEL2_5206_out0;
wire v$SEL2_5207_out0;
wire v$SEL2_5208_out0;
wire v$SEL2_5209_out0;
wire v$SEL2_5210_out0;
wire v$SEL2_5211_out0;
wire v$SEL2_5212_out0;
wire v$SEL2_5213_out0;
wire v$SEL2_5214_out0;
wire v$SEL2_5215_out0;
wire v$SEL2_5216_out0;
wire v$SEL2_5217_out0;
wire v$SEL2_5218_out0;
wire v$SEL2_5219_out0;
wire v$SEL2_5220_out0;
wire v$SEL2_5221_out0;
wire v$SEL2_5222_out0;
wire v$SEL2_5223_out0;
wire v$SEL2_5224_out0;
wire v$SEL2_5225_out0;
wire v$SEL2_5226_out0;
wire v$SEL2_5227_out0;
wire v$SEL2_5228_out0;
wire v$SEL2_5229_out0;
wire v$SEL2_5230_out0;
wire v$SEL2_5231_out0;
wire v$SEL2_5232_out0;
wire v$SEL2_5233_out0;
wire v$SEL2_5234_out0;
wire v$SEL2_5235_out0;
wire v$SEL2_5236_out0;
wire v$SEL2_5237_out0;
wire v$SEL2_5238_out0;
wire v$SEL2_5239_out0;
wire v$SEL2_5240_out0;
wire v$SEL2_5241_out0;
wire v$SEL2_5242_out0;
wire v$SEL2_5243_out0;
wire v$SEL2_5244_out0;
wire v$SEL2_5245_out0;
wire v$SEL2_5246_out0;
wire v$SEL2_5247_out0;
wire v$SEL2_5248_out0;
wire v$SEL2_5249_out0;
wire v$SEL2_5250_out0;
wire v$SEL2_5251_out0;
wire v$SEL2_5252_out0;
wire v$SEL2_5253_out0;
wire v$SEL2_5254_out0;
wire v$SEL2_5255_out0;
wire v$SEL2_5256_out0;
wire v$SEL2_5257_out0;
wire v$SEL2_5258_out0;
wire v$SEL2_5259_out0;
wire v$SEL2_5260_out0;
wire v$SEL2_6423_out0;
wire v$SEL2_6424_out0;
wire v$SEL2_7442_out0;
wire v$SEL2_7443_out0;
wire v$SEL2_7444_out0;
wire v$SEL2_7445_out0;
wire v$SEL2_7446_out0;
wire v$SEL2_7447_out0;
wire v$SEL2_7448_out0;
wire v$SEL2_7449_out0;
wire v$SEL2_7450_out0;
wire v$SEL2_7451_out0;
wire v$SEL2_7452_out0;
wire v$SEL2_7453_out0;
wire v$SEL2_7454_out0;
wire v$SEL2_7455_out0;
wire v$SEL2_7456_out0;
wire v$SEL2_7457_out0;
wire v$SEL2_7458_out0;
wire v$SEL2_7459_out0;
wire v$SEL2_7460_out0;
wire v$SEL2_7461_out0;
wire v$SEL2_7462_out0;
wire v$SEL2_7463_out0;
wire v$SEL2_8895_out0;
wire v$SEL2_8896_out0;
wire v$SEL2_8897_out0;
wire v$SEL2_8898_out0;
wire v$SEL2_9004_out0;
wire v$SEL2_9005_out0;
wire v$SEL2_9793_out0;
wire v$SEL2_9794_out0;
wire v$SEL3_1217_out0;
wire v$SEL3_1218_out0;
wire v$SEL3_1219_out0;
wire v$SEL3_12208_out0;
wire v$SEL3_12209_out0;
wire v$SEL3_1220_out0;
wire v$SEL3_1221_out0;
wire v$SEL3_1222_out0;
wire v$SEL3_1223_out0;
wire v$SEL3_1224_out0;
wire v$SEL3_1225_out0;
wire v$SEL3_1226_out0;
wire v$SEL3_1227_out0;
wire v$SEL3_1228_out0;
wire v$SEL3_1229_out0;
wire v$SEL3_1230_out0;
wire v$SEL3_1231_out0;
wire v$SEL3_1232_out0;
wire v$SEL3_1233_out0;
wire v$SEL3_1234_out0;
wire v$SEL3_1235_out0;
wire v$SEL3_1236_out0;
wire v$SEL3_1237_out0;
wire v$SEL3_1238_out0;
wire v$SEL3_1239_out0;
wire v$SEL3_1240_out0;
wire v$SEL3_1241_out0;
wire v$SEL3_1242_out0;
wire v$SEL3_1243_out0;
wire v$SEL3_1244_out0;
wire v$SEL3_1245_out0;
wire v$SEL3_1246_out0;
wire v$SEL3_1247_out0;
wire v$SEL3_1248_out0;
wire v$SEL3_1249_out0;
wire v$SEL3_1250_out0;
wire v$SEL3_1251_out0;
wire v$SEL3_1252_out0;
wire v$SEL3_1253_out0;
wire v$SEL3_1254_out0;
wire v$SEL3_1255_out0;
wire v$SEL3_1256_out0;
wire v$SEL3_1257_out0;
wire v$SEL3_1258_out0;
wire v$SEL3_1259_out0;
wire v$SEL3_1260_out0;
wire v$SEL3_1261_out0;
wire v$SEL3_1262_out0;
wire v$SEL3_1263_out0;
wire v$SEL3_1264_out0;
wire v$SEL3_1265_out0;
wire v$SEL3_1266_out0;
wire v$SEL3_1267_out0;
wire v$SEL3_1268_out0;
wire v$SEL3_1269_out0;
wire v$SEL3_1270_out0;
wire v$SEL3_1271_out0;
wire v$SEL3_1272_out0;
wire v$SEL3_1273_out0;
wire v$SEL3_1274_out0;
wire v$SEL3_1275_out0;
wire v$SEL3_1276_out0;
wire v$SEL3_1872_out0;
wire v$SEL3_437_out0;
wire v$SEL3_438_out0;
wire v$SEL3_439_out0;
wire v$SEL3_440_out0;
wire v$SEL3_441_out0;
wire v$SEL3_442_out0;
wire v$SEL3_443_out0;
wire v$SEL3_444_out0;
wire v$SEL3_5880_out0;
wire v$SEL3_5881_out0;
wire v$SEL3_5882_out0;
wire v$SEL3_5883_out0;
wire v$SEL3_5884_out0;
wire v$SEL3_5885_out0;
wire v$SEL3_5886_out0;
wire v$SEL3_5887_out0;
wire v$SEL3_5888_out0;
wire v$SEL3_5889_out0;
wire v$SEL3_5890_out0;
wire v$SEL3_5891_out0;
wire v$SEL3_5892_out0;
wire v$SEL3_5893_out0;
wire v$SEL3_5894_out0;
wire v$SEL3_5895_out0;
wire v$SEL3_5896_out0;
wire v$SEL3_5897_out0;
wire v$SEL3_5898_out0;
wire v$SEL3_5899_out0;
wire v$SEL3_5900_out0;
wire v$SEL3_5901_out0;
wire v$SEL3_5902_out0;
wire v$SEL3_5903_out0;
wire v$SEL3_7544_out0;
wire v$SEL3_7545_out0;
wire v$SEL3_7546_out0;
wire v$SEL3_7547_out0;
wire v$SEL3_887_out0;
wire v$SEL3_888_out0;
wire v$SEL3_9405_out0;
wire v$SEL3_9406_out0;
wire v$SEL3_9407_out0;
wire v$SEL3_9408_out0;
wire v$SEL4_1017_out0;
wire v$SEL4_1018_out0;
wire v$SEL4_1019_out0;
wire v$SEL4_1020_out0;
wire v$SEL4_11518_out0;
wire v$SEL4_3330_out0;
wire v$SEL4_3331_out0;
wire v$SEL4_3332_out0;
wire v$SEL4_3333_out0;
wire v$SEL4_3334_out0;
wire v$SEL4_3335_out0;
wire v$SEL4_3336_out0;
wire v$SEL4_3337_out0;
wire v$SEL4_4081_out0;
wire v$SEL4_4082_out0;
wire v$SEL4_4083_out0;
wire v$SEL4_4084_out0;
wire v$SEL4_4085_out0;
wire v$SEL4_4086_out0;
wire v$SEL4_4087_out0;
wire v$SEL4_4088_out0;
wire v$SEL4_4089_out0;
wire v$SEL4_4090_out0;
wire v$SEL4_4091_out0;
wire v$SEL4_4092_out0;
wire v$SEL4_4093_out0;
wire v$SEL4_4094_out0;
wire v$SEL4_4095_out0;
wire v$SEL4_4096_out0;
wire v$SEL4_4097_out0;
wire v$SEL4_4098_out0;
wire v$SEL4_4099_out0;
wire v$SEL4_4100_out0;
wire v$SEL4_4101_out0;
wire v$SEL4_4102_out0;
wire v$SEL4_4103_out0;
wire v$SEL4_4104_out0;
wire v$SEL4_4105_out0;
wire v$SEL4_4106_out0;
wire v$SEL4_4107_out0;
wire v$SEL4_4108_out0;
wire v$SEL4_4109_out0;
wire v$SEL4_4110_out0;
wire v$SEL4_4111_out0;
wire v$SEL4_4112_out0;
wire v$SEL4_4113_out0;
wire v$SEL4_4114_out0;
wire v$SEL4_4115_out0;
wire v$SEL4_4116_out0;
wire v$SEL4_4117_out0;
wire v$SEL4_4118_out0;
wire v$SEL4_4119_out0;
wire v$SEL4_4120_out0;
wire v$SEL4_4121_out0;
wire v$SEL4_4122_out0;
wire v$SEL4_4123_out0;
wire v$SEL4_4124_out0;
wire v$SEL4_4125_out0;
wire v$SEL4_4126_out0;
wire v$SEL4_4127_out0;
wire v$SEL4_4128_out0;
wire v$SEL4_4129_out0;
wire v$SEL4_4130_out0;
wire v$SEL4_4131_out0;
wire v$SEL4_4132_out0;
wire v$SEL4_4133_out0;
wire v$SEL4_4134_out0;
wire v$SEL4_4135_out0;
wire v$SEL4_4136_out0;
wire v$SEL4_4137_out0;
wire v$SEL4_4138_out0;
wire v$SEL4_4139_out0;
wire v$SEL4_4140_out0;
wire v$SEL4_475_out0;
wire v$SEL4_476_out0;
wire v$SEL4_4802_out0;
wire v$SEL4_4803_out0;
wire v$SEL4_4919_out0;
wire v$SEL4_4920_out0;
wire v$SEL4_4921_out0;
wire v$SEL4_4922_out0;
wire v$SEL4_4932_out0;
wire v$SEL4_4933_out0;
wire v$SEL4_4934_out0;
wire v$SEL4_4935_out0;
wire v$SEL4_4936_out0;
wire v$SEL4_4937_out0;
wire v$SEL4_4938_out0;
wire v$SEL4_4939_out0;
wire v$SEL4_4940_out0;
wire v$SEL4_4941_out0;
wire v$SEL4_4942_out0;
wire v$SEL4_4943_out0;
wire v$SEL4_4944_out0;
wire v$SEL4_4945_out0;
wire v$SEL4_4946_out0;
wire v$SEL4_4947_out0;
wire v$SEL4_4948_out0;
wire v$SEL4_4949_out0;
wire v$SEL4_4950_out0;
wire v$SEL4_4951_out0;
wire v$SEL4_4952_out0;
wire v$SEL4_4953_out0;
wire v$SEL4_4954_out0;
wire v$SEL4_4955_out0;
wire v$SEL5_10744_out0;
wire v$SEL5_10745_out0;
wire v$SEL5_10746_out0;
wire v$SEL5_10747_out0;
wire v$SEL5_260_out0;
wire v$SEL5_261_out0;
wire v$SEL5_7466_out0;
wire v$SEL5_7496_out0;
wire v$SEL5_7497_out0;
wire v$SEL5_7498_out0;
wire v$SEL5_7499_out0;
wire v$SEL5_783_out0;
wire v$SEL5_784_out0;
wire v$SEL5_7988_out0;
wire v$SEL5_7989_out0;
wire v$SEL5_7990_out0;
wire v$SEL5_7991_out0;
wire v$SEL5_7992_out0;
wire v$SEL5_7993_out0;
wire v$SEL5_7994_out0;
wire v$SEL5_7995_out0;
wire v$SEL5_8430_out0;
wire v$SEL5_8431_out0;
wire v$SEL5_8432_out0;
wire v$SEL5_8433_out0;
wire v$SEL5_8434_out0;
wire v$SEL5_8435_out0;
wire v$SEL5_8436_out0;
wire v$SEL5_8437_out0;
wire v$SEL5_8438_out0;
wire v$SEL5_8439_out0;
wire v$SEL5_8440_out0;
wire v$SEL5_8441_out0;
wire v$SEL5_8442_out0;
wire v$SEL5_8443_out0;
wire v$SEL5_8444_out0;
wire v$SEL5_8445_out0;
wire v$SEL5_8446_out0;
wire v$SEL5_8447_out0;
wire v$SEL5_8448_out0;
wire v$SEL5_8449_out0;
wire v$SEL5_8450_out0;
wire v$SEL5_8451_out0;
wire v$SEL5_8452_out0;
wire v$SEL5_8453_out0;
wire v$SEL6_3825_out0;
wire v$SEL6_3826_out0;
wire v$SEL6_3827_out0;
wire v$SEL6_3828_out0;
wire v$SEL6_6178_out0;
wire v$SEL6_6179_out0;
wire v$SEL6_6180_out0;
wire v$SEL6_6181_out0;
wire v$SEL6_8113_out0;
wire v$SEL6_8114_out0;
wire v$SEL6_8115_out0;
wire v$SEL6_8116_out0;
wire v$SEL6_9304_out0;
wire v$SEL6_9305_out0;
wire v$SEL6_9306_out0;
wire v$SEL6_9307_out0;
wire v$SEL6_9308_out0;
wire v$SEL6_9309_out0;
wire v$SEL6_9310_out0;
wire v$SEL6_9311_out0;
wire v$SEL6_9641_out0;
wire v$SEL6_9839_out0;
wire v$SEL6_9840_out0;
wire v$SEL7_10884_out0;
wire v$SEL7_10885_out0;
wire v$SEL7_12068_out0;
wire v$SEL7_2856_out0;
wire v$SEL7_2857_out0;
wire v$SEL7_2858_out0;
wire v$SEL7_2859_out0;
wire v$SEL7_2860_out0;
wire v$SEL7_2861_out0;
wire v$SEL7_2862_out0;
wire v$SEL7_2863_out0;
wire v$SEL7_2864_out0;
wire v$SEL7_2865_out0;
wire v$SEL7_2866_out0;
wire v$SEL7_2867_out0;
wire v$SEL7_2868_out0;
wire v$SEL7_2869_out0;
wire v$SEL7_2870_out0;
wire v$SEL7_2871_out0;
wire v$SEL7_2872_out0;
wire v$SEL7_2873_out0;
wire v$SEL7_2874_out0;
wire v$SEL7_2875_out0;
wire v$SEL7_2876_out0;
wire v$SEL7_2877_out0;
wire v$SEL7_2878_out0;
wire v$SEL7_2879_out0;
wire v$SEL7_4357_out0;
wire v$SEL7_4358_out0;
wire v$SEL7_4359_out0;
wire v$SEL7_4360_out0;
wire v$SEL7_4361_out0;
wire v$SEL7_4362_out0;
wire v$SEL7_4363_out0;
wire v$SEL7_4364_out0;
wire v$SEL7_491_out0;
wire v$SEL7_492_out0;
wire v$SEL7_9719_out0;
wire v$SEL7_9720_out0;
wire v$SEL7_9721_out0;
wire v$SEL7_9722_out0;
wire v$SEL8_1110_out0;
wire v$SEL8_11646_out0;
wire v$SEL8_11647_out0;
wire v$SEL8_11648_out0;
wire v$SEL8_11649_out0;
wire v$SEL8_11650_out0;
wire v$SEL8_11651_out0;
wire v$SEL8_11652_out0;
wire v$SEL8_11653_out0;
wire v$SEL8_12507_out0;
wire v$SEL8_12508_out0;
wire v$SEL8_12509_out0;
wire v$SEL8_12510_out0;
wire v$SEL8_8559_out0;
wire v$SEL8_8560_out0;
wire v$SEL8_8561_out0;
wire v$SEL8_8562_out0;
wire v$SEL8_8563_out0;
wire v$SEL8_8564_out0;
wire v$SEL8_8565_out0;
wire v$SEL8_8566_out0;
wire v$SEL8_8567_out0;
wire v$SEL8_8568_out0;
wire v$SEL8_8569_out0;
wire v$SEL8_8570_out0;
wire v$SEL8_8571_out0;
wire v$SEL8_8572_out0;
wire v$SEL8_8573_out0;
wire v$SEL8_8574_out0;
wire v$SEL8_8575_out0;
wire v$SEL8_8576_out0;
wire v$SEL8_8577_out0;
wire v$SEL8_8578_out0;
wire v$SEL8_8579_out0;
wire v$SEL8_8580_out0;
wire v$SEL8_8581_out0;
wire v$SEL8_8582_out0;
wire v$SEL9_3639_out0;
wire v$SEL9_3640_out0;
wire v$SEL9_6829_out0;
wire v$SEL9_6830_out0;
wire v$SEL9_6831_out0;
wire v$SEL9_6832_out0;
wire v$SEL9_7128_out0;
wire v$SEL9_7129_out0;
wire v$SEL9_7130_out0;
wire v$SEL9_7131_out0;
wire v$SEL9_7132_out0;
wire v$SEL9_7133_out0;
wire v$SEL9_7134_out0;
wire v$SEL9_7135_out0;
wire v$SEL9_7136_out0;
wire v$SEL9_7137_out0;
wire v$SEL9_7138_out0;
wire v$SEL9_7139_out0;
wire v$SEL9_7140_out0;
wire v$SEL9_7141_out0;
wire v$SEL9_7142_out0;
wire v$SEL9_7143_out0;
wire v$SEL9_7144_out0;
wire v$SEL9_7145_out0;
wire v$SEL9_7146_out0;
wire v$SEL9_7147_out0;
wire v$SEL9_7148_out0;
wire v$SEL9_7149_out0;
wire v$SEL9_7150_out0;
wire v$SEL9_7151_out0;
wire v$SELIN$VIEWER_7303_out0;
wire v$SELIN_12946_out0;
wire v$SELOUTVIEWER_4876_out0;
wire v$SELOUT_900_out0;
wire v$SERIALIN_3766_out0;
wire v$SERIALIN_3767_out0;
wire v$SHIFTEN_4821_out0;
wire v$SHIFTEN_4822_out0;
wire v$SHIFTEN_6401_out0;
wire v$SHIFTEN_6402_out0;
wire v$SHIFTEN_6403_out0;
wire v$SHIFTEN_6404_out0;
wire v$SHIFTEN_6405_out0;
wire v$SHIFTEN_6406_out0;
wire v$SHIFTEN_6407_out0;
wire v$SHIFTEN_6408_out0;
wire v$SHIFTEN_6409_out0;
wire v$SHIFTEN_6410_out0;
wire v$SHIFTEN_6411_out0;
wire v$SHIFTEN_6412_out0;
wire v$SHIFTEN_6847_out0;
wire v$SHIFTEN_6848_out0;
wire v$SHIFTEN_8420_out0;
wire v$SHIFTEN_8421_out0;
wire v$SIGN_591_out0;
wire v$SIGN_592_out0;
wire v$SIGN_593_out0;
wire v$SIGN_594_out0;
wire v$SIGN_8414_out0;
wire v$SIGN_8415_out0;
wire v$SIN_84_out0;
wire v$SIN_85_out0;
wire v$SIN_86_out0;
wire v$SIN_87_out0;
wire v$SIN_88_out0;
wire v$SIN_89_out0;
wire v$SIN_90_out0;
wire v$SIN_91_out0;
wire v$SIN_92_out0;
wire v$SIN_93_out0;
wire v$SIN_94_out0;
wire v$SIN_95_out0;
wire v$SOUT1_1068_out0;
wire v$SOUT1_1069_out0;
wire v$SOUT1_1070_out0;
wire v$SOUT1_1071_out0;
wire v$SOUT1_1072_out0;
wire v$SOUT1_1073_out0;
wire v$SOUT1_1074_out0;
wire v$SOUT1_1075_out0;
wire v$SOUT1_1076_out0;
wire v$SOUT1_1077_out0;
wire v$SOUT1_1078_out0;
wire v$SOUT1_1079_out0;
wire v$SOUT_12929_out0;
wire v$SOUT_12930_out0;
wire v$STALL$FETCH$OCCURRED_1549_out0;
wire v$STALL$FETCH$OCCURRED_1550_out0;
wire v$STALL$IN$PREV_8808_out0;
wire v$STALL$IN$PREV_8809_out0;
wire v$STALL$PREV$CYCLE_3798_out0;
wire v$STALL$PREV$CYCLE_3799_out0;
wire v$STALL$PREV$PREV_3829_out0;
wire v$STALL$PREV$PREV_3830_out0;
wire v$STALL$VIEWER_12825_out0;
wire v$STALL$VIEWER_12826_out0;
wire v$STALL_10775_out0;
wire v$STALL_10776_out0;
wire v$STALL_12672_out0;
wire v$STALL_12673_out0;
wire v$STALL_8002_out0;
wire v$STALL_8003_out0;
wire v$STALL_8758_out0;
wire v$STALL_8759_out0;
wire v$STATE_11196_out0;
wire v$STATE_11197_out0;
wire v$STATE_11198_out0;
wire v$STATUSCLR_3955_out0;
wire v$STATUSCLR_3956_out0;
wire v$STATUSREAD_835_out0;
wire v$STATUSREAD_836_out0;
wire v$STClr_6793_out0;
wire v$STClr_6794_out0;
wire v$STOP$1_5336_out0;
wire v$STOP$1_5337_out0;
wire v$STOP$2_5722_out0;
wire v$STOP$2_5723_out0;
wire v$STOPBITERROR_7542_out0;
wire v$STOPBITERROR_7543_out0;
wire v$STOPERROR_246_out0;
wire v$STOPERROR_247_out0;
wire v$STP$DECODED_11614_out0;
wire v$STP$DECODED_11615_out0;
wire v$STP$SAVED_5106_out0;
wire v$STP$SAVED_5107_out0;
wire v$STPHALT_12859_out0;
wire v$STPHALT_12860_out0;
wire v$STPHALT_2988_out0;
wire v$STPHALT_2989_out0;
wire v$STPHALT_8583_out0;
wire v$STPHALT_8584_out0;
wire v$STP_12552_out0;
wire v$STP_12553_out0;
wire v$STP_4222_out0;
wire v$STP_4223_out0;
wire v$STP_7120_out0;
wire v$STP_7121_out0;
wire v$STP_7534_out0;
wire v$STP_7535_out0;
wire v$STRead_6652_out0;
wire v$STRead_6653_out0;
wire v$SUBEN_8502_out0;
wire v$SUBEN_8503_out0;
wire v$SUBTRACTION$SIGN_7667_out0;
wire v$SUBTRACTION$SIGN_7668_out0;
wire v$SUB_9314_out0;
wire v$SUB_9315_out0;
wire v$SUM$0_8097_out0;
wire v$SUM$0_8098_out0;
wire v$SUM$10_9699_out0;
wire v$SUM$10_9700_out0;
wire v$SUM$11_12086_out0;
wire v$SUM$11_12087_out0;
wire v$SUM$1_6901_out0;
wire v$SUM$1_6902_out0;
wire v$SUM$2_6320_out0;
wire v$SUM$2_6321_out0;
wire v$SUM$3_5420_out0;
wire v$SUM$3_5421_out0;
wire v$SUM$4_10567_out0;
wire v$SUM$4_10568_out0;
wire v$SUM$5_5344_out0;
wire v$SUM$5_5345_out0;
wire v$SUM$6_8556_out0;
wire v$SUM$6_8557_out0;
wire v$SUM$7_5287_out0;
wire v$SUM$7_5288_out0;
wire v$SUM$8_11009_out0;
wire v$SUM$8_11010_out0;
wire v$SUM$9_184_out0;
wire v$SUM$9_185_out0;
wire v$S_10768_out0;
wire v$S_10769_out0;
wire v$S_11488_out0;
wire v$S_11489_out0;
wire v$S_11983_out0;
wire v$S_11984_out0;
wire v$S_11985_out0;
wire v$S_11986_out0;
wire v$S_11987_out0;
wire v$S_11988_out0;
wire v$S_11989_out0;
wire v$S_11990_out0;
wire v$S_11991_out0;
wire v$S_11992_out0;
wire v$S_11993_out0;
wire v$S_11994_out0;
wire v$S_11995_out0;
wire v$S_11996_out0;
wire v$S_11997_out0;
wire v$S_11998_out0;
wire v$S_11999_out0;
wire v$S_12000_out0;
wire v$S_12001_out0;
wire v$S_12002_out0;
wire v$S_12003_out0;
wire v$S_12004_out0;
wire v$S_12723_out0;
wire v$S_12724_out0;
wire v$S_1371_out0;
wire v$S_1372_out0;
wire v$S_2742_out0;
wire v$S_2743_out0;
wire v$S_2914_out0;
wire v$S_2915_out0;
wire v$S_3770_out0;
wire v$S_3771_out0;
wire v$S_406_out0;
wire v$S_407_out0;
wire v$S_495_out0;
wire v$S_5522_out0;
wire v$S_5523_out0;
wire v$S_5524_out0;
wire v$S_5664_out0;
wire v$S_5665_out0;
wire v$S_6419_out0;
wire v$S_6420_out0;
wire v$S_6897_out0;
wire v$S_6898_out0;
wire v$S_6988_out0;
wire v$S_6989_out0;
wire v$S_7016_out0;
wire v$S_7017_out0;
wire v$S_8290_out0;
wire v$S_8291_out0;
wire v$S_8468_out0;
wire v$S_8469_out0;
wire v$SetError_12380_out0;
wire v$SetError_12381_out0;
wire v$ShiftEN_3842_out0;
wire v$ShiftEN_3843_out0;
wire v$ShiftEN_5265_out0;
wire v$ShiftEN_5266_out0;
wire v$ShiftOut_11458_out0;
wire v$ShiftOut_11459_out0;
wire v$Shift_6566_out0;
wire v$Shift_6567_out0;
wire v$StatRegAdd1_9943_out0;
wire v$StatRegAdd1_9944_out0;
wire v$StatRegAdd_5285_out0;
wire v$StatRegAdd_5286_out0;
wire v$TAKEJUMP_7106_out0;
wire v$TAKEJUMP_7107_out0;
wire v$THRESHOLD$WRITE_4845_out0;
wire v$THRESHOLD$WRITE_4846_out0;
wire v$TWOS$COMPLEMENT$ADDER$COUT_2137_out0;
wire v$TWOS$COMPLEMENT$ADDER$COUT_2138_out0;
wire v$TXFLAG_10050_out0;
wire v$TXFLAG_10051_out0;
wire v$TXFLAG_2586_out0;
wire v$TXFLAG_2587_out0;
wire v$TXFlag_10569_out0;
wire v$TXFlag_10570_out0;
wire v$TXFlag_5261_out0;
wire v$TXFlag_5262_out0;
wire v$TXINTERRUPT_2342_out0;
wire v$TXINTERRUPT_2343_out0;
wire v$TXINT_3304_out0;
wire v$TXINT_3305_out0;
wire v$TXLast_7426_out0;
wire v$TXLast_7427_out0;
wire v$TXRST_11484_out0;
wire v$TXRST_11485_out0;
wire v$TXRST_5553_out0;
wire v$TXRST_5554_out0;
wire v$TXRegAdd_10869_out0;
wire v$TXRegAdd_10870_out0;
wire v$TXReset_12625_out0;
wire v$TXReset_12626_out0;
wire v$TXSet_8294_out0;
wire v$TXSet_8295_out0;
wire v$TXSet_9724_out0;
wire v$TXSet_9725_out0;
wire v$TXWRITE_11277_out0;
wire v$TXWRITE_11278_out0;
wire v$TXWRITE_7348_out0;
wire v$TXWRITE_7349_out0;
wire v$TXWrite_12290_out0;
wire v$TXWrite_12291_out0;
wire v$TX_12978_out0;
wire v$TX_12979_out0;
wire v$TX_349_out0;
wire v$TX_350_out0;
wire v$TX_534_out0;
wire v$TX_535_out0;
wire v$TX_7506_out0;
wire v$TX_7507_out0;
wire v$TXoverflow_2807_out0;
wire v$TXoverflow_2808_out0;
wire v$V0_5005_out0;
wire v$V0_6376_out0;
wire v$V1_11769_out0;
wire v$V1_12627_out0;
wire v$VALID$PREV_9000_out0;
wire v$VALID$PREV_9001_out0;
wire v$VALID0_8975_out0;
wire v$VALID1_6051_out0;
wire v$VALID_12693_out0;
wire v$VALID_12694_out0;
wire v$VALID_13300_out0;
wire v$VALID_13301_out0;
wire v$VALID_2425_out0;
wire v$VALID_2426_out0;
wire v$VALID_9883_out0;
wire v$VALID_9884_out0;
wire v$WB$HAZARD_6143_out0;
wire v$WB$HAZARD_6144_out0;
wire v$WEN$FPU_5786_out0;
wire v$WEN$FPU_5787_out0;
wire v$WEN3_1021_out0;
wire v$WEN3_1022_out0;
wire v$WEN3_1983_out0;
wire v$WEN3_1984_out0;
wire v$WENALU_11482_out0;
wire v$WENALU_11483_out0;
wire v$WENALU_13296_out0;
wire v$WENALU_13297_out0;
wire v$WENALU_2782_out0;
wire v$WENALU_2783_out0;
wire v$WENFPU_2200_out0;
wire v$WENFPU_2201_out0;
wire v$WENFPU_9279_out0;
wire v$WENFPU_9280_out0;
wire v$WENLDST_13265_out0;
wire v$WENLDST_13266_out0;
wire v$WENLDST_4677_out0;
wire v$WENLDST_4678_out0;
wire v$WENLDST_8125_out0;
wire v$WENLDST_8126_out0;
wire v$WENRAM0_6651_out0;
wire v$WENRAM1_899_out0;
wire v$WENRAM_12116_out0;
wire v$WENRAM_12117_out0;
wire v$WENRAM_1277_out0;
wire v$WENRAM_1278_out0;
wire v$WENRAM_3362_out0;
wire v$WENRAM_3363_out0;
wire v$WEN_13084_out0;
wire v$WEN_13085_out0;
wire v$WEN_2398_out0;
wire v$WEN_2399_out0;
wire v$WEN_2509_out0;
wire v$WEN_2510_out0;
wire v$WEN_7946_out0;
wire v$WEN_7947_out0;
wire v$WEN_8101_out0;
wire v$WEN_8102_out0;
wire v$WEN_9615_out0;
wire v$WEN_9616_out0;
wire v$WR0VIEWER_11107_out0;
wire v$WR0_546_out0;
wire v$WR0_9664_out0;
wire v$WR1VIEWER_11120_out0;
wire v$WR1_255_out0;
wire v$WR1_9723_out0;
wire v$WREN_1443_out0;
wire v$WREN_1444_out0;
wire v$WREN_7251_out0;
wire v$WREN_7252_out0;
wire v$Wordlength_3514_out0;
wire v$Wordlength_3515_out0;
wire v$Write_1959_out0;
wire v$Write_1960_out0;
wire v$Write_1961_out0;
wire v$Write_1962_out0;
wire v$Write_1963_out0;
wire v$Write_1964_out0;
wire v$Write_1965_out0;
wire v$Write_1966_out0;
wire v$Write_1967_out0;
wire v$Write_1968_out0;
wire v$Write_1969_out0;
wire v$Write_1970_out0;
wire v$Z1_12048_out0;
wire v$Z1_12049_out0;
wire v$Z1_12050_out0;
wire v$Z1_12051_out0;
wire v$Z1_12052_out0;
wire v$Z1_12053_out0;
wire v$Z1_12054_out0;
wire v$Z1_12055_out0;
wire v$Z1_12056_out0;
wire v$Z1_12057_out0;
wire v$Z1_12058_out0;
wire v$Z1_12059_out0;
wire v$Z1_12060_out0;
wire v$Z1_12061_out0;
wire v$Z1_12062_out0;
wire v$Z1_12063_out0;
wire v$Z1_12534_out0;
wire v$Z1_12535_out0;
wire v$Z1_3792_out0;
wire v$Z1_3793_out0;
wire v$Z1_3794_out0;
wire v$Z1_3795_out0;
wire v$Z1_3796_out0;
wire v$Z1_3797_out0;
wire v$Z2_1177_out0;
wire v$Z2_1178_out0;
wire v$Z2_168_out0;
wire v$Z2_169_out0;
wire v$Z2_170_out0;
wire v$Z2_171_out0;
wire v$Z2_172_out0;
wire v$Z2_173_out0;
wire v$Z2_4333_out0;
wire v$Z2_4334_out0;
wire v$Z2_4335_out0;
wire v$Z2_4336_out0;
wire v$Z2_4337_out0;
wire v$Z2_4338_out0;
wire v$Z2_4339_out0;
wire v$Z2_4340_out0;
wire v$Z2_4341_out0;
wire v$Z2_4342_out0;
wire v$Z2_4343_out0;
wire v$Z2_4344_out0;
wire v$Z2_4345_out0;
wire v$Z2_4346_out0;
wire v$Z2_4347_out0;
wire v$Z2_4348_out0;
wire v$Z3_12567_out0;
wire v$Z3_12568_out0;
wire v$Z3_12569_out0;
wire v$Z3_12570_out0;
wire v$Z3_12571_out0;
wire v$Z3_12572_out0;
wire v$Z3_12573_out0;
wire v$Z3_12574_out0;
wire v$Z3_12575_out0;
wire v$Z3_12576_out0;
wire v$Z3_12577_out0;
wire v$Z3_12578_out0;
wire v$Z3_12579_out0;
wire v$Z3_12580_out0;
wire v$Z3_12581_out0;
wire v$Z3_12582_out0;
wire v$Z3_7758_out0;
wire v$Z3_7759_out0;
wire v$Z4_5426_out0;
wire v$Z4_5427_out0;
wire v$Z4_5428_out0;
wire v$Z4_5429_out0;
wire v$Z4_5430_out0;
wire v$Z4_5431_out0;
wire v$Z4_5432_out0;
wire v$Z4_5433_out0;
wire v$Z4_5434_out0;
wire v$Z4_5435_out0;
wire v$Z4_5436_out0;
wire v$Z4_5437_out0;
wire v$Z_11031_out0;
wire v$Z_11032_out0;
wire v$Z_11033_out0;
wire v$Z_11034_out0;
wire v$Z_1460_out0;
wire v$Z_1461_out0;
wire v$Z_1462_out0;
wire v$Z_1463_out0;
wire v$Z_1464_out0;
wire v$Z_1465_out0;
wire v$Z_1466_out0;
wire v$Z_1467_out0;
wire v$Z_1468_out0;
wire v$Z_1469_out0;
wire v$Z_1470_out0;
wire v$Z_1471_out0;
wire v$Z_1472_out0;
wire v$Z_1473_out0;
wire v$Z_1474_out0;
wire v$Z_1475_out0;
wire v$Z_6883_out0;
wire v$Z_6884_out0;
wire v$Z_6885_out0;
wire v$Z_6886_out0;
wire v$Z_6887_out0;
wire v$Z_6888_out0;
wire v$Z_8188_out0;
wire v$Z_8189_out0;
wire v$Z_8190_out0;
wire v$Z_8191_out0;
wire v$Z_8192_out0;
wire v$Z_8193_out0;
wire v$Z_8194_out0;
wire v$Z_8195_out0;
wire v$Z_8196_out0;
wire v$Z_8197_out0;
wire v$Z_8198_out0;
wire v$Z_8199_out0;
wire v$Z_8200_out0;
wire v$Z_8201_out0;
wire v$Z_8202_out0;
wire v$Z_8203_out0;
wire v$Z_8204_out0;
wire v$Z_8205_out0;
wire v$Z_8206_out0;
wire v$Z_8207_out0;
wire v$Z_8208_out0;
wire v$Z_8209_out0;
wire v$Z_8210_out0;
wire v$Z_8211_out0;
wire v$Z_8212_out0;
wire v$Z_8213_out0;
wire v$Z_8214_out0;
wire v$Z_8215_out0;
wire v$Z_8216_out0;
wire v$Z_8217_out0;
wire v$Z_8218_out0;
wire v$Z_8219_out0;
wire v$Z_8220_out0;
wire v$Z_8221_out0;
wire v$Z_8222_out0;
wire v$Z_8223_out0;
wire v$Z_8224_out0;
wire v$Z_8225_out0;
wire v$Z_8226_out0;
wire v$Z_8227_out0;
wire v$Z_8228_out0;
wire v$Z_8229_out0;
wire v$Z_8230_out0;
wire v$Z_8231_out0;
wire v$Z_8232_out0;
wire v$Z_8233_out0;
wire v$Z_8234_out0;
wire v$Z_8235_out0;
wire v$Z_8236_out0;
wire v$Z_8237_out0;
wire v$Z_8238_out0;
wire v$Z_8239_out0;
wire v$Z_8240_out0;
wire v$Z_8241_out0;
wire v$Z_8242_out0;
wire v$Z_8243_out0;
wire v$Z_8244_out0;
wire v$Z_8245_out0;
wire v$Z_8246_out0;
wire v$Z_8247_out0;
wire v$Z_9121_out0;
wire v$Z_9122_out0;
wire v$_10014_out0;
wire v$_10014_out1;
wire v$_10015_out0;
wire v$_10015_out1;
wire v$_10441_out0;
wire v$_10442_out0;
wire v$_10491_out0;
wire v$_10491_out1;
wire v$_10492_out0;
wire v$_10492_out1;
wire v$_10493_out0;
wire v$_10493_out1;
wire v$_10494_out0;
wire v$_10494_out1;
wire v$_10627_out0;
wire v$_10627_out1;
wire v$_10628_out0;
wire v$_10628_out1;
wire v$_11057_out0;
wire v$_11057_out1;
wire v$_11058_out0;
wire v$_11058_out1;
wire v$_1108_out0;
wire v$_1109_out0;
wire v$_11302_out0;
wire v$_11302_out1;
wire v$_11303_out0;
wire v$_11303_out1;
wire v$_11630_out0;
wire v$_11630_out1;
wire v$_11631_out0;
wire v$_11631_out1;
wire v$_12039_out0;
wire v$_12039_out1;
wire v$_12040_out0;
wire v$_12040_out1;
wire v$_12741_out0;
wire v$_12741_out1;
wire v$_12742_out0;
wire v$_12742_out1;
wire v$_12787_out0;
wire v$_12788_out0;
wire v$_13007_out0;
wire v$_13008_out0;
wire v$_1375_out0;
wire v$_1376_out0;
wire v$_1554_out0;
wire v$_1555_out0;
wire v$_1743_out0;
wire v$_1744_out0;
wire v$_1864_out0;
wire v$_1864_out1;
wire v$_1865_out0;
wire v$_1865_out1;
wire v$_1868_out0;
wire v$_1868_out1;
wire v$_1869_out0;
wire v$_1869_out1;
wire v$_2193_out0;
wire v$_2193_out1;
wire v$_2194_out0;
wire v$_2194_out1;
wire v$_2400_out0;
wire v$_2400_out1;
wire v$_2401_out0;
wire v$_2401_out1;
wire v$_2495_out0;
wire v$_2495_out1;
wire v$_2496_out0;
wire v$_2496_out1;
wire v$_266_out0;
wire v$_266_out1;
wire v$_267_out0;
wire v$_267_out1;
wire v$_2714_out0;
wire v$_2714_out1;
wire v$_2715_out0;
wire v$_2715_out1;
wire v$_2732_out0;
wire v$_2732_out1;
wire v$_2733_out0;
wire v$_2733_out1;
wire v$_2736_out0;
wire v$_2736_out1;
wire v$_2737_out0;
wire v$_2737_out1;
wire v$_3183_out0;
wire v$_3183_out1;
wire v$_3184_out0;
wire v$_3184_out1;
wire v$_3284_out0;
wire v$_3284_out1;
wire v$_3285_out0;
wire v$_3285_out1;
wire v$_3288_out1;
wire v$_3289_out1;
wire v$_3433_out0;
wire v$_3433_out1;
wire v$_3434_out0;
wire v$_3434_out1;
wire v$_3451_out0;
wire v$_3451_out1;
wire v$_3452_out0;
wire v$_3452_out1;
wire v$_3651_out0;
wire v$_3651_out1;
wire v$_3652_out0;
wire v$_3652_out1;
wire v$_3805_out0;
wire v$_3805_out1;
wire v$_3806_out0;
wire v$_3806_out1;
wire v$_38_out0;
wire v$_398_out0;
wire v$_399_out0;
wire v$_39_out0;
wire v$_4077_out0;
wire v$_4078_out0;
wire v$_4743_out0;
wire v$_4743_out1;
wire v$_4744_out0;
wire v$_4744_out1;
wire v$_4849_out0;
wire v$_4849_out1;
wire v$_4850_out0;
wire v$_4850_out1;
wire v$_485_out0;
wire v$_486_out0;
wire v$_4885_out0;
wire v$_4885_out1;
wire v$_4886_out0;
wire v$_4886_out1;
wire v$_4887_out0;
wire v$_4888_out0;
wire v$_4988_out0;
wire v$_4988_out1;
wire v$_4989_out0;
wire v$_4989_out1;
wire v$_5052_out0;
wire v$_5053_out0;
wire v$_5187_out0;
wire v$_5187_out1;
wire v$_5188_out0;
wire v$_5188_out1;
wire v$_5189_out0;
wire v$_5189_out1;
wire v$_5190_out0;
wire v$_5190_out1;
wire v$_5191_out0;
wire v$_5191_out1;
wire v$_5192_out0;
wire v$_5192_out1;
wire v$_5193_out0;
wire v$_5193_out1;
wire v$_5194_out0;
wire v$_5194_out1;
wire v$_5195_out0;
wire v$_5195_out1;
wire v$_5196_out0;
wire v$_5196_out1;
wire v$_5197_out0;
wire v$_5197_out1;
wire v$_5198_out0;
wire v$_5198_out1;
wire v$_5488_out0;
wire v$_5488_out1;
wire v$_5489_out0;
wire v$_5489_out1;
wire v$_5597_out0;
wire v$_5597_out1;
wire v$_5598_out0;
wire v$_5598_out1;
wire v$_5720_out0;
wire v$_5721_out0;
wire v$_6015_out0;
wire v$_6016_out0;
wire v$_6017_out0;
wire v$_6017_out1;
wire v$_6018_out0;
wire v$_6018_out1;
wire v$_6057_out0;
wire v$_6057_out1;
wire v$_6058_out0;
wire v$_6058_out1;
wire v$_6308_out0;
wire v$_6308_out1;
wire v$_6309_out0;
wire v$_6309_out1;
wire v$_6349_out0;
wire v$_6349_out1;
wire v$_6350_out0;
wire v$_6350_out1;
wire v$_6383_out0;
wire v$_6383_out1;
wire v$_6384_out0;
wire v$_6384_out1;
wire v$_6473_out0;
wire v$_6473_out1;
wire v$_6474_out0;
wire v$_6474_out1;
wire v$_6546_out0;
wire v$_6547_out0;
wire v$_6815_out0;
wire v$_6815_out1;
wire v$_6816_out0;
wire v$_6816_out1;
wire v$_6843_out0;
wire v$_6844_out0;
wire v$_6962_out0;
wire v$_6963_out0;
wire v$_7094_out0;
wire v$_7095_out0;
wire v$_7294_out0;
wire v$_7294_out1;
wire v$_7295_out0;
wire v$_7295_out1;
wire v$_7432_out0;
wire v$_7433_out0;
wire v$_7576_out0;
wire v$_7577_out0;
wire v$_7653_out0;
wire v$_7653_out1;
wire v$_7654_out0;
wire v$_7654_out1;
wire v$_7655_out0;
wire v$_7655_out1;
wire v$_7656_out0;
wire v$_7656_out1;
wire v$_7657_out0;
wire v$_7657_out1;
wire v$_7658_out0;
wire v$_7658_out1;
wire v$_7659_out0;
wire v$_7659_out1;
wire v$_765_out0;
wire v$_7660_out0;
wire v$_7660_out1;
wire v$_7661_out0;
wire v$_7661_out1;
wire v$_7662_out0;
wire v$_7662_out1;
wire v$_7663_out0;
wire v$_7663_out1;
wire v$_7664_out0;
wire v$_7664_out1;
wire v$_766_out0;
wire v$_7862_out0;
wire v$_7862_out1;
wire v$_7863_out0;
wire v$_7863_out1;
wire v$_7866_out0;
wire v$_7866_out1;
wire v$_7867_out0;
wire v$_7867_out1;
wire v$_837_out0;
wire v$_837_out1;
wire v$_838_out0;
wire v$_838_out1;
wire v$_839_out0;
wire v$_839_out1;
wire v$_840_out0;
wire v$_840_out1;
wire v$_8418_out0;
wire v$_8419_out0;
wire v$_841_out0;
wire v$_841_out1;
wire v$_8426_out0;
wire v$_8427_out0;
wire v$_842_out0;
wire v$_842_out1;
wire v$_843_out0;
wire v$_843_out1;
wire v$_844_out0;
wire v$_844_out1;
wire v$_845_out0;
wire v$_845_out1;
wire v$_846_out0;
wire v$_846_out1;
wire v$_847_out0;
wire v$_847_out1;
wire v$_848_out0;
wire v$_848_out1;
wire v$_8852_out0;
wire v$_8855_out0;
wire v$_8872_out0;
wire v$_8873_out0;
wire v$_9112_out0;
wire v$_9113_out0;
wire v$_9237_out0;
wire v$_9238_out0;
wire v$_9360_out0;
wire v$_9360_out1;
wire v$_9361_out0;
wire v$_9361_out1;
wire v$_9470_out0;
wire v$_9470_out1;
wire v$_9471_out0;
wire v$_9471_out1;
wire v$_9644_out0;
wire v$_9644_out1;
wire v$_9645_out0;
wire v$_9645_out1;
wire v$_9711_out0;
wire v$_9712_out0;
wire v$_9897_out0;
wire v$_9897_out1;
wire v$_9898_out0;
wire v$_9898_out1;
wire v$_9899_out0;
wire v$_9899_out1;
wire v$_9900_out0;
wire v$_9900_out1;
wire v$_9901_out0;
wire v$_9901_out1;
wire v$_9902_out0;
wire v$_9902_out1;
wire v$_9903_out0;
wire v$_9903_out1;
wire v$_9904_out0;
wire v$_9904_out1;
wire v$_9905_out0;
wire v$_9905_out1;
wire v$_9906_out0;
wire v$_9906_out1;
wire v$_9907_out0;
wire v$_9907_out1;
wire v$_9908_out0;
wire v$_9908_out1;
wire v$_9909_out0;
wire v$_9909_out1;
wire v$_9910_out0;
wire v$_9910_out1;
wire v$increment_12632_out0;
wire v$increment_12633_out0;

always @(posedge clk) v$FF1_2_out0 <= v$NEWINTERRUPT_4784_out0;
always @(posedge clk) v$FF1_3_out0 <= v$NEWINTERRUPT_4785_out0;
always @(posedge clk) v$FF1_178_out0 <= v$G3_5549_out0;
always @(posedge clk) v$FF1_179_out0 <= v$G3_5550_out0;
always @(posedge clk) v$INT2_221_out0 <= v$I2EN_10989_out0 ? v$SEL1_7748_out0 : v$INT2_221_out0;
always @(posedge clk) v$INT2_222_out0 <= v$I2EN_10990_out0 ? v$SEL1_7749_out0 : v$INT2_222_out0;
always @(posedge clk) v$FF3_227_out0 <= v$ShiftEN_5265_out0 ? v$MUX3_12536_out0 : v$FF3_227_out0;
always @(posedge clk) v$FF3_228_out0 <= v$ShiftEN_5266_out0 ? v$MUX3_12537_out0 : v$FF3_228_out0;
always @(posedge clk) v$INT3_233_out0 <= v$I3EN_12565_out0 ? v$SEL1_7748_out0 : v$INT3_233_out0;
always @(posedge clk) v$INT3_234_out0 <= v$I3EN_12566_out0 ? v$SEL1_7749_out0 : v$INT3_234_out0;
always @(posedge clk) v$REG13_248_out0 <= v$HALT0_290_out0;
always @(posedge clk) v$FF0_374_out0 <= v$CLK4_7986_out0 ? v$G1_10609_out0 : v$FF0_374_out0;
always @(posedge clk) v$FF0_375_out0 <= v$CLK4_7987_out0 ? v$G1_10610_out0 : v$FF0_375_out0;
always @(posedge clk) v$REG2_376_out0 <= v$increment_12632_out0 ? v$A2_10173_out0 : v$REG2_376_out0;
always @(posedge clk) v$REG2_377_out0 <= v$increment_12633_out0 ? v$A2_10174_out0 : v$REG2_377_out0;
always @(posedge clk) v$REG1_457_out0 <= v$G14_11038_out0 ? v$A_7280_out0 : v$REG1_457_out0;
always @(posedge clk) v$REG1_458_out0 <= v$G14_11039_out0 ? v$A_7281_out0 : v$REG1_458_out0;
always @(posedge clk) v$FF1_467_out0 <= v$CLK4_7986_out0 ? v$G21_12498_out0 : v$FF1_467_out0;
always @(posedge clk) v$FF1_468_out0 <= v$CLK4_7987_out0 ? v$G21_12499_out0 : v$FF1_468_out0;
always @(posedge clk) v$FF2_469_out0 <= v$LDMAIN_9330_out0;
always @(posedge clk) v$FF2_470_out0 <= v$LDMAIN_9331_out0;
always @(posedge clk) v$FF3_532_out0 <= v$Shift_6566_out0 ? v$FF1_11343_out0 : v$FF3_532_out0;
always @(posedge clk) v$FF3_533_out0 <= v$Shift_6567_out0 ? v$FF1_11344_out0 : v$FF3_533_out0;
always @(posedge clk) v$FF1_601_out0 <= v$NEWINTERRUPT_3080_out0;
always @(posedge clk) v$FF1_602_out0 <= v$NEWINTERRUPT_3081_out0;
always @(posedge clk) v$FF2_779_out0 <= v$Shift_6566_out0 ? v$FF7_9941_out0 : v$FF2_779_out0;
always @(posedge clk) v$FF2_780_out0 <= v$Shift_6567_out0 ? v$FF7_9942_out0 : v$FF2_780_out0;
always @(posedge clk) v$FF5_933_out0 <= v$SHIFTEN_6401_out0 ? v$MUX1_1489_out0 : v$FF5_933_out0;
always @(posedge clk) v$FF5_934_out0 <= v$SHIFTEN_6402_out0 ? v$MUX1_1490_out0 : v$FF5_934_out0;
always @(posedge clk) v$FF5_935_out0 <= v$SHIFTEN_6403_out0 ? v$MUX1_1491_out0 : v$FF5_935_out0;
always @(posedge clk) v$FF5_936_out0 <= v$SHIFTEN_6404_out0 ? v$MUX1_1492_out0 : v$FF5_936_out0;
always @(posedge clk) v$FF5_937_out0 <= v$SHIFTEN_6405_out0 ? v$MUX1_1493_out0 : v$FF5_937_out0;
always @(posedge clk) v$FF5_938_out0 <= v$SHIFTEN_6406_out0 ? v$MUX1_1494_out0 : v$FF5_938_out0;
always @(posedge clk) v$FF5_939_out0 <= v$SHIFTEN_6407_out0 ? v$MUX1_1495_out0 : v$FF5_939_out0;
always @(posedge clk) v$FF5_940_out0 <= v$SHIFTEN_6408_out0 ? v$MUX1_1496_out0 : v$FF5_940_out0;
always @(posedge clk) v$FF5_941_out0 <= v$SHIFTEN_6409_out0 ? v$MUX1_1497_out0 : v$FF5_941_out0;
always @(posedge clk) v$FF5_942_out0 <= v$SHIFTEN_6410_out0 ? v$MUX1_1498_out0 : v$FF5_942_out0;
always @(posedge clk) v$FF5_943_out0 <= v$SHIFTEN_6411_out0 ? v$MUX1_1499_out0 : v$FF5_943_out0;
always @(posedge clk) v$FF5_944_out0 <= v$SHIFTEN_6412_out0 ? v$MUX1_1500_out0 : v$FF5_944_out0;
always @(posedge clk) v$FF4_1281_out0 <= v$ShiftEN_5265_out0 ? v$MUX4_10904_out0 : v$FF4_1281_out0;
always @(posedge clk) v$FF4_1282_out0 <= v$ShiftEN_5266_out0 ? v$MUX4_10905_out0 : v$FF4_1282_out0;
always @(posedge clk) v$FF11_1377_out0 <= v$G50_11471_out0;
always @(posedge clk) v$FF11_1378_out0 <= v$G50_11472_out0;
always @(posedge clk) v$FF1_1433_out0 <= v$G4_10044_out0;
always @(posedge clk) v$FF1_1434_out0 <= v$G4_10045_out0;
always @(posedge clk) v$FF6_1523_out0 <= v$SHIFTEN_6401_out0 ? v$MUX3_6670_out0 : v$FF6_1523_out0;
always @(posedge clk) v$FF6_1524_out0 <= v$SHIFTEN_6402_out0 ? v$MUX3_6671_out0 : v$FF6_1524_out0;
always @(posedge clk) v$FF6_1525_out0 <= v$SHIFTEN_6403_out0 ? v$MUX3_6672_out0 : v$FF6_1525_out0;
always @(posedge clk) v$FF6_1526_out0 <= v$SHIFTEN_6404_out0 ? v$MUX3_6673_out0 : v$FF6_1526_out0;
always @(posedge clk) v$FF6_1527_out0 <= v$SHIFTEN_6405_out0 ? v$MUX3_6674_out0 : v$FF6_1527_out0;
always @(posedge clk) v$FF6_1528_out0 <= v$SHIFTEN_6406_out0 ? v$MUX3_6675_out0 : v$FF6_1528_out0;
always @(posedge clk) v$FF6_1529_out0 <= v$SHIFTEN_6407_out0 ? v$MUX3_6676_out0 : v$FF6_1529_out0;
always @(posedge clk) v$FF6_1530_out0 <= v$SHIFTEN_6408_out0 ? v$MUX3_6677_out0 : v$FF6_1530_out0;
always @(posedge clk) v$FF6_1531_out0 <= v$SHIFTEN_6409_out0 ? v$MUX3_6678_out0 : v$FF6_1531_out0;
always @(posedge clk) v$FF6_1532_out0 <= v$SHIFTEN_6410_out0 ? v$MUX3_6679_out0 : v$FF6_1532_out0;
always @(posedge clk) v$FF6_1533_out0 <= v$SHIFTEN_6411_out0 ? v$MUX3_6680_out0 : v$FF6_1533_out0;
always @(posedge clk) v$FF6_1534_out0 <= v$SHIFTEN_6412_out0 ? v$MUX3_6681_out0 : v$FF6_1534_out0;
always @(posedge clk) v$REG3_1589_out0 <= v$G55_12935_out0 ? v$MUX5_7734_out0 : v$REG3_1589_out0;
always @(posedge clk) v$REG3_1590_out0 <= v$G55_12936_out0 ? v$MUX5_7735_out0 : v$REG3_1590_out0;
always @(posedge clk) v$FF2_1717_out0 <= v$ShiftEN_5265_out0 ? v$MUX2_8870_out0 : v$FF2_1717_out0;
always @(posedge clk) v$FF2_1718_out0 <= v$ShiftEN_5266_out0 ? v$MUX2_8871_out0 : v$FF2_1718_out0;
always @(posedge clk) v$REG12_2023_out0 <= v$HALT1_2849_out0 ? v$RAMADDR1_8300_out0 : v$REG12_2023_out0;
always @(posedge clk) v$FF3_2072_out0 <= v$G53_12287_out0;
always @(posedge clk) v$FF4_2489_out0 <= v$CAPTURE_207_out0 ? v$G6_7901_out0 : v$FF4_2489_out0;
always @(posedge clk) v$FF4_2490_out0 <= v$CAPTURE_208_out0 ? v$G6_7902_out0 : v$FF4_2490_out0;
always @(posedge clk) v$REG1_2760_out0 <= v$EN_11112_out0 ? v$MODE_7108_out0 : v$REG1_2760_out0;
always @(posedge clk) v$REG1_2761_out0 <= v$EN_11113_out0 ? v$MODE_7109_out0 : v$REG1_2761_out0;
always @(posedge clk) v$REG8_2804_out0 <= v$SELIN_12946_out0;
always @(posedge clk) v$FF0_2992_out0 <= v$CLK4_12743_out0 ? v$MUX1_5175_out0 : v$FF0_2992_out0;
always @(posedge clk) v$FF0_2993_out0 <= v$CLK4_12744_out0 ? v$MUX1_5176_out0 : v$FF0_2993_out0;
always @(posedge clk) v$FF2_3000_out0 <= v$CLK4_12743_out0 ? v$MUX3_4145_out0 : v$FF2_3000_out0;
always @(posedge clk) v$FF2_3001_out0 <= v$CLK4_12744_out0 ? v$MUX3_4146_out0 : v$FF2_3001_out0;
always @(posedge clk) v$FF5_3159_out0 <= v$EQ2_7440_out0;
always @(posedge clk) v$FF5_3160_out0 <= v$EQ2_7441_out0;
always @(posedge clk) v$REG1_3286_out0 <= v$D1_9486_out1 ? v$DIN3_9801_out0 : v$REG1_3286_out0;
always @(posedge clk) v$REG1_3287_out0 <= v$D1_9487_out1 ? v$DIN3_9802_out0 : v$REG1_3287_out0;
always @(posedge clk) v$FF0_3399_out0 <= v$G1_8760_out0;
always @(posedge clk) v$FF0_3400_out0 <= v$G1_8761_out0;
always @(posedge clk) v$REG2_3503_out0 <= v$HALT_11481_out0 ? v$G8_10979_out0 : v$REG2_3503_out0;
always @(posedge clk) v$FF1_3605_out0 <= v$NEXTSTATE_9107_out0;
always @(posedge clk) v$FF1_3606_out0 <= v$NEXTSTATE_9108_out0;
always @(posedge clk) v$FF1_3695_out0 <= v$G45_10651_out0;
always @(posedge clk) v$REG14_3705_out0 <= v$HALT1_2849_out0;
always @(posedge clk) v$FF1_4029_out0 <= v$INTERRUPT0_7520_out0;
always @(posedge clk) v$FF1_4030_out0 <= v$INTERRUPT0_7521_out0;
always @(posedge clk) v$FF1_4163_out0 <= v$CAPTURE_207_out0 ? v$I3_3228_out0 : v$FF1_4163_out0;
always @(posedge clk) v$FF1_4164_out0 <= v$CAPTURE_208_out0 ? v$I3_3229_out0 : v$FF1_4164_out0;
always @(posedge clk) v$REG7_4199_out0 <= v$G84_504_out0;
always @(posedge clk) v$REG4_4650_out0 <= v$G66_5924_out0 ? v$MUX1_10579_out0 : v$REG4_4650_out0;
always @(posedge clk) v$REG4_4651_out0 <= v$G66_5925_out0 ? v$MUX1_10580_out0 : v$REG4_4651_out0;
always @(posedge clk) v$REG3_4759_out0 <= v$EXEC1_13169_out0 ? v$_809_out0 : v$REG3_4759_out0;
always @(posedge clk) v$REG3_4760_out0 <= v$EXEC1_13170_out0 ? v$_810_out0 : v$REG3_4760_out0;
always @(posedge clk) v$FF4_4776_out0 <= v$EQ1_9709_out0;
always @(posedge clk) v$FF4_4777_out0 <= v$EQ1_9710_out0;
always @(posedge clk) v$REG1_4808_out0 <= v$HALTVALID_5289_out0 ? v$NEXTSTATE_9109_out0 : v$REG1_4808_out0;
always @(posedge clk) v$FF3_4929_out0 <= v$RX_40_out0;
always @(posedge clk) v$FF3_4930_out0 <= v$RX_41_out0;
always @(posedge clk) v$FF3_5109_out0 <= v$CAPTURE_207_out0 ? v$G9_10813_out0 : v$FF3_5109_out0;
always @(posedge clk) v$FF3_5110_out0 <= v$CAPTURE_208_out0 ? v$G9_10814_out0 : v$FF3_5110_out0;
always @(posedge clk) v$FF10_5406_out0 <= v$HALT_8544_out0;
always @(posedge clk) v$FF10_5407_out0 <= v$HALT_8545_out0;
always @(posedge clk) v$FF8_5529_out0 <= v$ShiftEN_5265_out0 ? v$MUX8_725_out0 : v$FF8_5529_out0;
always @(posedge clk) v$FF8_5530_out0 <= v$ShiftEN_5266_out0 ? v$MUX8_726_out0 : v$FF8_5530_out0;
always @(posedge clk) v$FF4_5562_out0 <= v$G68_10489_out0;
always @(posedge clk) v$FF4_5563_out0 <= v$G68_10490_out0;
always @(posedge clk) v$FF7_5594_out0 <= v$G62_7570_out0 ? v$R_6019_out0 : v$FF7_5594_out0;
always @(posedge clk) v$FF7_5595_out0 <= v$G62_7571_out0 ? v$R_6020_out0 : v$FF7_5595_out0;
always @(posedge clk) v$FF1_5716_out0 <= v$EXEC2_5557_out0 ? v$S_12723_out0 : v$FF1_5716_out0;
always @(posedge clk) v$FF1_5717_out0 <= v$EXEC2_5558_out0 ? v$S_12724_out0 : v$FF1_5717_out0;
always @(posedge clk) v$FF4_5735_out0 <= v$Shift_6566_out0 ? v$RX_1727_out0 : v$FF4_5735_out0;
always @(posedge clk) v$FF4_5736_out0 <= v$Shift_6567_out0 ? v$RX_1728_out0 : v$FF4_5736_out0;
always @(posedge clk) v$FF7_5772_out0 <= v$SHIFTEN_6401_out0 ? v$MUX8_2316_out0 : v$FF7_5772_out0;
always @(posedge clk) v$FF7_5773_out0 <= v$SHIFTEN_6402_out0 ? v$MUX8_2317_out0 : v$FF7_5773_out0;
always @(posedge clk) v$FF7_5774_out0 <= v$SHIFTEN_6403_out0 ? v$MUX8_2318_out0 : v$FF7_5774_out0;
always @(posedge clk) v$FF7_5775_out0 <= v$SHIFTEN_6404_out0 ? v$MUX8_2319_out0 : v$FF7_5775_out0;
always @(posedge clk) v$FF7_5776_out0 <= v$SHIFTEN_6405_out0 ? v$MUX8_2320_out0 : v$FF7_5776_out0;
always @(posedge clk) v$FF7_5777_out0 <= v$SHIFTEN_6406_out0 ? v$MUX8_2321_out0 : v$FF7_5777_out0;
always @(posedge clk) v$FF7_5778_out0 <= v$SHIFTEN_6407_out0 ? v$MUX8_2322_out0 : v$FF7_5778_out0;
always @(posedge clk) v$FF7_5779_out0 <= v$SHIFTEN_6408_out0 ? v$MUX8_2323_out0 : v$FF7_5779_out0;
always @(posedge clk) v$FF7_5780_out0 <= v$SHIFTEN_6409_out0 ? v$MUX8_2324_out0 : v$FF7_5780_out0;
always @(posedge clk) v$FF7_5781_out0 <= v$SHIFTEN_6410_out0 ? v$MUX8_2325_out0 : v$FF7_5781_out0;
always @(posedge clk) v$FF7_5782_out0 <= v$SHIFTEN_6411_out0 ? v$MUX8_2326_out0 : v$FF7_5782_out0;
always @(posedge clk) v$FF7_5783_out0 <= v$SHIFTEN_6412_out0 ? v$MUX8_2327_out0 : v$FF7_5783_out0;
always @(posedge clk) v$REG1_6069_out0 <= v$G6_2205_out0;
always @(posedge clk) v$REG1_6141_out0 <= v$EXEC2_6435_out0 ? v$MUX5_9877_out0 : v$REG1_6141_out0;
always @(posedge clk) v$REG1_6142_out0 <= v$EXEC2_6436_out0 ? v$MUX5_9878_out0 : v$REG1_6142_out0;
always @(posedge clk) v$FF6_6215_out0 <= v$Shift_6566_out0 ? v$FF8_11778_out0 : v$FF6_6215_out0;
always @(posedge clk) v$FF6_6216_out0 <= v$Shift_6567_out0 ? v$FF8_11779_out0 : v$FF6_6216_out0;
always @(posedge clk) v$FF0_6397_out0 <= v$G12_1148_out0;
always @(posedge clk) v$FF0_6398_out0 <= v$G12_1149_out0;
always @(posedge clk) v$FF2_6413_out0 <= v$STATUSREAD_835_out0;
always @(posedge clk) v$FF2_6414_out0 <= v$STATUSREAD_836_out0;
always @(posedge clk) v$FF1_6417_out0 <= v$ShiftEN_5265_out0 ? v$MUX1_345_out0 : v$FF1_6417_out0;
always @(posedge clk) v$FF1_6418_out0 <= v$ShiftEN_5266_out0 ? v$MUX1_346_out0 : v$FF1_6418_out0;
always @(posedge clk) v$FF1_6568_out0 <= v$CLK4_12743_out0 ? v$MUX2_4675_out0 : v$FF1_6568_out0;
always @(posedge clk) v$FF1_6569_out0 <= v$CLK4_12744_out0 ? v$MUX2_4676_out0 : v$FF1_6569_out0;
always @(posedge clk) v$REG11_6578_out0 <= v$HALT1_2849_out0 ? v$DATAIN1_6590_out0 : v$REG11_6578_out0;
always @(posedge clk) v$FF1_6586_out0 <= v$G2_3619_out0;
always @(posedge clk) v$FF1_6587_out0 <= v$G2_3620_out0;
always @(posedge clk) v$FF3_6686_out0 <= v$SHIFTEN_6401_out0 ? v$MUX5_6500_out0 : v$FF3_6686_out0;
always @(posedge clk) v$FF3_6687_out0 <= v$SHIFTEN_6402_out0 ? v$MUX5_6501_out0 : v$FF3_6687_out0;
always @(posedge clk) v$FF3_6688_out0 <= v$SHIFTEN_6403_out0 ? v$MUX5_6502_out0 : v$FF3_6688_out0;
always @(posedge clk) v$FF3_6689_out0 <= v$SHIFTEN_6404_out0 ? v$MUX5_6503_out0 : v$FF3_6689_out0;
always @(posedge clk) v$FF3_6690_out0 <= v$SHIFTEN_6405_out0 ? v$MUX5_6504_out0 : v$FF3_6690_out0;
always @(posedge clk) v$FF3_6691_out0 <= v$SHIFTEN_6406_out0 ? v$MUX5_6505_out0 : v$FF3_6691_out0;
always @(posedge clk) v$FF3_6692_out0 <= v$SHIFTEN_6407_out0 ? v$MUX5_6506_out0 : v$FF3_6692_out0;
always @(posedge clk) v$FF3_6693_out0 <= v$SHIFTEN_6408_out0 ? v$MUX5_6507_out0 : v$FF3_6693_out0;
always @(posedge clk) v$FF3_6694_out0 <= v$SHIFTEN_6409_out0 ? v$MUX5_6508_out0 : v$FF3_6694_out0;
always @(posedge clk) v$FF3_6695_out0 <= v$SHIFTEN_6410_out0 ? v$MUX5_6509_out0 : v$FF3_6695_out0;
always @(posedge clk) v$FF3_6696_out0 <= v$SHIFTEN_6411_out0 ? v$MUX5_6510_out0 : v$FF3_6696_out0;
always @(posedge clk) v$FF3_6697_out0 <= v$SHIFTEN_6412_out0 ? v$MUX5_6511_out0 : v$FF3_6697_out0;
always @(posedge clk) v$REG1_6863_out0 <= v$EXEC2_5557_out0 ? v$MUX6_9251_out0 : v$REG1_6863_out0;
always @(posedge clk) v$REG1_6864_out0 <= v$EXEC2_5558_out0 ? v$MUX6_9252_out0 : v$REG1_6864_out0;
always @(posedge clk) v$FF1_6867_out0 <= v$G5_5122_out0 ? v$A1_6425_out1 : v$FF1_6867_out0;
always @(posedge clk) v$FF1_6868_out0 <= v$G5_5123_out0 ? v$A1_6426_out1 : v$FF1_6868_out0;
always @(posedge clk) v$FF8_6889_out0 <= v$EQ3_2888_out0;
always @(posedge clk) v$FF8_6890_out0 <= v$EQ3_2889_out0;
always @(posedge clk) v$FF9_6996_out0 <= v$STP$DECODED_11614_out0;
always @(posedge clk) v$FF9_6997_out0 <= v$STP$DECODED_11615_out0;
always @(posedge clk) v$S$FF_7118_out0 <= v$EXEC2_461_out0 ? v$S_7016_out0 : v$S$FF_7118_out0;
always @(posedge clk) v$S$FF_7119_out0 <= v$EXEC2_462_out0 ? v$S_7017_out0 : v$S$FF_7119_out0;
always @(posedge clk) v$REG1_7183_out0 <= v$EXEC2_701_out0 ? v$MUX5_5450_out0 : v$REG1_7183_out0;
always @(posedge clk) v$REG1_7184_out0 <= v$EXEC2_702_out0 ? v$MUX5_5451_out0 : v$REG1_7184_out0;
always @(posedge clk) v$FF14_7185_out0 <= v$VALID_2425_out0;
always @(posedge clk) v$FF14_7186_out0 <= v$VALID_2426_out0;
always @(posedge clk) v$FF3_7189_out0 <= v$CLK4_12743_out0 ? v$MUX4_12118_out0 : v$FF3_7189_out0;
always @(posedge clk) v$FF3_7190_out0 <= v$CLK4_12744_out0 ? v$MUX4_12119_out0 : v$FF3_7190_out0;
always @(posedge clk) v$REG4_7248_out0 <= v$G88_4994_out0;
always @(posedge clk) v$REG3_7255_out0 <= v$D1_9486_out3 ? v$DIN3_9801_out0 : v$REG3_7255_out0;
always @(posedge clk) v$REG3_7256_out0 <= v$D1_9487_out3 ? v$DIN3_9802_out0 : v$REG3_7256_out0;
always @(posedge clk) v$FF1_7292_out0 <= v$G1_2894_out0;
always @(posedge clk) v$FF1_7293_out0 <= v$G1_2895_out0;
always @(posedge clk) v$REG3_7578_out0 <= v$G18_5076_out0 ? v$SEL4_6522_out0 : v$REG3_7578_out0;
always @(posedge clk) v$REG3_7579_out0 <= v$G18_5077_out0 ? v$SEL4_6523_out0 : v$REG3_7579_out0;
always @(posedge clk) v$REG2_7598_out0 <= v$IR2$VALID_8838_out0 ? v$_6015_out0 : v$REG2_7598_out0;
always @(posedge clk) v$REG2_7599_out0 <= v$IR2$VALID_8839_out0 ? v$_6016_out0 : v$REG2_7599_out0;
always @(posedge clk) v$FF15_8373_out0 <= v$HALT$PREV$PREV_12829_out0;
always @(posedge clk) v$FF15_8374_out0 <= v$HALT$PREV$PREV_12830_out0;
always @(posedge clk) v$FF7_8410_out0 <= v$STALL_12672_out0;
always @(posedge clk) v$FF7_8411_out0 <= v$STALL_12673_out0;
always @(posedge clk) v$PCNORMAL_8422_out0 <= v$G33_7075_out0 ? v$SUM_9219_out0 : v$PCNORMAL_8422_out0;
always @(posedge clk) v$PCNORMAL_8423_out0 <= v$G33_7076_out0 ? v$SUM_9220_out0 : v$PCNORMAL_8423_out0;
v$RAM1_8558 I8558 (v$RAM1_8558_out0, v$RAMADDR_9169_out0, v$MUX2_11061_out0, v$RAMWEN_12732_out0, clk);
always @(posedge clk) v$FF2_8662_out0 <= v$G7_9511_out0;
always @(posedge clk) v$FF2_8663_out0 <= v$G7_9512_out0;
always @(posedge clk) v$FF2_8664_out0 <= v$G7_9513_out0;
always @(posedge clk) v$FF2_8665_out0 <= v$G7_9514_out0;
always @(posedge clk) v$FF2_8666_out0 <= v$G7_9515_out0;
always @(posedge clk) v$FF2_8667_out0 <= v$G7_9516_out0;
always @(posedge clk) v$FF2_8668_out0 <= v$G4_7633_out0;
always @(posedge clk) v$FF2_8669_out0 <= v$G4_7634_out0;
always @(posedge clk) v$FF2_8670_out0 <= v$G4_7635_out0;
always @(posedge clk) v$FF2_8671_out0 <= v$G4_7636_out0;
always @(posedge clk) v$FF2_8672_out0 <= v$G4_7637_out0;
always @(posedge clk) v$FF2_8673_out0 <= v$G7_9517_out0;
always @(posedge clk) v$FF2_8674_out0 <= v$G7_9518_out0;
always @(posedge clk) v$FF2_8675_out0 <= v$G7_9519_out0;
always @(posedge clk) v$FF2_8676_out0 <= v$G7_9520_out0;
always @(posedge clk) v$FF2_8677_out0 <= v$G7_9521_out0;
always @(posedge clk) v$FF2_8678_out0 <= v$G7_9522_out0;
always @(posedge clk) v$FF2_8679_out0 <= v$G4_7638_out0;
always @(posedge clk) v$FF2_8680_out0 <= v$G4_7639_out0;
always @(posedge clk) v$FF2_8681_out0 <= v$G4_7640_out0;
always @(posedge clk) v$FF2_8682_out0 <= v$G4_7641_out0;
always @(posedge clk) v$FF2_8683_out0 <= v$G4_7642_out0;
always @(posedge clk) v$FF1_8718_out0 <= v$G16_4405_out0 ? v$G7_1007_out0 : v$FF1_8718_out0;
always @(posedge clk) v$FF1_8719_out0 <= v$G16_4406_out0 ? v$G7_1008_out0 : v$FF1_8719_out0;
always @(posedge clk) v$FF2_9024_out0 <= v$G51_13389_out0;
always @(posedge clk) v$FF4_9118_out0 <= v$G54_8868_out0;
always @(posedge clk) v$REG1_9161_out0 <= v$MUX1_13028_out0;
always @(posedge clk) v$REG1_9162_out0 <= v$MUX1_13029_out0;
always @(posedge clk) v$FF1_9226_out0 <= v$EXEC2_6435_out0 ? v$S_6897_out0 : v$FF1_9226_out0;
always @(posedge clk) v$FF1_9227_out0 <= v$EXEC2_6436_out0 ? v$S_6898_out0 : v$FF1_9227_out0;
always @(posedge clk) v$REG1_9488_out0 <= v$IR1$VALID_58_out0 ? v$RM_12933_out0 : v$REG1_9488_out0;
always @(posedge clk) v$REG1_9489_out0 <= v$IR1$VALID_59_out0 ? v$RM_12934_out0 : v$REG1_9489_out0;
always @(posedge clk) v$FF10_9601_out0 <= v$WREN_7251_out0;
always @(posedge clk) v$FF10_9602_out0 <= v$WREN_7252_out0;
always @(posedge clk) v$FF8_9843_out0 <= v$SHIFTEN_6401_out0 ? v$MUX4_11896_out0 : v$FF8_9843_out0;
always @(posedge clk) v$FF8_9844_out0 <= v$SHIFTEN_6402_out0 ? v$MUX4_11897_out0 : v$FF8_9844_out0;
always @(posedge clk) v$FF8_9845_out0 <= v$SHIFTEN_6403_out0 ? v$MUX4_11898_out0 : v$FF8_9845_out0;
always @(posedge clk) v$FF8_9846_out0 <= v$SHIFTEN_6404_out0 ? v$MUX4_11899_out0 : v$FF8_9846_out0;
always @(posedge clk) v$FF8_9847_out0 <= v$SHIFTEN_6405_out0 ? v$MUX4_11900_out0 : v$FF8_9847_out0;
always @(posedge clk) v$FF8_9848_out0 <= v$SHIFTEN_6406_out0 ? v$MUX4_11901_out0 : v$FF8_9848_out0;
always @(posedge clk) v$FF8_9849_out0 <= v$SHIFTEN_6407_out0 ? v$MUX4_11902_out0 : v$FF8_9849_out0;
always @(posedge clk) v$FF8_9850_out0 <= v$SHIFTEN_6408_out0 ? v$MUX4_11903_out0 : v$FF8_9850_out0;
always @(posedge clk) v$FF8_9851_out0 <= v$SHIFTEN_6409_out0 ? v$MUX4_11904_out0 : v$FF8_9851_out0;
always @(posedge clk) v$FF8_9852_out0 <= v$SHIFTEN_6410_out0 ? v$MUX4_11905_out0 : v$FF8_9852_out0;
always @(posedge clk) v$FF8_9853_out0 <= v$SHIFTEN_6411_out0 ? v$MUX4_11906_out0 : v$FF8_9853_out0;
always @(posedge clk) v$FF8_9854_out0 <= v$SHIFTEN_6412_out0 ? v$MUX4_11907_out0 : v$FF8_9854_out0;
always @(posedge clk) v$FF7_9941_out0 <= v$Shift_6566_out0 ? v$FF6_6215_out0 : v$FF7_9941_out0;
always @(posedge clk) v$FF7_9942_out0 <= v$Shift_6567_out0 ? v$FF6_6216_out0 : v$FF7_9942_out0;
always @(posedge clk) v$FF2_9998_out0 <= v$CLK4_7986_out0 ? v$G24_6574_out0 : v$FF2_9998_out0;
always @(posedge clk) v$FF2_9999_out0 <= v$CLK4_7987_out0 ? v$G24_6575_out0 : v$FF2_9999_out0;
always @(posedge clk) v$FF2_10133_out0 <= v$SHIFTEN_6401_out0 ? v$MUX6_6937_out0 : v$FF2_10133_out0;
always @(posedge clk) v$FF2_10134_out0 <= v$SHIFTEN_6402_out0 ? v$MUX6_6938_out0 : v$FF2_10134_out0;
always @(posedge clk) v$FF2_10135_out0 <= v$SHIFTEN_6403_out0 ? v$MUX6_6939_out0 : v$FF2_10135_out0;
always @(posedge clk) v$FF2_10136_out0 <= v$SHIFTEN_6404_out0 ? v$MUX6_6940_out0 : v$FF2_10136_out0;
always @(posedge clk) v$FF2_10137_out0 <= v$SHIFTEN_6405_out0 ? v$MUX6_6941_out0 : v$FF2_10137_out0;
always @(posedge clk) v$FF2_10138_out0 <= v$SHIFTEN_6406_out0 ? v$MUX6_6942_out0 : v$FF2_10138_out0;
always @(posedge clk) v$FF2_10139_out0 <= v$SHIFTEN_6407_out0 ? v$MUX6_6943_out0 : v$FF2_10139_out0;
always @(posedge clk) v$FF2_10140_out0 <= v$SHIFTEN_6408_out0 ? v$MUX6_6944_out0 : v$FF2_10140_out0;
always @(posedge clk) v$FF2_10141_out0 <= v$SHIFTEN_6409_out0 ? v$MUX6_6945_out0 : v$FF2_10141_out0;
always @(posedge clk) v$FF2_10142_out0 <= v$SHIFTEN_6410_out0 ? v$MUX6_6946_out0 : v$FF2_10142_out0;
always @(posedge clk) v$FF2_10143_out0 <= v$SHIFTEN_6411_out0 ? v$MUX6_6947_out0 : v$FF2_10143_out0;
always @(posedge clk) v$FF2_10144_out0 <= v$SHIFTEN_6412_out0 ? v$MUX6_6948_out0 : v$FF2_10144_out0;
always @(posedge clk) v$REG1_10179_out0 <= v$MUX1_6647_out0;
always @(posedge clk) v$REG1_10180_out0 <= v$MUX1_6648_out0;
always @(posedge clk) v$REG2_10321_out0 <= v$R_13054_out0;
always @(posedge clk) v$REG2_10322_out0 <= v$R_13055_out0;
always @(posedge clk) v$FF3_10341_out0 <= v$INTERRUPT2_857_out0;
always @(posedge clk) v$FF3_10342_out0 <= v$INTERRUPT2_858_out0;
always @(posedge clk) v$FF6_10631_out0 <= v$ShiftEN_5265_out0 ? v$MUX6_6364_out0 : v$FF6_10631_out0;
always @(posedge clk) v$FF6_10632_out0 <= v$ShiftEN_5266_out0 ? v$MUX6_6365_out0 : v$FF6_10632_out0;
always @(posedge clk) v$FF2_10772_out0 <= v$G1_3667_out0;
always @(posedge clk) v$FF2_10773_out0 <= v$G1_3668_out0;
always @(posedge clk) v$REG2_10886_out0 <= v$G13_5410_out0 ? v$B_2056_out0 : v$REG2_10886_out0;
always @(posedge clk) v$REG2_10887_out0 <= v$G13_5411_out0 ? v$B_2057_out0 : v$REG2_10887_out0;
always @(posedge clk) v$INT0_11100_out0 <= v$I0EN_5551_out0 ? v$SEL1_7748_out0 : v$INT0_11100_out0;
always @(posedge clk) v$INT0_11101_out0 <= v$I0EN_5552_out0 ? v$SEL1_7749_out0 : v$INT0_11101_out0;
always @(posedge clk) v$FF3_11154_out0 <= v$CLK4_7986_out0 ? v$G32_11448_out0 : v$FF3_11154_out0;
always @(posedge clk) v$FF3_11155_out0 <= v$CLK4_7987_out0 ? v$G32_11449_out0 : v$FF3_11155_out0;
always @(posedge clk) v$FF4_11162_out0 <= v$SHIFTEN_6401_out0 ? v$MUX2_9342_out0 : v$FF4_11162_out0;
always @(posedge clk) v$FF4_11163_out0 <= v$SHIFTEN_6402_out0 ? v$MUX2_9343_out0 : v$FF4_11163_out0;
always @(posedge clk) v$FF4_11164_out0 <= v$SHIFTEN_6403_out0 ? v$MUX2_9344_out0 : v$FF4_11164_out0;
always @(posedge clk) v$FF4_11165_out0 <= v$SHIFTEN_6404_out0 ? v$MUX2_9345_out0 : v$FF4_11165_out0;
always @(posedge clk) v$FF4_11166_out0 <= v$SHIFTEN_6405_out0 ? v$MUX2_9346_out0 : v$FF4_11166_out0;
always @(posedge clk) v$FF4_11167_out0 <= v$SHIFTEN_6406_out0 ? v$MUX2_9347_out0 : v$FF4_11167_out0;
always @(posedge clk) v$FF4_11168_out0 <= v$SHIFTEN_6407_out0 ? v$MUX2_9348_out0 : v$FF4_11168_out0;
always @(posedge clk) v$FF4_11169_out0 <= v$SHIFTEN_6408_out0 ? v$MUX2_9349_out0 : v$FF4_11169_out0;
always @(posedge clk) v$FF4_11170_out0 <= v$SHIFTEN_6409_out0 ? v$MUX2_9350_out0 : v$FF4_11170_out0;
always @(posedge clk) v$FF4_11171_out0 <= v$SHIFTEN_6410_out0 ? v$MUX2_9351_out0 : v$FF4_11171_out0;
always @(posedge clk) v$FF4_11172_out0 <= v$SHIFTEN_6411_out0 ? v$MUX2_9352_out0 : v$FF4_11172_out0;
always @(posedge clk) v$FF4_11173_out0 <= v$SHIFTEN_6412_out0 ? v$MUX2_9353_out0 : v$FF4_11173_out0;
always @(posedge clk) v$FF9_11201_out0 <= v$FF10_9601_out0 ? v$G26_11199_out0 : v$FF9_11201_out0;
always @(posedge clk) v$FF9_11202_out0 <= v$FF10_9602_out0 ? v$G26_11200_out0 : v$FF9_11202_out0;
always @(posedge clk) v$FF1_11255_out0 <= v$SHIFTEN_6401_out0 ? v$MUX7_12679_out0 : v$FF1_11255_out0;
always @(posedge clk) v$FF1_11256_out0 <= v$SHIFTEN_6402_out0 ? v$MUX7_12680_out0 : v$FF1_11256_out0;
always @(posedge clk) v$FF1_11257_out0 <= v$SHIFTEN_6403_out0 ? v$MUX7_12681_out0 : v$FF1_11257_out0;
always @(posedge clk) v$FF1_11258_out0 <= v$SHIFTEN_6404_out0 ? v$MUX7_12682_out0 : v$FF1_11258_out0;
always @(posedge clk) v$FF1_11259_out0 <= v$SHIFTEN_6405_out0 ? v$MUX7_12683_out0 : v$FF1_11259_out0;
always @(posedge clk) v$FF1_11260_out0 <= v$SHIFTEN_6406_out0 ? v$MUX7_12684_out0 : v$FF1_11260_out0;
always @(posedge clk) v$FF1_11261_out0 <= v$SHIFTEN_6407_out0 ? v$MUX7_12685_out0 : v$FF1_11261_out0;
always @(posedge clk) v$FF1_11262_out0 <= v$SHIFTEN_6408_out0 ? v$MUX7_12686_out0 : v$FF1_11262_out0;
always @(posedge clk) v$FF1_11263_out0 <= v$SHIFTEN_6409_out0 ? v$MUX7_12687_out0 : v$FF1_11263_out0;
always @(posedge clk) v$FF1_11264_out0 <= v$SHIFTEN_6410_out0 ? v$MUX7_12688_out0 : v$FF1_11264_out0;
always @(posedge clk) v$FF1_11265_out0 <= v$SHIFTEN_6411_out0 ? v$MUX7_12689_out0 : v$FF1_11265_out0;
always @(posedge clk) v$FF1_11266_out0 <= v$SHIFTEN_6412_out0 ? v$MUX7_12690_out0 : v$FF1_11266_out0;
always @(posedge clk) v$REG9_11269_out0 <= v$HALT0_290_out0 ? v$RAMADDR0_12041_out0 : v$REG9_11269_out0;
always @(posedge clk) v$FF6_11336_out0 <= v$PHALT1_6182_out0;
always @(posedge clk) v$FF1_11343_out0 <= v$Shift_6566_out0 ? v$FF2_779_out0 : v$FF1_11343_out0;
always @(posedge clk) v$FF1_11344_out0 <= v$Shift_6567_out0 ? v$FF2_780_out0 : v$FF1_11344_out0;
always @(posedge clk) v$REG0_11406_out0 <= v$D1_9486_out0 ? v$DIN3_9801_out0 : v$REG0_11406_out0;
always @(posedge clk) v$REG0_11407_out0 <= v$D1_9487_out0 ? v$DIN3_9802_out0 : v$REG0_11407_out0;
always @(posedge clk) v$FF1_11440_out0 <= v$EXEC2_701_out0 ? v$S_6988_out0 : v$FF1_11440_out0;
always @(posedge clk) v$FF1_11441_out0 <= v$EXEC2_702_out0 ? v$S_6989_out0 : v$FF1_11441_out0;
always @(posedge clk) v$FF2_11450_out0 <= v$CAPTURE_207_out0 ? v$G1_9116_out0 : v$FF2_11450_out0;
always @(posedge clk) v$FF2_11451_out0 <= v$CAPTURE_208_out0 ? v$G1_9117_out0 : v$FF2_11451_out0;
always @(posedge clk) v$FF5_11452_out0 <= v$ShiftEN_5265_out0 ? v$MUX5_13207_out0 : v$FF5_11452_out0;
always @(posedge clk) v$FF5_11453_out0 <= v$ShiftEN_5266_out0 ? v$MUX5_13208_out0 : v$FF5_11453_out0;
always @(posedge clk) v$REG2_11460_out0 <= v$THRESHOLD$WRITE_4845_out0 ? v$THRESHOLD_10815_out0 : v$REG2_11460_out0;
always @(posedge clk) v$REG2_11461_out0 <= v$THRESHOLD$WRITE_4846_out0 ? v$THRESHOLD_10816_out0 : v$REG2_11461_out0;
always @(posedge clk) v$FF5_11521_out0 <= v$PHALT0_7479_out0;
always @(posedge clk) v$FF12_11522_out0 <= v$FF10_5406_out0;
always @(posedge clk) v$FF12_11523_out0 <= v$FF10_5407_out0;
always @(posedge clk) v$REG10_11541_out0 <= v$HALT0_290_out0 ? v$DATAIN0_7296_out0 : v$REG10_11541_out0;
always @(posedge clk) v$FF2_11724_out0 <= v$INTERRUPT1_12516_out0;
always @(posedge clk) v$FF2_11725_out0 <= v$INTERRUPT1_12517_out0;
always @(posedge clk) v$FF8_11778_out0 <= v$Shift_6566_out0 ? v$FF4_5735_out0 : v$FF8_11778_out0;
always @(posedge clk) v$FF8_11779_out0 <= v$Shift_6567_out0 ? v$FF4_5736_out0 : v$FF8_11779_out0;
v$ROM1_12254 I12254 (v$ROM1_12254_out0, v$ADDRESS_10499_out0, clk);
v$ROM1_12255 I12255 (v$ROM1_12255_out0, v$ADDRESS_10500_out0, clk);
always @(posedge clk) v$REG2_12278_out0 <= v$D1_9486_out2 ? v$DIN3_9801_out0 : v$REG2_12278_out0;
always @(posedge clk) v$REG2_12279_out0 <= v$D1_9487_out2 ? v$DIN3_9802_out0 : v$REG2_12279_out0;
always @(posedge clk) v$REG3_12548_out0 <= v$IR2$VALID_8838_out0 ? v$EQ1_11412_out0 : v$REG3_12548_out0;
always @(posedge clk) v$REG3_12549_out0 <= v$IR2$VALID_8839_out0 ? v$EQ1_11413_out0 : v$REG3_12549_out0;
always @(posedge clk) v$PCINTERRUPT_12603_out0 <= v$ININTERRUPT_433_out0 ? v$SUM_9219_out0 : v$PCINTERRUPT_12603_out0;
always @(posedge clk) v$PCINTERRUPT_12604_out0 <= v$ININTERRUPT_434_out0 ? v$SUM_9220_out0 : v$PCINTERRUPT_12604_out0;
always @(posedge clk) v$FF4_12634_out0 <= v$C1_3681_out0;
always @(posedge clk) v$FF4_12635_out0 <= v$C1_3682_out0;
always @(posedge clk) v$FF3_12851_out0 <= v$G29_5378_out0;
always @(posedge clk) v$FF3_12852_out0 <= v$G29_5379_out0;
always @(posedge clk) v$FF7_12855_out0 <= v$ShiftEN_5265_out0 ? v$MUX7_6471_out0 : v$FF7_12855_out0;
always @(posedge clk) v$FF7_12856_out0 <= v$ShiftEN_5266_out0 ? v$MUX7_6472_out0 : v$FF7_12856_out0;
always @(posedge clk) v$REG2_13074_out0 <= v$EXEC1_13169_out0 ? v$COUT$EXEC1_796_out0 : v$REG2_13074_out0;
always @(posedge clk) v$REG2_13075_out0 <= v$EXEC1_13170_out0 ? v$COUT$EXEC1_797_out0 : v$REG2_13075_out0;
always @(posedge clk) v$FF4_13119_out0 <= v$INTERRUPT3_1583_out0;
always @(posedge clk) v$FF4_13120_out0 <= v$INTERRUPT3_1584_out0;
always @(posedge clk) v$FF5_13141_out0 <= v$Shift_6566_out0 ? v$FF3_532_out0 : v$FF5_13141_out0;
always @(posedge clk) v$FF5_13142_out0 <= v$Shift_6567_out0 ? v$FF3_533_out0 : v$FF5_13142_out0;
always @(posedge clk) v$LSB$FF_13171_out0 <= v$EXEC2_461_out0 ? v$MUX5_12110_out0 : v$LSB$FF_13171_out0;
always @(posedge clk) v$LSB$FF_13172_out0 <= v$EXEC2_462_out0 ? v$MUX5_12111_out0 : v$LSB$FF_13172_out0;
always @(posedge clk) v$INT1_13185_out0 <= v$I1EN_13089_out0 ? v$SEL1_7748_out0 : v$INT1_13185_out0;
always @(posedge clk) v$INT1_13186_out0 <= v$I1EN_13090_out0 ? v$SEL1_7749_out0 : v$INT1_13186_out0;
always @(posedge clk) v$FF13_13193_out0 <= v$FF7_8410_out0;
always @(posedge clk) v$FF13_13194_out0 <= v$FF7_8411_out0;
always @(posedge clk) v$REG1_13298_out0 <= v$MODEWRITE_10070_out0 ? v$SEL1_12970_out0 : v$REG1_13298_out0;
always @(posedge clk) v$REG1_13299_out0 <= v$MODEWRITE_10071_out0 ? v$SEL1_12971_out0 : v$REG1_13299_out0;
assign v$C9_13388_out0 = 16'h0;
assign v$C9_13387_out0 = 16'h0;
assign v$C3_13206_out0 = 1'h0;
assign v$C3_13205_out0 = 1'h0;
assign v$C2_13021_out0 = 1'h0;
assign v$C2_13020_out0 = 1'h0;
assign v$CIN_12959_out0 = 1'h1;
assign v$CIN_12958_out0 = 1'h1;
assign v$CIN_12957_out0 = 1'h1;
assign v$CIN_12956_out0 = 1'h1;
assign v$CIN_12955_out0 = 1'h1;
assign v$CIN_12954_out0 = 1'h1;
assign v$CIN_12953_out0 = 1'h1;
assign v$CIN_12952_out0 = 1'h1;
assign v$C1_12940_out0 = 16'h0;
assign v$C1_12939_out0 = 16'h0;
assign v$C3_12864_out0 = 1'h0;
assign v$C3_12863_out0 = 1'h0;
assign v$C2_12782_out0 = 15'h0;
assign v$C2_12781_out0 = 15'h0;
assign v$C1_12497_out0 = 1'h0;
assign v$C1_12496_out0 = 1'h0;
assign v$C1_12495_out0 = 1'h0;
assign v$C1_12494_out0 = 1'h0;
assign v$C1_12493_out0 = 1'h0;
assign v$C1_12492_out0 = 1'h0;
assign v$C1_12160_out0 = 1'h1;
assign v$C1_12159_out0 = 1'h1;
assign v$C1_12158_out0 = 1'h1;
assign v$C1_12157_out0 = 1'h1;
assign v$C2_12079_out0 = 1'h0;
assign v$C2_12078_out0 = 1'h0;
assign v$C5_11972_out0 = 2'h2;
assign v$C5_11971_out0 = 2'h2;
assign v$C5_11970_out0 = 2'h2;
assign v$C5_11969_out0 = 2'h1;
assign v$C5_11968_out0 = 2'h2;
assign v$C5_11967_out0 = 2'h2;
assign v$C5_11966_out0 = 2'h2;
assign v$C5_11965_out0 = 2'h1;
assign v$C5_11964_out0 = 2'h2;
assign v$C5_11963_out0 = 2'h2;
assign v$C5_11962_out0 = 2'h2;
assign v$C5_11961_out0 = 2'h1;
assign v$C5_11960_out0 = 2'h2;
assign v$C5_11959_out0 = 2'h2;
assign v$C5_11958_out0 = 2'h2;
assign v$C5_11957_out0 = 2'h1;
assign v$C1_11891_out0 = 3'h0;
assign v$C1_11890_out0 = 3'h0;
assign v$C4_11603_out0 = 2'h1;
assign v$C4_11602_out0 = 2'h1;
assign v$C4_11601_out0 = 2'h1;
assign v$C4_11600_out0 = 2'h0;
assign v$C4_11599_out0 = 2'h1;
assign v$C4_11598_out0 = 2'h1;
assign v$C4_11597_out0 = 2'h1;
assign v$C4_11596_out0 = 2'h0;
assign v$C4_11595_out0 = 2'h1;
assign v$C4_11594_out0 = 2'h1;
assign v$C4_11593_out0 = 2'h1;
assign v$C4_11592_out0 = 2'h0;
assign v$C4_11591_out0 = 2'h1;
assign v$C4_11590_out0 = 2'h1;
assign v$C4_11589_out0 = 2'h1;
assign v$C4_11588_out0 = 2'h0;
assign v$C2_11447_out0 = 1'h1;
assign v$C2_11446_out0 = 1'h1;
assign v$C2_11445_out0 = 1'h1;
assign v$C2_11444_out0 = 1'h1;
assign v$C1_11443_out0 = 16'h0;
assign v$C1_11442_out0 = 16'h0;
assign v$C4_11433_out0 = 2'h0;
assign v$C4_11432_out0 = 2'h0;
assign v$C2_11419_out0 = 1'h0;
assign v$C2_11418_out0 = 1'h0;
assign v$C2_11417_out0 = 1'h0;
assign v$C2_11416_out0 = 1'h0;
assign v$C2_11392_out0 = 1'h1;
assign v$C2_11391_out0 = 1'h1;
assign v$C1_11390_out0 = 24'h0;
assign v$C1_11389_out0 = 24'h0;
assign v$C2_11175_out0 = 6'h1;
assign v$C2_11174_out0 = 6'h1;
assign v$C1_11145_out0 = 12'h0;
assign v$C1_11144_out0 = 12'h0;
assign v$C1_11127_out0 = 1'h1;
assign v$C1_11126_out0 = 1'h1;
assign v$C4_11122_out0 = 12'h0;
assign v$C4_11121_out0 = 12'h0;
assign v$C1_11028_out0 = 11'h0;
assign v$C1_11027_out0 = 11'h0;
assign v$C1_10983_out0 = 5'h1f;
assign v$C1_10982_out0 = 5'h1f;
assign v$C1_10976_out0 = 1'h0;
assign v$C1_10975_out0 = 1'h0;
assign v$C1_10974_out0 = 1'h0;
assign v$C1_10973_out0 = 1'h0;
assign v$C5_10889_out0 = 23'h0;
assign v$C5_10888_out0 = 23'h0;
assign v$C9_10582_out0 = 24'hffffff;
assign v$C9_10581_out0 = 24'hffffff;
assign v$C1_10548_out0 = 32'h0;
assign v$C1_10547_out0 = 32'h0;
assign v$C2_10486_out0 = 1'h0;
assign v$C2_10485_out0 = 1'h0;
assign v$C2_10484_out0 = 1'h0;
assign v$C2_10483_out0 = 1'h0;
assign v$C4_10178_out0 = 1'h1;
assign v$C4_10177_out0 = 1'h1;
assign v$C4_10176_out0 = 1'h1;
assign v$C4_10175_out0 = 1'h1;
assign v$C1_10161_out0 = 8'h0;
assign v$C1_10160_out0 = 8'h0;
assign v$C7_10013_out0 = 24'h0;
assign v$C7_10012_out0 = 24'h0;
assign v$C1_9651_out0 = 2'h3;
assign v$C1_9650_out0 = 2'h3;
assign v$C4_9420_out0 = 32'h0;
assign v$C4_9419_out0 = 32'h0;
assign v$C1_9391_out0 = 8'h0;
assign v$C1_9390_out0 = 8'h0;
assign v$C8_9179_out0 = 24'hffffff;
assign v$C8_9178_out0 = 24'hffffff;
assign v$C1_9154_out0 = 8'hff;
assign v$C1_9153_out0 = 5'h1f;
assign v$C1_9152_out0 = 8'hff;
assign v$C1_9151_out0 = 5'h1f;
assign v$C1_9150_out0 = 8'hff;
assign v$C1_9149_out0 = 5'h1f;
assign v$C1_9148_out0 = 8'hff;
assign v$C1_9147_out0 = 5'h1f;
assign v$C10_9111_out0 = 3'h0;
assign v$C10_9110_out0 = 3'h0;
assign v$C3_9096_out0 = 1'h1;
assign v$C3_9095_out0 = 1'h1;
assign v$C3_9094_out0 = 1'h1;
assign v$C3_9093_out0 = 1'h1;
assign v$C2_9088_out0 = 1'h0;
assign v$C2_9087_out0 = 1'h0;
assign v$C1_9015_out0 = 8'h0;
assign v$C1_9014_out0 = 8'h0;
assign v$C2_8961_out0 = 2'h1;
assign v$C2_8960_out0 = 2'h1;
assign v$C2_8900_out0 = 3'h0;
assign v$C2_8899_out0 = 3'h0;
assign v$C3_8773_out0 = 6'h0;
assign v$C3_8772_out0 = 6'h0;
assign v$C1_8497_out0 = 1'h0;
assign v$C1_8496_out0 = 1'h0;
assign v$C1_8475_out0 = 4'h0;
assign v$C1_8474_out0 = 4'h0;
assign v$C6_8187_out0 = 1'h1;
assign v$C6_8186_out0 = 1'h1;
assign v$C2_7981_out0 = 16'hffff;
assign v$C2_7980_out0 = 16'hffff;
assign v$C3_7979_out0 = 16'h0;
assign v$C3_7978_out0 = 16'h0;
assign v$C3_7505_out0 = 1'h0;
assign v$C3_7504_out0 = 1'h0;
assign v$C6_7407_out0 = 1'h0;
assign v$C6_7406_out0 = 1'h0;
assign v$C6_7405_out0 = 1'h0;
assign v$C6_7404_out0 = 1'h0;
assign v$C6_7403_out0 = 1'h0;
assign v$C6_7402_out0 = 1'h0;
assign v$C6_7401_out0 = 1'h0;
assign v$C6_7400_out0 = 1'h0;
assign v$C6_7399_out0 = 1'h0;
assign v$C6_7398_out0 = 1'h0;
assign v$C6_7397_out0 = 1'h0;
assign v$C6_7396_out0 = 1'h0;
assign v$C6_7395_out0 = 1'h0;
assign v$C6_7394_out0 = 1'h0;
assign v$C6_7393_out0 = 1'h0;
assign v$C6_7392_out0 = 1'h0;
assign v$C6_7391_out0 = 1'h0;
assign v$C6_7390_out0 = 1'h0;
assign v$C6_7389_out0 = 1'h0;
assign v$C6_7388_out0 = 1'h0;
assign v$C6_7387_out0 = 1'h0;
assign v$C6_7386_out0 = 1'h0;
assign v$C6_7385_out0 = 1'h0;
assign v$C6_7384_out0 = 1'h0;
assign v$C2_6725_out0 = 16'hffff;
assign v$C2_6724_out0 = 16'hffff;
assign v$C10_6198_out0 = 13'h0;
assign v$C10_6197_out0 = 13'h0;
assign v$C5_6005_out0 = 1'h1;
assign v$C5_6004_out0 = 1'h1;
assign v$C5_6003_out0 = 1'h1;
assign v$C5_6002_out0 = 1'h1;
assign v$C4_5742_out0 = 31'h0;
assign v$C4_5741_out0 = 15'h0;
assign v$C4_5740_out0 = 31'h0;
assign v$C4_5739_out0 = 15'h0;
assign v$C8_5699_out0 = 13'h0;
assign v$C8_5698_out0 = 13'h0;
assign v$C6_5556_out0 = 6'h1;
assign v$C6_5555_out0 = 6'h1;
assign v$C1_5485_out0 = 8'h0;
assign v$C1_5484_out0 = 4'h0;
assign v$C1_5483_out0 = 2'h0;
assign v$C1_5482_out0 = 1'h0;
assign v$C1_5481_out0 = 8'h0;
assign v$C1_5480_out0 = 4'h0;
assign v$C1_5479_out0 = 2'h0;
assign v$C1_5478_out0 = 1'h0;
assign v$C2_5341_out0 = 24'h0;
assign v$C2_5340_out0 = 24'h0;
assign v$C1_5268_out0 = 2'h2;
assign v$C1_5267_out0 = 2'h2;
assign v$C2_5168_out0 = 1'h1;
assign v$C2_5167_out0 = 1'h1;
assign v$C2_5166_out0 = 1'h1;
assign v$C2_5165_out0 = 1'h1;
assign v$C2_5164_out0 = 1'h1;
assign v$C2_5163_out0 = 1'h1;
assign v$C1_5007_out0 = 5'h0;
assign v$C1_5006_out0 = 5'h0;
assign v$C8_4880_out0 = 4'h0;
assign v$C8_4879_out0 = 4'h0;
assign v$C4_4631_out0 = 3'h0;
assign v$C4_4630_out0 = 3'h0;
assign v$C6_4551_out0 = 2'h3;
assign v$C6_4550_out0 = 2'h3;
assign v$C6_4549_out0 = 2'h3;
assign v$C6_4548_out0 = 2'h2;
assign v$C6_4547_out0 = 2'h3;
assign v$C6_4546_out0 = 2'h3;
assign v$C6_4545_out0 = 2'h3;
assign v$C6_4544_out0 = 2'h2;
assign v$C6_4543_out0 = 2'h3;
assign v$C6_4542_out0 = 2'h3;
assign v$C6_4541_out0 = 2'h3;
assign v$C6_4540_out0 = 2'h2;
assign v$C6_4539_out0 = 2'h3;
assign v$C6_4538_out0 = 2'h3;
assign v$C6_4537_out0 = 2'h3;
assign v$C6_4536_out0 = 2'h2;
assign v$C1_4455_out0 = 1'h0;
assign v$C1_4454_out0 = 1'h0;
assign v$C10_4404_out0 = 16'h0;
assign v$C10_4403_out0 = 16'h0;
assign v$C4_4392_out0 = 1'h0;
assign v$C4_4391_out0 = 1'h0;
assign v$C7_4040_out0 = 13'h0;
assign v$C7_4039_out0 = 13'h0;
assign v$C1_4026_out0 = 2'h0;
assign v$C1_4025_out0 = 4'h0;
assign v$C1_4024_out0 = 1'h0;
assign v$C1_4023_out0 = 8'h0;
assign v$C1_4022_out0 = 16'h0;
assign v$C1_4021_out0 = 2'h0;
assign v$C1_4020_out0 = 4'h0;
assign v$C1_4019_out0 = 1'h0;
assign v$C1_4018_out0 = 8'h0;
assign v$C1_4017_out0 = 16'h0;
assign v$C1_4016_out0 = 2'h0;
assign v$C1_4015_out0 = 4'h0;
assign v$C1_4014_out0 = 1'h0;
assign v$C1_4013_out0 = 8'h0;
assign v$C1_4012_out0 = 16'h0;
assign v$C1_4011_out0 = 4'h0;
assign v$C1_4010_out0 = 1'h0;
assign v$C1_4009_out0 = 16'h0;
assign v$C1_4008_out0 = 2'h0;
assign v$C1_4007_out0 = 8'h0;
assign v$C1_4006_out0 = 32'h0;
assign v$C1_4005_out0 = 4'h0;
assign v$C1_4004_out0 = 1'h0;
assign v$C1_4003_out0 = 16'h0;
assign v$C1_4002_out0 = 2'h0;
assign v$C1_4001_out0 = 8'h0;
assign v$C1_4000_out0 = 32'h0;
assign v$C1_3999_out0 = 2'h0;
assign v$C1_3998_out0 = 4'h0;
assign v$C1_3997_out0 = 1'h0;
assign v$C1_3996_out0 = 8'h0;
assign v$C1_3995_out0 = 16'h0;
assign v$C1_3994_out0 = 2'h0;
assign v$C1_3993_out0 = 4'h0;
assign v$C1_3992_out0 = 1'h0;
assign v$C1_3991_out0 = 8'h0;
assign v$C1_3990_out0 = 16'h0;
assign v$C1_3989_out0 = 2'h0;
assign v$C1_3988_out0 = 4'h0;
assign v$C1_3987_out0 = 1'h0;
assign v$C1_3986_out0 = 8'h0;
assign v$C1_3985_out0 = 16'h0;
assign v$C1_3984_out0 = 2'h0;
assign v$C1_3983_out0 = 4'h0;
assign v$C1_3982_out0 = 1'h0;
assign v$C1_3981_out0 = 8'h0;
assign v$C1_3980_out0 = 16'h0;
assign v$C1_3979_out0 = 4'h0;
assign v$C1_3978_out0 = 1'h0;
assign v$C1_3977_out0 = 16'h0;
assign v$C1_3976_out0 = 2'h0;
assign v$C1_3975_out0 = 8'h0;
assign v$C1_3974_out0 = 32'h0;
assign v$C1_3973_out0 = 4'h0;
assign v$C1_3972_out0 = 1'h0;
assign v$C1_3971_out0 = 16'h0;
assign v$C1_3970_out0 = 2'h0;
assign v$C1_3969_out0 = 8'h0;
assign v$C1_3968_out0 = 32'h0;
assign v$C1_3967_out0 = 2'h0;
assign v$C1_3966_out0 = 4'h0;
assign v$C1_3965_out0 = 1'h0;
assign v$C1_3964_out0 = 8'h0;
assign v$C1_3963_out0 = 16'h0;
assign v$C1_3960_out0 = 8'h81;
assign v$C1_3959_out0 = 5'h11;
assign v$C1_3958_out0 = 8'h81;
assign v$C1_3957_out0 = 5'h11;
assign v$C1_3682_out0 = 1'h1;
assign v$C1_3681_out0 = 1'h1;
assign v$C1_3658_out0 = 4'h0;
assign v$C1_3657_out0 = 4'h0;
assign v$C3_3632_out0 = 1'h1;
assign v$C3_3631_out0 = 1'h1;
assign v$C1_3100_out0 = 24'h0;
assign v$C1_3099_out0 = 24'h0;
assign v$C1_3098_out0 = 24'h0;
assign v$C1_3097_out0 = 24'h0;
assign v$C1_3096_out0 = 24'h0;
assign v$C1_3095_out0 = 24'h0;
assign v$C1_3094_out0 = 24'h0;
assign v$C1_3093_out0 = 24'h0;
assign v$C1_3013_out0 = 1'h1;
assign v$C1_3012_out0 = 1'h1;
assign v$C5_2812_out0 = 32'h0;
assign v$C5_2811_out0 = 32'h0;
assign v$C5_2695_out0 = 24'h0;
assign v$C5_2694_out0 = 24'h0;
assign v$C5_2693_out0 = 24'h0;
assign v$C5_2692_out0 = 24'h0;
assign v$C5_2691_out0 = 24'h0;
assign v$C5_2690_out0 = 24'h0;
assign v$C5_2689_out0 = 24'h0;
assign v$C5_2688_out0 = 24'h0;
assign v$C5_2687_out0 = 24'h0;
assign v$C5_2686_out0 = 24'h0;
assign v$C5_2685_out0 = 24'h0;
assign v$C5_2684_out0 = 24'h0;
assign v$C5_2683_out0 = 24'h0;
assign v$C5_2682_out0 = 24'h0;
assign v$C5_2681_out0 = 24'h0;
assign v$C5_2680_out0 = 24'h0;
assign v$C5_2679_out0 = 24'h0;
assign v$C5_2678_out0 = 24'h0;
assign v$C5_2677_out0 = 24'h0;
assign v$C5_2676_out0 = 24'h0;
assign v$C5_2675_out0 = 24'h0;
assign v$C5_2674_out0 = 24'h0;
assign v$C5_2673_out0 = 24'h0;
assign v$C5_2672_out0 = 24'h0;
assign v$C4_2468_out0 = 1'h1;
assign v$C4_2467_out0 = 1'h1;
assign v$C11_2341_out0 = 1'h0;
assign v$C11_2340_out0 = 1'h0;
assign v$C2_2337_out0 = 1'h1;
assign v$C2_2336_out0 = 1'h1;
assign v$C3_2012_out0 = 2'h0;
assign v$C3_2011_out0 = 2'h0;
assign v$C3_2010_out0 = 2'h0;
assign v$C3_2009_out0 = 2'h0;
assign v$C3_2008_out0 = 2'h0;
assign v$C3_2007_out0 = 2'h0;
assign v$C3_2006_out0 = 2'h0;
assign v$C3_2005_out0 = 2'h0;
assign v$C3_2004_out0 = 2'h0;
assign v$C3_2003_out0 = 2'h0;
assign v$C3_2002_out0 = 2'h0;
assign v$C3_2001_out0 = 2'h0;
assign v$C9_2000_out0 = 16'h0;
assign v$C9_1999_out0 = 16'h0;
assign v$C1_1780_out0 = 2'h0;
assign v$C1_1779_out0 = 2'h0;
assign v$C2_1737_out0 = 1'h1;
assign v$C2_1736_out0 = 1'h1;
assign v$C4_1693_out0 = 1'h1;
assign v$C4_1692_out0 = 1'h1;
assign v$C2_1569_out0 = 1'h0;
assign v$C2_1568_out0 = 1'h0;
assign v$C1_1546_out0 = 1'h1;
assign v$C1_1545_out0 = 1'h1;
assign v$C1_1544_out0 = 1'h1;
assign v$C1_1543_out0 = 1'h1;
assign v$C1_1542_out0 = 1'h1;
assign v$C1_1541_out0 = 1'h1;
assign v$C1_1540_out0 = 1'h1;
assign v$C1_1539_out0 = 1'h1;
assign v$C1_1538_out0 = 1'h1;
assign v$C1_1537_out0 = 1'h1;
assign v$C1_1536_out0 = 1'h1;
assign v$C1_1535_out0 = 1'h1;
assign v$C4_1380_out0 = 13'h0;
assign v$C4_1379_out0 = 13'h0;
assign v$C6_1360_out0 = 1'h1;
assign v$C6_1359_out0 = 1'h1;
assign v$C6_1358_out0 = 1'h1;
assign v$C6_1357_out0 = 1'h1;
assign v$C7_894_out0 = 16'h0;
assign v$C7_893_out0 = 16'h0;
assign v$C6_776_out0 = 1'h1;
assign v$C6_775_out0 = 1'h1;
assign v$C1_768_out0 = 8'hff;
assign v$C1_767_out0 = 8'hff;
assign v$C6_758_out0 = 13'h0;
assign v$C6_757_out0 = 13'h0;
assign v$C1_740_out0 = 1'h0;
assign v$C1_739_out0 = 1'h0;
assign v$C1_704_out0 = 1'h0;
assign v$C1_703_out0 = 1'h0;
assign v$C2_694_out0 = 1'h1;
assign v$C2_693_out0 = 1'h1;
assign v$C3_588_out0 = 1'h1;
assign v$C3_587_out0 = 1'h1;
assign v$C2_466_out0 = 1'h1;
assign v$C2_465_out0 = 1'h1;
assign v$C7_275_out0 = 1'h0;
assign v$C7_274_out0 = 1'h0;
assign v$C2_159_out0 = 2'h0;
assign v$C2_158_out0 = 4'h0;
assign v$C2_157_out0 = 1'h0;
assign v$C2_156_out0 = 8'h0;
assign v$C2_155_out0 = 16'h0;
assign v$C2_154_out0 = 2'h0;
assign v$C2_153_out0 = 4'h0;
assign v$C2_152_out0 = 1'h0;
assign v$C2_151_out0 = 8'h0;
assign v$C2_150_out0 = 16'h0;
assign v$C2_149_out0 = 2'h0;
assign v$C2_148_out0 = 4'h0;
assign v$C2_147_out0 = 1'h0;
assign v$C2_146_out0 = 8'h0;
assign v$C2_145_out0 = 16'h0;
assign v$C2_144_out0 = 4'h0;
assign v$C2_143_out0 = 1'h0;
assign v$C2_142_out0 = 16'h0;
assign v$C2_141_out0 = 2'h0;
assign v$C2_140_out0 = 8'h0;
assign v$C2_139_out0 = 32'h0;
assign v$C2_138_out0 = 4'h0;
assign v$C2_137_out0 = 1'h0;
assign v$C2_136_out0 = 16'h0;
assign v$C2_135_out0 = 2'h0;
assign v$C2_134_out0 = 8'h0;
assign v$C2_133_out0 = 32'h0;
assign v$C2_132_out0 = 2'h0;
assign v$C2_131_out0 = 4'h0;
assign v$C2_130_out0 = 1'h0;
assign v$C2_129_out0 = 8'h0;
assign v$C2_128_out0 = 16'h0;
assign v$C2_127_out0 = 2'h0;
assign v$C2_126_out0 = 4'h0;
assign v$C2_125_out0 = 1'h0;
assign v$C2_124_out0 = 8'h0;
assign v$C2_123_out0 = 16'h0;
assign v$C2_122_out0 = 2'h0;
assign v$C2_121_out0 = 4'h0;
assign v$C2_120_out0 = 1'h0;
assign v$C2_119_out0 = 8'h0;
assign v$C2_118_out0 = 16'h0;
assign v$C2_117_out0 = 2'h0;
assign v$C2_116_out0 = 4'h0;
assign v$C2_115_out0 = 1'h0;
assign v$C2_114_out0 = 8'h0;
assign v$C2_113_out0 = 16'h0;
assign v$C2_112_out0 = 4'h0;
assign v$C2_111_out0 = 1'h0;
assign v$C2_110_out0 = 16'h0;
assign v$C2_109_out0 = 2'h0;
assign v$C2_108_out0 = 8'h0;
assign v$C2_107_out0 = 32'h0;
assign v$C2_106_out0 = 4'h0;
assign v$C2_105_out0 = 1'h0;
assign v$C2_104_out0 = 16'h0;
assign v$C2_103_out0 = 2'h0;
assign v$C2_102_out0 = 8'h0;
assign v$C2_101_out0 = 32'h0;
assign v$C2_100_out0 = 2'h0;
assign v$C2_99_out0 = 4'h0;
assign v$C2_98_out0 = 1'h0;
assign v$C2_97_out0 = 8'h0;
assign v$C2_96_out0 = 16'h0;
assign v$C5_7_out0 = 13'h0;
assign v$C5_6_out0 = 13'h0;
assign v$G3_22_out0 = !(v$FF0_3399_out0 || v$FF1_6586_out0);
assign v$G3_23_out0 = !(v$FF0_3400_out0 || v$FF1_6587_out0);
assign v$G2_62_out0 = ! v$FF1_178_out0;
assign v$G2_63_out0 = ! v$FF1_179_out0;
assign v$Q0_74_out0 = v$FF0_6397_out0;
assign v$Q0_75_out0 = v$FF0_6398_out0;
assign v$SIN_87_out0 = v$C7_274_out0;
assign v$SIN_93_out0 = v$C7_275_out0;
assign v$G58_162_out0 = ! v$FF5_3159_out0;
assign v$G58_163_out0 = ! v$FF5_3160_out0;
assign v$_525_out0 = { v$FF0_6397_out0,v$FF1_1433_out0 };
assign v$_526_out0 = { v$FF0_6398_out0,v$FF1_1434_out0 };
assign v$G2_529_out0 = ((v$FF5_13141_out0 && !v$FF3_532_out0) || (!v$FF5_13141_out0) && v$FF3_532_out0);
assign v$G2_530_out0 = ((v$FF5_13142_out0 && !v$FF3_533_out0) || (!v$FF5_13142_out0) && v$FF3_533_out0);
assign v$INITIAL$FETCH$OCCURRED_759_out0 = v$FF4_12634_out0;
assign v$INITIAL$FETCH$OCCURRED_760_out0 = v$FF4_12635_out0;
assign v$CIN$EXEC1_792_out0 = v$REG2_13074_out0;
assign v$CIN$EXEC1_793_out0 = v$REG2_13075_out0;
assign v$PHALT_834_out0 = v$REG2_3503_out0;
assign v$SELOUT_900_out0 = v$REG8_2804_out0;
assign v$SOUT1_1068_out0 = v$FF4_11162_out0;
assign v$SOUT1_1069_out0 = v$FF4_11163_out0;
assign v$SOUT1_1070_out0 = v$FF4_11164_out0;
assign v$SOUT1_1071_out0 = v$FF4_11165_out0;
assign v$SOUT1_1072_out0 = v$FF4_11166_out0;
assign v$SOUT1_1073_out0 = v$FF4_11167_out0;
assign v$SOUT1_1074_out0 = v$FF4_11168_out0;
assign v$SOUT1_1075_out0 = v$FF4_11169_out0;
assign v$SOUT1_1076_out0 = v$FF4_11170_out0;
assign v$SOUT1_1077_out0 = v$FF4_11171_out0;
assign v$SOUT1_1078_out0 = v$FF4_11172_out0;
assign v$SOUT1_1079_out0 = v$FF4_11173_out0;
assign v$I2P_1179_out0 = v$FF2_11450_out0;
assign v$I2P_1180_out0 = v$FF2_11451_out0;
assign v$_1185_out0 = { v$FF7_12855_out0,v$FF8_5529_out0 };
assign v$_1186_out0 = { v$FF7_12856_out0,v$FF8_5530_out0 };
assign v$PIPELINERESTART_1353_out0 = v$FF1_2_out0;
assign v$PIPELINERESTART_1354_out0 = v$FF1_3_out0;
assign v$G4_1665_out0 = ((v$FF7_9941_out0 && !v$FF6_6215_out0) || (!v$FF7_9941_out0) && v$FF6_6215_out0);
assign v$G4_1666_out0 = ((v$FF7_9942_out0 && !v$FF6_6216_out0) || (!v$FF7_9942_out0) && v$FF6_6216_out0);
assign v$LEFT$SHIT_1800_out0 = v$C6_1357_out0;
assign v$LEFT$SHIT_1801_out0 = v$C4_10175_out0;
assign v$LEFT$SHIT_1802_out0 = v$C2_11444_out0;
assign v$LEFT$SHIT_1803_out0 = v$C5_6002_out0;
assign v$LEFT$SHIT_1804_out0 = v$C1_12157_out0;
assign v$LEFT$SHIT_1805_out0 = v$C3_9093_out0;
assign v$LEFT$SHIT_1806_out0 = v$C6_1358_out0;
assign v$LEFT$SHIT_1807_out0 = v$C4_10176_out0;
assign v$LEFT$SHIT_1808_out0 = v$C2_11445_out0;
assign v$LEFT$SHIT_1809_out0 = v$C5_6003_out0;
assign v$LEFT$SHIT_1810_out0 = v$C1_12158_out0;
assign v$LEFT$SHIT_1811_out0 = v$C3_9094_out0;
assign v$LEFT$SHIT_1832_out0 = v$C6_1359_out0;
assign v$LEFT$SHIT_1833_out0 = v$C4_10177_out0;
assign v$LEFT$SHIT_1834_out0 = v$C2_11446_out0;
assign v$LEFT$SHIT_1835_out0 = v$C5_6004_out0;
assign v$LEFT$SHIT_1836_out0 = v$C1_12159_out0;
assign v$LEFT$SHIT_1837_out0 = v$C3_9095_out0;
assign v$LEFT$SHIT_1838_out0 = v$C6_1360_out0;
assign v$LEFT$SHIT_1839_out0 = v$C4_10178_out0;
assign v$LEFT$SHIT_1840_out0 = v$C2_11447_out0;
assign v$LEFT$SHIT_1841_out0 = v$C5_6005_out0;
assign v$LEFT$SHIT_1842_out0 = v$C1_12160_out0;
assign v$LEFT$SHIT_1843_out0 = v$C3_9096_out0;
assign v$Q2_1883_out0 = v$FF2_10772_out0;
assign v$Q2_1884_out0 = v$FF2_10773_out0;
assign v$R0_1977_out0 = v$REG0_11406_out0;
assign v$R0_1978_out0 = v$REG0_11407_out0;
assign v$S$REG_2143_out0 = v$REG1_7183_out0;
assign v$S$REG_2144_out0 = v$REG1_7184_out0;
assign v$A$SAVED_2413_out0 = v$REG1_457_out0;
assign v$A$SAVED_2414_out0 = v$REG1_458_out0;
assign v$_2493_out0 = { v$FF7_9941_out0,v$FF6_6215_out0 };
assign v$_2494_out0 = { v$FF7_9942_out0,v$FF6_6216_out0 };
assign {v$A1_2728_out1,v$A1_2728_out0 } = v$REG1_10179_out0 + v$C2_11174_out0 + v$C1_739_out0;
assign {v$A1_2729_out1,v$A1_2729_out0 } = v$REG1_10180_out0 + v$C2_11175_out0 + v$C1_740_out0;
assign v$Q1_3089_out0 = v$FF1_6568_out0;
assign v$Q1_3090_out0 = v$FF1_6569_out0;
assign v$B$SAVED_3161_out0 = v$REG2_10886_out0;
assign v$B$SAVED_3162_out0 = v$REG2_10887_out0;
assign v$_3288_out0 = v$REG1_13298_out0[2:0];
assign v$_3288_out1 = v$REG1_13298_out0[3:1];
assign v$_3289_out0 = v$REG1_13299_out0[2:0];
assign v$_3289_out1 = v$REG1_13299_out0[3:1];
assign v$Wordlength_3514_out0 = v$REG1_10179_out0 == 6'h27;
assign v$Wordlength_3515_out0 = v$REG1_10180_out0 == 6'h27;
assign v$G2_3619_out0 = ((v$FF0_3399_out0 && !v$FF1_6586_out0) || (!v$FF0_3399_out0) && v$FF1_6586_out0);
assign v$G2_3620_out0 = ((v$FF0_3400_out0 && !v$FF1_6587_out0) || (!v$FF0_3400_out0) && v$FF1_6587_out0);
assign v$OUT_3625_out0 = v$ROM1_12254_out0;
assign v$OUT_3626_out0 = v$ROM1_12255_out0;
assign v$Q2_3703_out0 = v$FF2_9998_out0;
assign v$Q2_3704_out0 = v$FF2_9999_out0;
assign v$G17_3720_out0 = ! v$FF2_11724_out0;
assign v$G17_3721_out0 = ! v$FF2_11725_out0;
assign v$STALL$PREV$CYCLE_3798_out0 = v$FF7_8410_out0;
assign v$STALL$PREV$CYCLE_3799_out0 = v$FF7_8411_out0;
assign v$STALL$PREV$PREV_3829_out0 = v$FF13_13193_out0;
assign v$STALL$PREV$PREV_3830_out0 = v$FF13_13194_out0;
assign v$IR$READ$IN$PREV$CYCLE_4206_out0 = v$REG2_10321_out0;
assign v$IR$READ$IN$PREV$CYCLE_4207_out0 = v$REG2_10322_out0;
assign v$I1P_4447_out0 = v$FF3_5109_out0;
assign v$I1P_4448_out0 = v$FF3_5110_out0;
assign v$EQ1_4702_out0 = v$REG2_11460_out0 == 16'h0;
assign v$EQ1_4703_out0 = v$REG2_11461_out0 == 16'h0;
assign v$PHALT1$PREV_4956_out0 = v$FF6_11336_out0;
assign v$G20_4995_out0 = ((v$FF7_12855_out0 && !v$FF8_5529_out0) || (!v$FF7_12855_out0) && v$FF8_5529_out0);
assign v$G20_4996_out0 = ((v$FF7_12856_out0 && !v$FF8_5530_out0) || (!v$FF7_12856_out0) && v$FF8_5530_out0);
assign v$PHALT0$PREV_5150_out0 = v$FF5_11521_out0;
assign v$HALT$PREV$PREV$PREV_5277_out0 = v$FF15_8373_out0;
assign v$HALT$PREV$PREV$PREV_5278_out0 = v$FF15_8374_out0;
assign v$_5279_out0 = { v$FF3_227_out0,v$FF4_1281_out0 };
assign v$_5280_out0 = { v$FF3_228_out0,v$FF4_1282_out0 };
assign v$LSB_5342_out0 = v$LSB$FF_13171_out0;
assign v$LSB_5343_out0 = v$LSB$FF_13172_out0;
assign v$LSBS_5438_out0 = v$REG1_6863_out0;
assign v$LSBS_5439_out0 = v$REG1_6864_out0;
assign v$R2_5454_out0 = v$REG2_12278_out0;
assign v$R2_5455_out0 = v$REG2_12279_out0;
assign v$PHALT1_6182_out0 = v$REG14_3705_out0;
assign v$I3P_6221_out0 = v$FF1_4163_out0;
assign v$I3P_6222_out0 = v$FF1_4164_out0;
assign v$G23_6381_out0 = ((v$FF1_6417_out0 && !v$FF2_1717_out0) || (!v$FF1_6417_out0) && v$FF2_1717_out0);
assign v$G23_6382_out0 = ((v$FF1_6418_out0 && !v$FF2_1718_out0) || (!v$FF1_6418_out0) && v$FF2_1718_out0);
assign v$SHIFTEN_6401_out0 = v$C1_1535_out0;
assign v$SHIFTEN_6402_out0 = v$C1_1536_out0;
assign v$SHIFTEN_6403_out0 = v$C1_1537_out0;
assign v$SHIFTEN_6404_out0 = v$C1_1538_out0;
assign v$SHIFTEN_6405_out0 = v$C1_1539_out0;
assign v$SHIFTEN_6406_out0 = v$C1_1540_out0;
assign v$SHIFTEN_6407_out0 = v$C1_1541_out0;
assign v$SHIFTEN_6408_out0 = v$C1_1542_out0;
assign v$SHIFTEN_6409_out0 = v$C1_1543_out0;
assign v$SHIFTEN_6410_out0 = v$C1_1544_out0;
assign v$SHIFTEN_6411_out0 = v$C1_1545_out0;
assign v$SHIFTEN_6412_out0 = v$C1_1546_out0;
assign v$_6431_out0 = { v$FF8_11778_out0,v$FF4_5735_out0 };
assign v$_6432_out0 = { v$FF8_11779_out0,v$FF4_5736_out0 };
assign v$RecievedParity_6514_out0 = v$FF7_5594_out0;
assign v$RecievedParity_6515_out0 = v$FF7_5595_out0;
assign v$G31_6588_out0 = ! v$FF4_13119_out0;
assign v$G31_6589_out0 = ! v$FF4_13120_out0;
assign v$G63_6734_out0 = ! v$FF8_6889_out0;
assign v$G63_6735_out0 = ! v$FF8_6890_out0;
assign v$I0P_6869_out0 = v$FF4_2489_out0;
assign v$I0P_6870_out0 = v$FF4_2490_out0;
assign v$OUTPUT_6891_out0 = v$FF1_3605_out0;
assign v$OUTPUT_6892_out0 = v$FF1_3606_out0;
assign v$HALT$PREV_6935_out0 = v$FF10_5406_out0;
assign v$HALT$PREV_6936_out0 = v$FF10_5407_out0;
assign v$R3_7072_out0 = v$REG3_7255_out0;
assign v$R3_7073_out0 = v$REG3_7256_out0;
assign v$Q1_7197_out0 = v$FF1_467_out0;
assign v$Q1_7198_out0 = v$FF1_468_out0;
assign v$PHALT0_7479_out0 = v$REG13_248_out0;
assign v$ISINTERRUPTED_7651_out0 = v$FF1_8718_out0;
assign v$ISINTERRUPTED_7652_out0 = v$FF1_8719_out0;
assign v$G21_7669_out0 = ((v$FF5_11452_out0 && !v$FF6_10631_out0) || (!v$FF5_11452_out0) && v$FF6_10631_out0);
assign v$G21_7670_out0 = ((v$FF5_11453_out0 && !v$FF6_10632_out0) || (!v$FF5_11453_out0) && v$FF6_10632_out0);
assign v$INT2_7675_out0 = v$C3_7504_out0;
assign v$INT2_7676_out0 = v$C3_7505_out0;
assign v$G24_7868_out0 = ! v$FF3_10341_out0;
assign v$G24_7869_out0 = ! v$FF3_10342_out0;
assign v$LASTQ_7873_out0 = v$FF2_8662_out0;
assign v$LASTQ_7874_out0 = v$FF2_8663_out0;
assign v$LASTQ_7875_out0 = v$FF2_8664_out0;
assign v$LASTQ_7876_out0 = v$FF2_8665_out0;
assign v$LASTQ_7877_out0 = v$FF2_8666_out0;
assign v$LASTQ_7878_out0 = v$FF2_8667_out0;
assign v$LASTQ_7879_out0 = v$FF2_8668_out0;
assign v$LASTQ_7880_out0 = v$FF2_8669_out0;
assign v$LASTQ_7881_out0 = v$FF2_8670_out0;
assign v$LASTQ_7882_out0 = v$FF2_8671_out0;
assign v$LASTQ_7883_out0 = v$FF2_8672_out0;
assign v$LASTQ_7884_out0 = v$FF2_8673_out0;
assign v$LASTQ_7885_out0 = v$FF2_8674_out0;
assign v$LASTQ_7886_out0 = v$FF2_8675_out0;
assign v$LASTQ_7887_out0 = v$FF2_8676_out0;
assign v$LASTQ_7888_out0 = v$FF2_8677_out0;
assign v$LASTQ_7889_out0 = v$FF2_8678_out0;
assign v$LASTQ_7890_out0 = v$FF2_8679_out0;
assign v$LASTQ_7891_out0 = v$FF2_8680_out0;
assign v$LASTQ_7892_out0 = v$FF2_8681_out0;
assign v$LASTQ_7893_out0 = v$FF2_8682_out0;
assign v$LASTQ_7894_out0 = v$FF2_8683_out0;
assign v$PCHALT_8399_out0 = v$REG1_6069_out0;
assign v$LEFT$SHIFT_8476_out0 = v$C3_12863_out0;
assign v$LEFT$SHIFT_8477_out0 = v$C11_2340_out0;
assign v$LEFT$SHIFT_8478_out0 = v$C2_12078_out0;
assign v$LEFT$SHIFT_8479_out0 = v$C3_587_out0;
assign v$LEFT$SHIFT_8480_out0 = v$C3_12864_out0;
assign v$LEFT$SHIFT_8481_out0 = v$C11_2341_out0;
assign v$LEFT$SHIFT_8482_out0 = v$C2_12079_out0;
assign v$LEFT$SHIFT_8483_out0 = v$C3_588_out0;
assign v$RMORIGINAL_8617_out0 = v$REG1_9488_out0;
assign v$RMORIGINAL_8618_out0 = v$REG1_9489_out0;
assign v$G1_8760_out0 = ! v$FF0_3399_out0;
assign v$G1_8761_out0 = ! v$FF0_3400_out0;
assign v$VALID$PREV_9000_out0 = v$FF14_7185_out0;
assign v$VALID$PREV_9001_out0 = v$FF14_7186_out0;
assign v$CARRY_9008_out0 = v$FF1_6867_out0;
assign v$CARRY_9009_out0 = v$FF1_6868_out0;
assign v$Q0_9249_out0 = v$FF0_374_out0;
assign v$Q0_9250_out0 = v$FF0_375_out0;
assign v$R1_9296_out0 = v$REG1_3286_out0;
assign v$R1_9297_out0 = v$REG1_3287_out0;
assign v$Q1_9713_out0 = v$FF1_1433_out0;
assign v$Q1_9714_out0 = v$FF1_1434_out0;
assign v$G1_9855_out0 = ! v$FF1_4029_out0;
assign v$G1_9856_out0 = ! v$FF1_4030_out0;
assign v$ADDRESS_9958_out0 = v$REG2_376_out0;
assign v$ADDRESS_9959_out0 = v$REG2_377_out0;
assign v$G5_10022_out0 = ((v$FF8_11778_out0 && !v$FF4_5735_out0) || (!v$FF8_11778_out0) && v$FF4_5735_out0);
assign v$G5_10023_out0 = ((v$FF8_11779_out0 && !v$FF4_5736_out0) || (!v$FF8_11779_out0) && v$FF4_5736_out0);
assign v$_10125_out0 = { v$FF1_6417_out0,v$FF2_1717_out0 };
assign v$_10126_out0 = { v$FF1_6418_out0,v$FF2_1718_out0 };
assign {v$A2_10173_out1,v$A2_10173_out0 } = v$REG2_376_out0 + v$C6_5555_out0 + v$C4_4391_out0;
assign {v$A2_10174_out1,v$A2_10174_out0 } = v$REG2_377_out0 + v$C6_5556_out0 + v$C4_4392_out0;
assign v$_10228_out0 = { v$FF1_11343_out0,v$FF2_779_out0 };
assign v$_10229_out0 = { v$FF1_11344_out0,v$FF2_780_out0 };
assign v$G71_10591_out0 = ! v$FF4_5562_out0;
assign v$G71_10592_out0 = ! v$FF4_5563_out0;
assign v$LSBS_10623_out0 = v$REG1_6141_out0;
assign v$LSBS_10624_out0 = v$REG1_6142_out0;
assign v$EQ1_10629_out0 = v$REG1_10179_out0 == 6'h1e;
assign v$EQ1_10630_out0 = v$REG1_10180_out0 == 6'h1e;
assign v$SAVED_10674_out0 = v$REG3_4759_out0;
assign v$SAVED_10675_out0 = v$REG3_4760_out0;
assign v$G3_11055_out0 = ((v$FF1_11343_out0 && !v$FF2_779_out0) || (!v$FF1_11343_out0) && v$FF2_779_out0);
assign v$G3_11056_out0 = ((v$FF1_11344_out0 && !v$FF2_780_out0) || (!v$FF1_11344_out0) && v$FF2_780_out0);
assign v$G52_11142_out0 = ! v$FF4_4776_out0;
assign v$G52_11143_out0 = ! v$FF4_4777_out0;
assign v$_11152_out0 = { v$FF5_11452_out0,v$FF6_10631_out0 };
assign v$_11153_out0 = { v$FF5_11453_out0,v$FF6_10632_out0 };
assign v$STATE_11196_out0 = v$FF1_3605_out0;
assign v$STATE_11197_out0 = v$FF1_3606_out0;
assign v$STATE_11198_out0 = v$REG1_4808_out0;
assign v$IR2_11640_out0 = v$REG4_4650_out0;
assign v$IR2_11641_out0 = v$REG4_4651_out0;
assign v$G24_12076_out0 = ((v$FF3_227_out0 && !v$FF4_1281_out0) || (!v$FF3_227_out0) && v$FF4_1281_out0);
assign v$G24_12077_out0 = ((v$FF3_228_out0 && !v$FF4_1282_out0) || (!v$FF3_228_out0) && v$FF4_1282_out0);
assign v$A_12094_out0 = v$REG1_9161_out0;
assign v$A_12095_out0 = v$REG1_9162_out0;
assign v$Q2_12285_out0 = v$FF2_3000_out0;
assign v$Q2_12286_out0 = v$FF2_3001_out0;
assign v$B_12739_out0 = v$REG2_11460_out0;
assign v$B_12740_out0 = v$REG2_11461_out0;
assign v$HALT$PREV$PREV_12829_out0 = v$FF12_11522_out0;
assign v$HALT$PREV$PREV_12830_out0 = v$FF12_11523_out0;
assign v$INT3_12861_out0 = v$C2_13020_out0;
assign v$INT3_12862_out0 = v$C2_13021_out0;
assign v$SOUT_12929_out0 = v$FF1_6417_out0;
assign v$SOUT_12930_out0 = v$FF1_6418_out0;
assign v$AUTODISABLE_12944_out0 = v$FF3_12851_out0;
assign v$AUTODISABLE_12945_out0 = v$FF3_12852_out0;
assign v$Q3_12999_out0 = v$FF3_11154_out0;
assign v$Q3_13000_out0 = v$FF3_11155_out0;
assign v$EPARITY_13014_out0 = v$FF9_11201_out0;
assign v$EPARITY_13015_out0 = v$FF9_11202_out0;
assign v$Q0_13018_out0 = v$FF0_2992_out0;
assign v$Q0_13019_out0 = v$FF0_2993_out0;
assign v$_13097_out0 = { v$FF5_13141_out0,v$FF3_532_out0 };
assign v$_13098_out0 = { v$FF5_13142_out0,v$FF3_533_out0 };
assign v$Q3_13107_out0 = v$FF3_7189_out0;
assign v$Q3_13108_out0 = v$FF3_7190_out0;
assign v$_13131_out0 = v$REG1_2760_out0[3:0];
assign v$_13131_out1 = v$REG1_2760_out0[7:4];
assign v$_13132_out0 = v$REG1_2761_out0[3:0];
assign v$_13132_out1 = v$REG1_2761_out0[7:4];
assign v$OUTPUT_13145_out0 = v$REG1_4808_out0;
assign v$G1_30_out0 = v$Wordlength_3514_out0 || v$G2_62_out0;
assign v$G1_31_out0 = v$Wordlength_3515_out0 || v$G2_63_out0;
assign v$SIN_84_out0 = v$SOUT1_1069_out0;
assign v$SIN_85_out0 = v$SOUT1_1072_out0;
assign v$SIN_86_out0 = v$SOUT1_1073_out0;
assign v$SIN_88_out0 = v$SOUT1_1071_out0;
assign v$SIN_89_out0 = v$SOUT1_1068_out0;
assign v$SIN_90_out0 = v$SOUT1_1075_out0;
assign v$SIN_91_out0 = v$SOUT1_1078_out0;
assign v$SIN_92_out0 = v$SOUT1_1079_out0;
assign v$SIN_94_out0 = v$SOUT1_1077_out0;
assign v$SIN_95_out0 = v$SOUT1_1074_out0;
assign v$_749_out0 = v$A_12094_out0[7:0];
assign v$_749_out1 = v$A_12094_out0[15:8];
assign v$_750_out0 = v$A_12095_out0[7:0];
assign v$_750_out1 = v$A_12095_out0[15:8];
assign v$G1_794_out0 = ! v$Q0_13018_out0;
assign v$G1_795_out0 = ! v$Q0_13019_out0;
assign v$IR2_929_out0 = v$IR2_11640_out0;
assign v$IR2_930_out0 = v$IR2_11641_out0;
assign v$_1005_out0 = { v$Q0_13018_out0,v$Q1_3089_out0 };
assign v$_1006_out0 = { v$Q0_13019_out0,v$Q1_3090_out0 };
assign v$G8_1189_out0 = ! v$Q1_9713_out0;
assign v$G8_1190_out0 = ! v$Q1_9714_out0;
assign v$I1P_1427_out0 = v$I1P_4447_out0;
assign v$I1P_1428_out0 = v$I1P_4448_out0;
assign v$IR2_1700_out0 = v$IR2_11640_out0;
assign v$IR2_1701_out0 = v$IR2_11641_out0;
assign v$G18_1749_out0 = ! v$ISINTERRUPTED_7651_out0;
assign v$G18_1750_out0 = ! v$ISINTERRUPTED_7652_out0;
assign v$END4_1971_out0 = v$LASTQ_7883_out0;
assign v$END4_1972_out0 = v$LASTQ_7894_out0;
assign v$G6_2050_out0 = ((v$Q0_74_out0 && !v$Q1_9713_out0) || (!v$Q0_74_out0) && v$Q1_9713_out0);
assign v$G6_2051_out0 = ((v$Q0_75_out0 && !v$Q1_9714_out0) || (!v$Q0_75_out0) && v$Q1_9714_out0);
assign v$INTERRUPT3_2210_out0 = v$INT3_12861_out0;
assign v$INTERRUPT3_2211_out0 = v$INT3_12862_out0;
assign v$INTERRUPT2_2562_out0 = v$INT2_7675_out0;
assign v$INTERRUPT2_2563_out0 = v$INT2_7676_out0;
assign v$B$SAVED_2592_out0 = v$B$SAVED_3161_out0;
assign v$B$SAVED_2593_out0 = v$B$SAVED_3162_out0;
assign v$CIN_2595_out0 = v$CIN$EXEC1_792_out0;
assign v$CIN_2607_out0 = v$CIN$EXEC1_793_out0;
assign v$OFF_2756_out0 = v$EQ1_4702_out0;
assign v$OFF_2757_out0 = v$EQ1_4703_out0;
assign v$G22_2984_out0 = ((v$Q1_7197_out0 && !v$Q0_9249_out0) || (!v$Q1_7197_out0) && v$Q0_9249_out0);
assign v$G22_2985_out0 = ((v$Q1_7198_out0 && !v$Q0_9250_out0) || (!v$Q1_7198_out0) && v$Q0_9250_out0);
assign v$G35_2986_out0 = v$Q1_3089_out0 && v$Q0_13018_out0;
assign v$G35_2987_out0 = v$Q1_3090_out0 && v$Q0_13019_out0;
assign v$I0P_3002_out0 = v$I0P_6869_out0;
assign v$I0P_3003_out0 = v$I0P_6870_out0;
assign v$B$SAVED_3014_out0 = v$B$SAVED_3161_out0;
assign v$B$SAVED_3015_out0 = v$B$SAVED_3162_out0;
assign v$G48_3270_out0 = ! v$STALL$PREV$CYCLE_3798_out0;
assign v$G48_3271_out0 = ! v$STALL$PREV$CYCLE_3799_out0;
assign v$G87_3518_out0 = ! v$PHALT0_7479_out0;
assign v$_3718_out0 = { v$_10125_out0,v$_5279_out0 };
assign v$_3719_out0 = { v$_10126_out0,v$_5280_out0 };
assign v$_3760_out0 = { v$_13097_out0,v$_10228_out0 };
assign v$_3761_out0 = { v$_13098_out0,v$_10229_out0 };
assign v$SERIALIN_3766_out0 = v$SOUT_12929_out0;
assign v$SERIALIN_3767_out0 = v$SOUT_12930_out0;
assign v$SEL6_3784_out0 = v$SAVED_10674_out0[35:12];
assign v$SEL6_3785_out0 = v$SAVED_10675_out0[35:12];
assign v$PIPELINE$RESTART_4073_out0 = v$PIPELINERESTART_1353_out0;
assign v$PIPELINE$RESTART_4074_out0 = v$PIPELINERESTART_1354_out0;
assign v$RECIEVEDPARITY_4231_out0 = v$RecievedParity_6514_out0;
assign v$RECIEVEDPARITY_4232_out0 = v$RecievedParity_6515_out0;
assign v$G64_4407_out0 = v$HALT$PREV_6935_out0 && v$STALL$PREV$PREV_3829_out0;
assign v$G64_4408_out0 = v$HALT$PREV_6936_out0 && v$STALL$PREV$PREV_3830_out0;
assign v$END1_4730_out0 = v$LASTQ_7882_out0;
assign v$END1_4731_out0 = v$LASTQ_7893_out0;
assign v$END1_4747_out0 = v$A2_10173_out1;
assign v$END1_4748_out0 = v$A2_10174_out1;
assign v$_4782_out0 = { v$_11152_out0,v$_1185_out0 };
assign v$_4783_out0 = { v$_11153_out0,v$_1186_out0 };
assign v$G22_4865_out0 = ((v$G21_7669_out0 && !v$G20_4995_out0) || (!v$G21_7669_out0) && v$G20_4995_out0);
assign v$G22_4866_out0 = ((v$G21_7670_out0 && !v$G20_4996_out0) || (!v$G21_7670_out0) && v$G20_4996_out0);
assign v$I2P_5068_out0 = v$I2P_1179_out0;
assign v$I2P_5069_out0 = v$I2P_1180_out0;
assign v$R3TEST_5094_out0 = v$R3_7072_out0;
assign v$R3TEST_5095_out0 = v$R3_7073_out0;
assign v$END6_5096_out0 = v$LASTQ_7877_out0;
assign v$END6_5097_out0 = v$LASTQ_7888_out0;
assign v$G2_5108_out0 = ! v$OUTPUT_13145_out0;
assign v$G7_5374_out0 = ! v$Q3_12999_out0;
assign v$G7_5375_out0 = ! v$Q3_13000_out0;
assign v$DM1_5380_out0 = v$SELOUT_900_out0 ? 16'h0 : v$RAM1_8558_out0;
assign v$DM1_5380_out1 = v$SELOUT_900_out0 ? v$RAM1_8558_out0 : 16'h0;
assign v$RXDISABLE_5404_out0 = v$_3288_out1;
assign v$RXDISABLE_5405_out0 = v$_3289_out1;
assign v$G3_5549_out0 = v$FF1_178_out0 || v$G2_62_out0;
assign v$G3_5550_out0 = v$FF1_179_out0 || v$G2_63_out0;
assign v$END_5603_out0 = v$A1_2728_out1;
assign v$END_5604_out0 = v$A1_2729_out1;
assign v$_5609_out0 = { v$_525_out0,v$Q2_1883_out0 };
assign v$_5610_out0 = { v$_526_out0,v$Q2_1884_out0 };
assign v$END4_5637_out0 = v$LASTQ_7874_out0;
assign v$END4_5638_out0 = v$LASTQ_7885_out0;
assign v$R0TEST_5724_out0 = v$R0_1977_out0;
assign v$R0TEST_5725_out0 = v$R0_1978_out0;
assign v$LEFT$SHIFT_6043_out0 = v$LEFT$SHIFT_8476_out0;
assign v$LEFT$SHIFT_6044_out0 = v$LEFT$SHIFT_8477_out0;
assign v$LEFT$SHIFT_6045_out0 = v$LEFT$SHIFT_8478_out0;
assign v$LEFT$SHIFT_6046_out0 = v$LEFT$SHIFT_8479_out0;
assign v$LEFT$SHIFT_6047_out0 = v$LEFT$SHIFT_8480_out0;
assign v$LEFT$SHIFT_6048_out0 = v$LEFT$SHIFT_8481_out0;
assign v$LEFT$SHIFT_6049_out0 = v$LEFT$SHIFT_8482_out0;
assign v$LEFT$SHIFT_6050_out0 = v$LEFT$SHIFT_8483_out0;
assign v$_6223_out0 = v$B_12739_out0[7:0];
assign v$_6223_out1 = v$B_12739_out0[15:8];
assign v$_6224_out0 = v$B_12740_out0[7:0];
assign v$_6224_out1 = v$B_12740_out0[15:8];
assign v$G6_6314_out0 = ! v$Q2_3703_out0;
assign v$G6_6315_out0 = ! v$Q2_3704_out0;
assign v$MODE_6360_out0 = v$_3288_out0;
assign v$MODE_6361_out0 = v$_3289_out0;
assign v$A$SAVED_6682_out0 = v$A$SAVED_2413_out0;
assign v$A$SAVED_6683_out0 = v$A$SAVED_2414_out0;
assign v$G38_6823_out0 = v$Q0_13018_out0 || v$Q1_3089_out0;
assign v$G38_6824_out0 = v$Q0_13019_out0 || v$Q1_3090_out0;
assign v$INIT_7077_out0 = v$G2_62_out0;
assign v$INIT_7078_out0 = v$G2_63_out0;
assign v$_7112_out0 = v$_13131_out0[1:0];
assign v$_7112_out1 = v$_13131_out0[3:2];
assign v$_7113_out0 = v$_13132_out0[1:0];
assign v$_7113_out1 = v$_13132_out0[3:2];
assign v$I3P_7124_out0 = v$I3P_6221_out0;
assign v$I3P_7125_out0 = v$I3P_6222_out0;
assign v$CARRY_7187_out0 = v$CARRY_9008_out0;
assign v$CARRY_7188_out0 = v$CARRY_9009_out0;
assign v$TXLast_7426_out0 = v$LASTQ_7879_out0;
assign v$TXLast_7427_out0 = v$LASTQ_7890_out0;
assign v$G57_7492_out0 = ! v$HALT$PREV_6935_out0;
assign v$G57_7493_out0 = ! v$HALT$PREV_6936_out0;
assign v$G27_7526_out0 = v$Q0_9249_out0 && v$Q1_7197_out0;
assign v$G27_7527_out0 = v$Q0_9250_out0 && v$Q1_7198_out0;
assign v$_7616_out0 = v$_13131_out1[1:0];
assign v$_7616_out1 = v$_13131_out1[3:2];
assign v$_7617_out0 = v$_13132_out1[1:0];
assign v$_7617_out1 = v$_13132_out1[3:2];
assign v$HALTED_7627_out0 = v$OUTPUT_6891_out0;
assign v$HALTED_7628_out0 = v$OUTPUT_6892_out0;
assign v$INSTR$READ1_7747_out0 = v$OUT_3626_out0;
assign v$SEL8_8402_out0 = v$SAVED_10674_out0[11:0];
assign v$SEL8_8403_out0 = v$SAVED_10675_out0[11:0];
assign v$RXlast_8470_out0 = v$LASTQ_7880_out0;
assign v$RXlast_8471_out0 = v$LASTQ_7891_out0;
assign v$G6_8632_out0 = ((v$G2_529_out0 && !v$G3_11055_out0) || (!v$G2_529_out0) && v$G3_11055_out0);
assign v$G6_8633_out0 = ((v$G2_530_out0 && !v$G3_11056_out0) || (!v$G2_530_out0) && v$G3_11056_out0);
assign v$_8980_out0 = { v$Q2_12285_out0,v$Q3_13107_out0 };
assign v$_8981_out0 = { v$Q2_12286_out0,v$Q3_13108_out0 };
assign v$G7_9002_out0 = ((v$G4_1665_out0 && !v$G5_10022_out0) || (!v$G4_1665_out0) && v$G5_10022_out0);
assign v$G7_9003_out0 = ((v$G4_1666_out0 && !v$G5_10023_out0) || (!v$G4_1666_out0) && v$G5_10023_out0);
assign v$G86_9099_out0 = ! v$PHALT1_6182_out0;
assign v$EVENPARITY_9157_out0 = v$EPARITY_13014_out0;
assign v$EVENPARITY_9158_out0 = v$EPARITY_13015_out0;
assign v$G4_9398_out0 = ! v$Q0_9249_out0;
assign v$G4_9399_out0 = ! v$Q0_9250_out0;
assign v$G51_9413_out0 = ! v$HALT$PREV_6935_out0;
assign v$G51_9414_out0 = ! v$HALT$PREV_6936_out0;
assign v$G25_9422_out0 = ((v$Q0_13018_out0 && !v$Q1_3089_out0) || (!v$Q0_13018_out0) && v$Q1_3089_out0);
assign v$G25_9423_out0 = ((v$Q0_13019_out0 && !v$Q1_3090_out0) || (!v$Q0_13019_out0) && v$Q1_3090_out0);
assign v$INSTR$READ0_9560_out0 = v$OUT_3625_out0;
assign v$G7_9703_out0 = ! v$Q2_1883_out0;
assign v$G7_9704_out0 = ! v$Q2_1884_out0;
assign v$A$SAVED_10000_out0 = v$A$SAVED_2413_out0;
assign v$A$SAVED_10001_out0 = v$A$SAVED_2414_out0;
assign v$PHALT_10440_out0 = v$PHALT_834_out0;
assign v$R1TEST_10449_out0 = v$R1_9296_out0;
assign v$R1TEST_10450_out0 = v$R1_9297_out0;
assign v$R2TEST_10971_out0 = v$R2_5454_out0;
assign v$R2TEST_10972_out0 = v$R2_5455_out0;
assign v$G2_10999_out0 = ! v$Q1_3089_out0;
assign v$G2_11000_out0 = ! v$Q1_3090_out0;
assign v$G25_11283_out0 = ((v$G23_6381_out0 && !v$G24_12076_out0) || (!v$G23_6381_out0) && v$G24_12076_out0);
assign v$G25_11284_out0 = ((v$G23_6382_out0 && !v$G24_12077_out0) || (!v$G23_6382_out0) && v$G24_12077_out0);
assign v$_11296_out0 = { v$_2493_out0,v$_6431_out0 };
assign v$_11297_out0 = { v$_2494_out0,v$_6432_out0 };
assign v$G5_11318_out0 = ! v$Q1_7197_out0;
assign v$G5_11319_out0 = ! v$Q1_7198_out0;
v$AROM1_11322 I11322 (v$AROM1_11322_out0, v$ADDRESS_9958_out0);
v$AROM1_11323 I11323 (v$AROM1_11323_out0, v$ADDRESS_9959_out0);
assign v$G61_11531_out0 = ! v$HALT$PREV_6935_out0;
assign v$G61_11532_out0 = ! v$HALT$PREV_6936_out0;
assign v$G9_11572_out0 = ! v$Q0_74_out0;
assign v$G9_11573_out0 = ! v$Q0_75_out0;
assign v$PCHALT_11644_out0 = v$PCHALT_8399_out0;
assign v$CLK4_11784_out0 = v$G3_22_out0;
assign v$CLK4_11785_out0 = v$G3_23_out0;
assign v$END_12098_out0 = v$LASTQ_7881_out0;
assign v$END_12099_out0 = v$LASTQ_7892_out0;
assign v$G4_12393_out0 = ! v$Q3_13107_out0;
assign v$G4_12394_out0 = ! v$Q3_13108_out0;
assign v$increment_12632_out0 = v$EQ1_10629_out0;
assign v$increment_12633_out0 = v$EQ1_10630_out0;
assign v$G55_12935_out0 = ! v$HALT$PREV_6935_out0;
assign v$G55_12936_out0 = ! v$HALT$PREV_6936_out0;
assign v$_13026_out0 = { v$Q2_3703_out0,v$Q3_12999_out0 };
assign v$_13027_out0 = { v$Q2_3704_out0,v$Q3_13000_out0 };
assign v$G3_13101_out0 = ! v$Q2_12285_out0;
assign v$G3_13102_out0 = ! v$Q2_12286_out0;
assign v$G41_13147_out0 = v$Q0_13018_out0 && v$Q1_3089_out0;
assign v$G41_13148_out0 = v$Q0_13019_out0 && v$Q1_3090_out0;
assign v$_13175_out0 = { v$Q0_9249_out0,v$Q1_7197_out0 };
assign v$_13176_out0 = { v$Q0_9250_out0,v$Q1_7198_out0 };
assign v$NQ1_219_out0 = v$G5_11318_out0;
assign v$NQ1_220_out0 = v$G5_11319_out0;
assign v$SEL5_368_out0 = v$IR2_929_out0[11:10];
assign v$SEL5_369_out0 = v$IR2_930_out0[11:10];
assign v$G1_483_out0 = ! v$OFF_2756_out0;
assign v$G1_484_out0 = ! v$OFF_2757_out0;
assign v$NQ3_721_out0 = v$G7_5374_out0;
assign v$NQ3_722_out0 = v$G7_5375_out0;
assign v$MODE_821_out0 = v$MODE_6360_out0;
assign v$MODE_822_out0 = v$MODE_6361_out0;
assign v$IR2_1150_out0 = v$IR2_1700_out0;
assign v$IR2_1151_out0 = v$IR2_1701_out0;
assign v$_1279_out0 = v$_6223_out0[3:0];
assign v$_1279_out1 = v$_6223_out0[7:4];
assign v$_1280_out0 = v$_6224_out0[3:0];
assign v$_1280_out1 = v$_6224_out0[7:4];
assign v$G58_1431_out0 = v$FF11_1377_out0 && v$G57_7492_out0;
assign v$G58_1432_out0 = v$FF11_1378_out0 && v$G57_7493_out0;
assign v$_1673_out0 = v$_6223_out1[3:0];
assign v$_1673_out1 = v$_6223_out1[7:4];
assign v$_1674_out0 = v$_6224_out1[3:0];
assign v$_1674_out1 = v$_6224_out1[7:4];
assign v$NQ2_1741_out0 = v$G6_6314_out0;
assign v$NQ2_1742_out0 = v$G6_6315_out0;
assign v$NQ3_1759_out0 = v$G4_12393_out0;
assign v$NQ3_1760_out0 = v$G4_12394_out0;
assign v$LEFT$SHIT_1795_out0 = v$LEFT$SHIFT_6043_out0;
assign v$LEFT$SHIT_1796_out0 = v$LEFT$SHIFT_6043_out0;
assign v$LEFT$SHIT_1797_out0 = v$LEFT$SHIFT_6043_out0;
assign v$LEFT$SHIT_1798_out0 = v$LEFT$SHIFT_6043_out0;
assign v$LEFT$SHIT_1799_out0 = v$LEFT$SHIFT_6043_out0;
assign v$LEFT$SHIT_1812_out0 = v$LEFT$SHIFT_6044_out0;
assign v$LEFT$SHIT_1813_out0 = v$LEFT$SHIFT_6044_out0;
assign v$LEFT$SHIT_1814_out0 = v$LEFT$SHIFT_6044_out0;
assign v$LEFT$SHIT_1815_out0 = v$LEFT$SHIFT_6044_out0;
assign v$LEFT$SHIT_1816_out0 = v$LEFT$SHIFT_6044_out0;
assign v$LEFT$SHIT_1817_out0 = v$LEFT$SHIFT_6045_out0;
assign v$LEFT$SHIT_1818_out0 = v$LEFT$SHIFT_6045_out0;
assign v$LEFT$SHIT_1819_out0 = v$LEFT$SHIFT_6045_out0;
assign v$LEFT$SHIT_1820_out0 = v$LEFT$SHIFT_6045_out0;
assign v$LEFT$SHIT_1821_out0 = v$LEFT$SHIFT_6045_out0;
assign v$LEFT$SHIT_1822_out0 = v$LEFT$SHIFT_6046_out0;
assign v$LEFT$SHIT_1823_out0 = v$LEFT$SHIFT_6046_out0;
assign v$LEFT$SHIT_1824_out0 = v$LEFT$SHIFT_6046_out0;
assign v$LEFT$SHIT_1825_out0 = v$LEFT$SHIFT_6046_out0;
assign v$LEFT$SHIT_1826_out0 = v$LEFT$SHIFT_6046_out0;
assign v$LEFT$SHIT_1827_out0 = v$LEFT$SHIFT_6047_out0;
assign v$LEFT$SHIT_1828_out0 = v$LEFT$SHIFT_6047_out0;
assign v$LEFT$SHIT_1829_out0 = v$LEFT$SHIFT_6047_out0;
assign v$LEFT$SHIT_1830_out0 = v$LEFT$SHIFT_6047_out0;
assign v$LEFT$SHIT_1831_out0 = v$LEFT$SHIFT_6047_out0;
assign v$LEFT$SHIT_1844_out0 = v$LEFT$SHIFT_6048_out0;
assign v$LEFT$SHIT_1845_out0 = v$LEFT$SHIFT_6048_out0;
assign v$LEFT$SHIT_1846_out0 = v$LEFT$SHIFT_6048_out0;
assign v$LEFT$SHIT_1847_out0 = v$LEFT$SHIFT_6048_out0;
assign v$LEFT$SHIT_1848_out0 = v$LEFT$SHIFT_6048_out0;
assign v$LEFT$SHIT_1849_out0 = v$LEFT$SHIFT_6049_out0;
assign v$LEFT$SHIT_1850_out0 = v$LEFT$SHIFT_6049_out0;
assign v$LEFT$SHIT_1851_out0 = v$LEFT$SHIFT_6049_out0;
assign v$LEFT$SHIT_1852_out0 = v$LEFT$SHIFT_6049_out0;
assign v$LEFT$SHIT_1853_out0 = v$LEFT$SHIFT_6049_out0;
assign v$LEFT$SHIT_1854_out0 = v$LEFT$SHIFT_6050_out0;
assign v$LEFT$SHIT_1855_out0 = v$LEFT$SHIFT_6050_out0;
assign v$LEFT$SHIT_1856_out0 = v$LEFT$SHIFT_6050_out0;
assign v$LEFT$SHIT_1857_out0 = v$LEFT$SHIFT_6050_out0;
assign v$LEFT$SHIT_1858_out0 = v$LEFT$SHIFT_6050_out0;
assign v$_1864_out0 = v$_7616_out1[0:0];
assign v$_1864_out1 = v$_7616_out1[1:1];
assign v$_1865_out0 = v$_7617_out1[0:0];
assign v$_1865_out1 = v$_7617_out1[1:1];
assign v$_2400_out0 = v$_7112_out1[0:0];
assign v$_2400_out1 = v$_7112_out1[1:1];
assign v$_2401_out0 = v$_7113_out1[0:0];
assign v$_2401_out1 = v$_7113_out1[1:1];
assign v$SEL13_3246_out0 = v$IR2_929_out0[9:8];
assign v$SEL13_3247_out0 = v$IR2_930_out0[9:8];
assign v$CARRY_3395_out0 = v$CARRY_7187_out0;
assign v$CARRY_3396_out0 = v$CARRY_7188_out0;
assign v$_3451_out0 = v$_7616_out0[0:0];
assign v$_3451_out1 = v$_7616_out0[1:1];
assign v$_3452_out0 = v$_7617_out0[0:0];
assign v$_3452_out1 = v$_7617_out0[1:1];
assign v$_4458_out0 = v$_749_out1[3:0];
assign v$_4458_out1 = v$_749_out1[7:4];
assign v$_4459_out0 = v$_750_out1[3:0];
assign v$_4459_out1 = v$_750_out1[7:4];
assign v$_4743_out0 = v$_7112_out0[0:0];
assign v$_4743_out1 = v$_7112_out0[1:1];
assign v$_4744_out0 = v$_7113_out0[0:0];
assign v$_4744_out1 = v$_7113_out0[1:1];
assign v$EDGE2_4761_out0 = v$INTERRUPT2_2562_out0;
assign v$EDGE2_4762_out0 = v$INTERRUPT2_2563_out0;
assign v$SEL4_4802_out0 = v$IR2_929_out0[15:15];
assign v$SEL4_4803_out0 = v$IR2_930_out0[15:15];
assign v$CLK4_4804_out0 = v$CLK4_11784_out0;
assign v$CLK4_4805_out0 = v$CLK4_11785_out0;
assign v$INSTR$READ_4830_out0 = v$INSTR$READ0_9560_out0;
assign v$INSTR$READ_4831_out0 = v$INSTR$READ1_7747_out0;
assign v$SEL10_4877_out0 = v$IR2_929_out0[9:9];
assign v$SEL10_4878_out0 = v$IR2_930_out0[9:9];
assign v$NQ0_5322_out0 = v$G4_9398_out0;
assign v$NQ0_5323_out0 = v$G4_9399_out0;
assign v$RAMDOUT1_5788_out0 = v$DM1_5380_out1;
assign v$SEL11_5832_out0 = v$IR2_929_out0[8:8];
assign v$SEL11_5833_out0 = v$IR2_930_out0[8:8];
assign v$_5874_out0 = v$_749_out0[3:0];
assign v$_5874_out1 = v$_749_out0[7:4];
assign v$_5875_out0 = v$_750_out0[3:0];
assign v$_5875_out1 = v$_750_out0[7:4];
assign v$G65_6054_out0 = ! v$PHALT_10440_out0;
assign v$_6183_out0 = { v$_13175_out0,v$_13026_out0 };
assign v$_6184_out0 = { v$_13176_out0,v$_13027_out0 };
assign v$RAMDOUT0_6338_out0 = v$DM1_5380_out0;
assign v$G3_6429_out0 = ! v$RXDISABLE_5404_out0;
assign v$G3_6430_out0 = ! v$RXDISABLE_5405_out0;
assign v$_6656_out0 = v$AROM1_11322_out0[27:0];
assign v$_6656_out1 = v$AROM1_11322_out0[43:16];
assign v$_6657_out0 = v$AROM1_11323_out0[27:0];
assign v$_6657_out1 = v$AROM1_11323_out0[43:16];
assign v$_6821_out0 = { v$_1005_out0,v$_8980_out0 };
assign v$_6822_out0 = { v$_1006_out0,v$_8981_out0 };
assign v$Mode_7235_out0 = v$MODE_6360_out0;
assign v$Mode_7236_out0 = v$MODE_6361_out0;
assign v$G3_7242_out0 = ! v$OFF_2756_out0;
assign v$G3_7243_out0 = ! v$OFF_2757_out0;
assign v$NQ1_7276_out0 = v$G2_10999_out0;
assign v$NQ1_7277_out0 = v$G2_11000_out0;
assign v$G8_8068_out0 = ((v$G6_8632_out0 && !v$G7_9002_out0) || (!v$G6_8632_out0) && v$G7_9002_out0);
assign v$G8_8069_out0 = ((v$G6_8633_out0 && !v$G7_9003_out0) || (!v$G6_8633_out0) && v$G7_9003_out0);
assign v$SEL12_8456_out0 = v$IR2_929_out0[15:12];
assign v$SEL12_8457_out0 = v$IR2_930_out0[15:12];
assign v$Mode_8796_out0 = v$MODE_6360_out0;
assign v$Mode_8797_out0 = v$MODE_6361_out0;
assign v$EQ1_8927_out0 = v$_5609_out0 == 3'h0;
assign v$EQ1_8928_out0 = v$_5610_out0 == 3'h0;
assign v$G67_9285_out0 = ! v$PHALT_10440_out0;
assign v$G70_9421_out0 = v$PCHALT_11644_out0 && v$PHALT_10440_out0;
assign v$G67_9496_out0 = v$HALTED_7627_out0 && v$VALID$PREV_9000_out0;
assign v$G67_9497_out0 = v$HALTED_7628_out0 && v$VALID$PREV_9001_out0;
assign v$G4_9611_out0 = v$SOUT1_1070_out0 || v$INIT_7077_out0;
assign v$G4_9612_out0 = v$SOUT1_1076_out0 || v$INIT_7078_out0;
assign v$_10020_out0 = { v$_3718_out0,v$_4782_out0 };
assign v$_10021_out0 = { v$_3719_out0,v$_4783_out0 };
assign v$HALTSEL_10098_out0 = v$G2_5108_out0;
assign v$NQ0_10672_out0 = v$G9_11572_out0;
assign v$NQ0_10673_out0 = v$G9_11573_out0;
assign v$NQ0_10890_out0 = v$G1_794_out0;
assign v$NQ0_10891_out0 = v$G1_795_out0;
assign v$_10934_out0 = { v$_3760_out0,v$_11296_out0 };
assign v$_10935_out0 = { v$_3761_out0,v$_11297_out0 };
assign v$G69_11035_out0 = v$PCHALT_11644_out0 && v$PHALT_10440_out0;
assign v$G26_11199_out0 = ((v$G25_11283_out0 && !v$G22_4865_out0) || (!v$G25_11283_out0) && v$G22_4865_out0);
assign v$G26_11200_out0 = ((v$G25_11284_out0 && !v$G22_4866_out0) || (!v$G25_11284_out0) && v$G22_4866_out0);
assign v$NQ2_11764_out0 = v$G7_9703_out0;
assign v$NQ2_11765_out0 = v$G7_9704_out0;
assign v$NQ1_11780_out0 = v$G8_1189_out0;
assign v$NQ1_11781_out0 = v$G8_1190_out0;
assign v$CIN_11850_out0 = v$CIN_2595_out0;
assign v$CIN_11862_out0 = v$CIN_2607_out0;
assign v$PHALT_12284_out0 = v$G2_5108_out0;
assign v$CLEAR_13091_out0 = v$G1_30_out0;
assign v$CLEAR_13092_out0 = v$G1_31_out0;
assign v$RceivedParity_13191_out0 = v$RECIEVEDPARITY_4231_out0;
assign v$RceivedParity_13192_out0 = v$RECIEVEDPARITY_4232_out0;
assign v$NQ2_13211_out0 = v$G3_13101_out0;
assign v$NQ2_13212_out0 = v$G3_13102_out0;
assign v$PIPELINE$RESTART_13261_out0 = v$PIPELINE$RESTART_4073_out0;
assign v$PIPELINE$RESTART_13262_out0 = v$PIPELINE$RESTART_4074_out0;
assign v$_192_out0 = v$_5874_out1[1:0];
assign v$_192_out1 = v$_5874_out1[3:2];
assign v$_193_out0 = v$_5875_out1[1:0];
assign v$_193_out1 = v$_5875_out1[3:2];
assign v$G43_319_out0 = v$NQ2_13211_out0 && v$Q3_13107_out0;
assign v$G43_320_out0 = v$NQ2_13212_out0 && v$Q3_13108_out0;
assign v$G37_394_out0 = v$NQ0_5322_out0 || v$NQ1_219_out0;
assign v$G37_395_out0 = v$NQ0_5323_out0 || v$NQ1_220_out0;
assign v$S_495_out0 = v$PHALT_12284_out0;
assign v$RXCLK_507_out0 = v$EQ1_8927_out0;
assign v$RXCLK_508_out0 = v$EQ1_8928_out0;
assign v$EQ12_761_out0 = v$SEL12_8456_out0 == 4'h0;
assign v$EQ12_762_out0 = v$SEL12_8457_out0 == 4'h0;
assign v$_807_out0 = v$_4458_out1[1:0];
assign v$_807_out1 = v$_4458_out1[3:2];
assign v$_808_out0 = v$_4459_out1[1:0];
assign v$_808_out1 = v$_4459_out1[3:2];
assign v$INTERRUPT2_857_out0 = v$EDGE2_4761_out0;
assign v$INTERRUPT2_858_out0 = v$EDGE2_4762_out0;
assign v$_865_out0 = v$_6656_out1[7:0];
assign v$_865_out1 = v$_6656_out1[15:8];
assign v$_866_out0 = v$_6657_out1[7:0];
assign v$_866_out1 = v$_6657_out1[15:8];
assign v$G54_1052_out0 = v$NQ1_219_out0 && v$NQ0_5322_out0;
assign v$G54_1053_out0 = v$NQ1_220_out0 && v$NQ0_5323_out0;
assign v$G23_1199_out0 = v$NQ3_721_out0 || v$NQ2_1741_out0;
assign v$G23_1200_out0 = v$NQ3_722_out0 || v$NQ2_1742_out0;
assign v$_1213_out0 = v$_1279_out0[1:0];
assign v$_1213_out1 = v$_1279_out0[3:2];
assign v$_1214_out0 = v$_1280_out0[1:0];
assign v$_1214_out1 = v$_1280_out0[3:2];
assign v$G19_1347_out0 = v$NQ1_219_out0 && v$NQ2_1741_out0;
assign v$G19_1348_out0 = v$NQ1_220_out0 && v$NQ2_1742_out0;
assign v$G51_1633_out0 = v$Q3_12999_out0 && v$NQ2_1741_out0;
assign v$G51_1634_out0 = v$Q3_13000_out0 && v$NQ2_1742_out0;
assign v$G16_1783_out0 = v$NQ1_11780_out0 && v$Q2_1883_out0;
assign v$G16_1784_out0 = v$NQ1_11781_out0 && v$Q2_1884_out0;
assign v$G56_1877_out0 = v$NQ3_721_out0 && v$Q0_9249_out0;
assign v$G56_1878_out0 = v$NQ3_722_out0 && v$Q0_9250_out0;
assign v$Write_1959_out0 = v$CLEAR_13091_out0;
assign v$Write_1960_out0 = v$CLEAR_13091_out0;
assign v$Write_1961_out0 = v$CLEAR_13091_out0;
assign v$Write_1962_out0 = v$CLEAR_13091_out0;
assign v$Write_1963_out0 = v$CLEAR_13091_out0;
assign v$Write_1964_out0 = v$CLEAR_13091_out0;
assign v$Write_1965_out0 = v$CLEAR_13092_out0;
assign v$Write_1966_out0 = v$CLEAR_13092_out0;
assign v$Write_1967_out0 = v$CLEAR_13092_out0;
assign v$Write_1968_out0 = v$CLEAR_13092_out0;
assign v$Write_1969_out0 = v$CLEAR_13092_out0;
assign v$Write_1970_out0 = v$CLEAR_13092_out0;
assign v$F1_2195_out0 = v$_3451_out1;
assign v$F1_2196_out0 = v$_3452_out1;
assign v$C_2344_out0 = v$CARRY_3395_out0;
assign v$C_2345_out0 = v$CARRY_3396_out0;
assign v$CLK4_2409_out0 = v$CLK4_4804_out0;
assign v$CLK4_2410_out0 = v$CLK4_4805_out0;
assign v$RXENABLE_2429_out0 = v$G3_6429_out0;
assign v$RXENABLE_2430_out0 = v$G3_6430_out0;
assign v$G59_2552_out0 = v$Q2_12285_out0 && v$NQ3_1759_out0;
assign v$G59_2553_out0 = v$Q2_12286_out0 && v$NQ3_1760_out0;
assign v$R2_2554_out0 = v$_2400_out0;
assign v$R2_2555_out0 = v$_2401_out0;
assign v$IR2_2660_out0 = v$IR2_1150_out0;
assign v$IR2_2661_out0 = v$IR2_1151_out0;
assign v$G26_2796_out0 = v$G27_7526_out0 && v$NQ2_1741_out0;
assign v$G26_2797_out0 = v$G27_7527_out0 && v$NQ2_1742_out0;
assign v$G15_2890_out0 = v$NQ0_10890_out0 && v$Q1_3089_out0;
assign v$G15_2891_out0 = v$NQ0_10891_out0 && v$Q1_3090_out0;
assign v$G11_3264_out0 = v$NQ2_1741_out0 && v$NQ1_219_out0;
assign v$G11_3265_out0 = v$NQ2_1742_out0 && v$NQ1_220_out0;
assign v$_3516_out0 = v$_1279_out1[1:0];
assign v$_3516_out1 = v$_1279_out1[3:2];
assign v$_3517_out0 = v$_1280_out1[1:0];
assign v$_3517_out1 = v$_1280_out1[3:2];
assign v$EQ13_3617_out0 = v$SEL12_8456_out0 == 4'h1;
assign v$EQ13_3618_out0 = v$SEL12_8457_out0 == 4'h1;
assign v$_4077_out0 = v$Mode_7235_out0[0:0];
assign v$_4077_out1 = v$Mode_7235_out0[2:2];
assign v$_4078_out0 = v$Mode_7236_out0[0:0];
assign v$_4078_out1 = v$Mode_7236_out0[2:2];
assign v$Q_4167_out0 = v$_6821_out0;
assign v$Q_4168_out0 = v$_6822_out0;
assign v$IR2$REG$IMMEDIATE_4213_out0 = v$SEL10_4877_out0;
assign v$IR2$REG$IMMEDIATE_4214_out0 = v$SEL10_4878_out0;
assign v$G16_4419_out0 = v$NQ3_721_out0 && v$Q2_3703_out0;
assign v$G16_4420_out0 = v$NQ3_722_out0 && v$Q2_3704_out0;
assign v$_4973_out0 = v$_1673_out0[1:0];
assign v$_4973_out1 = v$_1673_out0[3:2];
assign v$_4974_out0 = v$_1674_out0[1:0];
assign v$_4974_out1 = v$_1674_out0[3:2];
assign v$G29_5042_out0 = v$NQ1_219_out0 || v$NQ0_5322_out0;
assign v$G29_5043_out0 = v$NQ1_220_out0 || v$NQ0_5323_out0;
assign v$IR2$FPU$OP_5098_out0 = v$SEL13_3246_out0;
assign v$IR2$FPU$OP_5099_out0 = v$SEL13_3247_out0;
assign v$_5700_out0 = v$_5874_out0[1:0];
assign v$_5700_out1 = v$_5874_out0[3:2];
assign v$_5701_out0 = v$_5875_out0[1:0];
assign v$_5701_out1 = v$_5875_out0[3:2];
assign v$G11_5718_out0 = v$NQ1_11780_out0 && v$NQ0_10672_out0;
assign v$G11_5719_out0 = v$NQ1_11781_out0 && v$NQ0_10673_out0;
assign v$F3_5730_out0 = v$_1864_out1;
assign v$F3_5731_out0 = v$_1865_out1;
assign v$G66_6177_out0 = v$PCHALT_11644_out0 && v$G65_6054_out0;
assign v$G32_6353_out0 = v$NQ1_7276_out0 || v$NQ0_10890_out0;
assign v$G32_6354_out0 = v$NQ1_7277_out0 || v$NQ0_10891_out0;
assign v$_6415_out0 = v$_1673_out1[1:0];
assign v$_6415_out1 = v$_1673_out1[3:2];
assign v$_6416_out0 = v$_1674_out1[1:0];
assign v$_6416_out1 = v$_1674_out1[3:2];
assign v$G42_6544_out0 = v$Q2_12285_out0 && v$NQ3_1759_out0;
assign v$G42_6545_out0 = v$Q2_12286_out0 && v$NQ3_1760_out0;
assign v$MUX1_6647_out0 = v$CLEAR_13091_out0 ? v$C3_8772_out0 : v$A1_2728_out0;
assign v$MUX1_6648_out0 = v$CLEAR_13092_out0 ? v$C3_8773_out0 : v$A1_2729_out0;
assign v$IS$IR2$DATA$PROCESSING_6664_out0 = v$SEL4_4802_out0;
assign v$IS$IR2$DATA$PROCESSING_6665_out0 = v$SEL4_4803_out0;
assign v$G49_6992_out0 = v$NQ3_721_out0 && v$Q1_7197_out0;
assign v$G49_6993_out0 = v$NQ3_722_out0 && v$Q1_7198_out0;
assign v$G5_7012_out0 = v$NQ2_11764_out0 && v$G6_2050_out0;
assign v$G5_7013_out0 = v$NQ2_11765_out0 && v$G6_2051_out0;
assign v$G36_7154_out0 = v$NQ2_1741_out0 && v$Q3_12999_out0;
assign v$G36_7155_out0 = v$NQ2_1742_out0 && v$Q3_13000_out0;
assign v$G17_7508_out0 = v$NQ2_1741_out0 && v$Q1_7197_out0;
assign v$G17_7509_out0 = v$NQ2_1742_out0 && v$Q1_7198_out0;
assign v$F2_7871_out0 = v$_1864_out0;
assign v$F2_7872_out0 = v$_1865_out0;
assign v$DATA$OUT0_8072_out0 = v$RAMDOUT0_6338_out0;
assign v$Q_8619_out0 = v$_6183_out0;
assign v$Q_8620_out0 = v$_6184_out0;
assign v$G50_8804_out0 = v$NQ3_721_out0 && v$Q2_3703_out0;
assign v$G50_8805_out0 = v$NQ3_722_out0 && v$Q2_3704_out0;
assign v$_8866_out0 = v$_4458_out0[1:0];
assign v$_8866_out1 = v$_4458_out0[3:2];
assign v$_8867_out0 = v$_4459_out0[1:0];
assign v$_8867_out1 = v$_4459_out0[3:2];
assign v$_8872_out0 = v$Mode_8796_out0[0:0];
assign v$_8872_out1 = v$Mode_8796_out0[2:2];
assign v$_8873_out0 = v$Mode_8797_out0[0:0];
assign v$_8873_out1 = v$Mode_8797_out0[2:2];
assign v$G9_9012_out0 = v$NQ2_13211_out0 && v$NQ1_7276_out0;
assign v$G9_9013_out0 = v$NQ2_13212_out0 && v$NQ1_7277_out0;
assign v$MUX6_9127_out0 = v$PIPELINE$RESTART_13261_out0 ? v$C2_9087_out0 : v$FF9_6996_out0;
assign v$MUX6_9128_out0 = v$PIPELINE$RESTART_13262_out0 ? v$C2_9088_out0 : v$FF9_6997_out0;
assign v$POut_9234_out0 = v$_10934_out0;
assign v$POut_9235_out0 = v$_10935_out0;
assign v$G68_10170_out0 = v$PCHALT_11644_out0 && v$G67_9285_out0;
assign v$INSTR$READ_10224_out0 = v$INSTR$READ_4830_out0;
assign v$INSTR$READ_10225_out0 = v$INSTR$READ_4831_out0;
assign v$G62_10313_out0 = v$Q3_13107_out0 && v$NQ2_13211_out0;
assign v$G62_10314_out0 = v$Q3_13108_out0 && v$NQ2_13212_out0;
assign v$R1_10327_out0 = v$_4743_out1;
assign v$R1_10328_out0 = v$_4744_out1;
assign v$R0_10497_out0 = v$_4743_out0;
assign v$R0_10498_out0 = v$_4744_out0;
assign v$R3_10621_out0 = v$_2400_out1;
assign v$R3_10622_out0 = v$_2401_out1;
assign v$DATA$OUT1_10871_out0 = v$RAMDOUT1_5788_out0;
assign v$F0_11052_out0 = v$_3451_out0;
assign v$F0_11053_out0 = v$_3452_out0;
assign v$G3_11270_out0 = ! v$PHALT_12284_out0;
assign v$IR2$RD_11468_out0 = v$SEL5_368_out0;
assign v$IR2$RD_11469_out0 = v$SEL5_369_out0;
assign v$_11477_out0 = v$_6656_out0[11:0];
assign v$_11477_out1 = v$_6656_out0[27:16];
assign v$_11478_out0 = v$_6657_out0[11:0];
assign v$_11478_out1 = v$_6657_out0[27:16];
assign v$G50_12147_out0 = v$Q2_12285_out0 && v$NQ3_1759_out0;
assign v$G50_12148_out0 = v$Q2_12286_out0 && v$NQ3_1760_out0;
assign v$IR2$S$WB_12240_out0 = v$SEL11_5832_out0;
assign v$IR2$S$WB_12241_out0 = v$SEL11_5833_out0;
assign v$_12276_out0 = { v$G1_483_out0,v$C2_12781_out0 };
assign v$_12277_out0 = { v$G1_484_out0,v$C2_12782_out0 };
assign v$CLK4_12743_out0 = v$CLK4_4804_out0;
assign v$CLK4_12744_out0 = v$CLK4_4805_out0;
assign v$G68_12849_out0 = v$HALT$PREV$PREV_12829_out0 || v$G67_9496_out0;
assign v$G68_12850_out0 = v$HALT$PREV$PREV_12830_out0 || v$G67_9497_out0;
assign v$TX_12978_out0 = v$G4_9611_out0;
assign v$TX_12979_out0 = v$G4_9612_out0;
assign v$_13007_out0 = v$MODE_821_out0[0:0];
assign v$_13007_out1 = v$MODE_821_out0[2:2];
assign v$_13008_out0 = v$MODE_822_out0[0:0];
assign v$_13008_out1 = v$MODE_822_out0[2:2];
assign v$G14_13117_out0 = v$NQ0_10672_out0 && v$NQ2_11764_out0;
assign v$G14_13118_out0 = v$NQ0_10673_out0 && v$NQ2_11765_out0;
assign v$G42_13143_out0 = v$Q0_9249_out0 && v$NQ3_721_out0;
assign v$G42_13144_out0 = v$Q0_9250_out0 && v$NQ3_722_out0;
assign v$G60_13385_out0 = v$NQ3_1759_out0 && v$Q1_3089_out0;
assign v$G60_13386_out0 = v$NQ3_1760_out0 && v$Q1_3090_out0;
assign v$R_56_out0 = v$INSTR$READ_10224_out0;
assign v$R_57_out0 = v$INSTR$READ_10225_out0;
assign v$EQ7_201_out0 = v$Q_4167_out0 == 4'hc;
assign v$EQ7_202_out0 = v$Q_4168_out0 == 4'hc;
assign v$END_317_out0 = v$_8872_out1;
assign v$END_318_out0 = v$_8873_out1;
assign v$8_481_out0 = v$IR2_2660_out0[11:10];
assign v$8_482_out0 = v$IR2_2661_out0[11:10];
assign v$SEL12_581_out0 = v$IR2_2660_out0[6:6];
assign v$SEL12_582_out0 = v$IR2_2661_out0[6:6];
assign v$EQ6_773_out0 = v$Q_4167_out0 == 4'hb;
assign v$EQ6_774_out0 = v$Q_4168_out0 == 4'hb;
assign v$6_1094_out0 = v$IR2_2660_out0[15:15];
assign v$6_1095_out0 = v$IR2_2661_out0[15:15];
assign v$G48_1203_out0 = v$G51_1633_out0 && v$G54_1052_out0;
assign v$G48_1204_out0 = v$G51_1634_out0 && v$G54_1053_out0;
assign v$EQ3_1515_out0 = v$Q_4167_out0 == 4'hb;
assign v$EQ3_1516_out0 = v$Q_4168_out0 == 4'hb;
assign v$EQ4_1519_out0 = v$Q_8619_out0 == 4'h9;
assign v$EQ4_1520_out0 = v$Q_8620_out0 == 4'h9;
assign v$IR2_1985_out0 = v$IR2_2660_out0;
assign v$IR2_1986_out0 = v$IR2_2661_out0;
assign v$_2495_out0 = v$_4973_out0[0:0];
assign v$_2495_out1 = v$_4973_out0[1:1];
assign v$_2496_out0 = v$_4974_out0[0:0];
assign v$_2496_out1 = v$_4974_out0[1:1];
assign v$_2714_out0 = v$_4077_out1[0:0];
assign v$_2714_out1 = v$_4077_out1[1:1];
assign v$_2715_out0 = v$_4078_out1[0:0];
assign v$_2715_out1 = v$_4078_out1[1:1];
assign v$_2732_out0 = v$_5700_out0[0:0];
assign v$_2732_out1 = v$_5700_out0[1:1];
assign v$_2733_out0 = v$_5701_out0[0:0];
assign v$_2733_out1 = v$_5701_out0[1:1];
assign v$SEL10_2841_out0 = v$IR2_2660_out0[5:5];
assign v$SEL10_2842_out0 = v$IR2_2661_out0[5:5];
assign v$EQ3_2888_out0 = v$Q_8619_out0 == 4'hb;
assign v$EQ3_2889_out0 = v$Q_8620_out0 == 4'hb;
assign v$IR2$IS$LDST_3050_out0 = v$EQ12_761_out0;
assign v$IR2$IS$LDST_3051_out0 = v$EQ12_762_out0;
assign v$_3183_out0 = v$_192_out1[0:0];
assign v$_3183_out1 = v$_192_out1[1:1];
assign v$_3184_out0 = v$_193_out1[0:0];
assign v$_3184_out1 = v$_193_out1[1:1];
assign v$G47_3665_out0 = v$G49_6992_out0 || v$G50_8804_out0;
assign v$G47_3666_out0 = v$G49_6993_out0 || v$G50_8805_out0;
assign v$EQ14_3730_out0 = v$IR2$FPU$OP_5098_out0 == 2'h3;
assign v$EQ14_3731_out0 = v$IR2$FPU$OP_5099_out0 == 2'h3;
assign v$_3805_out0 = v$_192_out0[0:0];
assign v$_3805_out1 = v$_192_out0[1:1];
assign v$_3806_out0 = v$_193_out0[0:0];
assign v$_3806_out1 = v$_193_out0[1:1];
assign v$RX_4204_out0 = v$TX_12978_out0;
assign v$RX_4205_out0 = v$TX_12979_out0;
assign v$PIN_4636_out0 = v$_865_out1;
assign v$PIN_4639_out0 = v$_865_out0;
assign v$PIN_4642_out0 = v$_866_out1;
assign v$PIN_4645_out0 = v$_866_out0;
assign v$G21_4790_out0 = ! v$INTERRUPT2_857_out0;
assign v$G21_4791_out0 = ! v$INTERRUPT2_858_out0;
assign v$G58_4796_out0 = v$G60_13385_out0 || v$G59_2552_out0;
assign v$G58_4797_out0 = v$G60_13386_out0 || v$G59_2553_out0;
assign v$IR2$IS$FPU_4798_out0 = v$EQ13_3617_out0;
assign v$IR2$IS$FPU_4799_out0 = v$EQ13_3618_out0;
assign v$_4885_out0 = v$_8866_out1[0:0];
assign v$_4885_out1 = v$_8866_out1[1:1];
assign v$_4886_out0 = v$_8867_out1[0:0];
assign v$_4886_out1 = v$_8867_out1[1:1];
assign v$EQ1_5014_out0 = v$Q_4167_out0 == 4'h9;
assign v$EQ1_5015_out0 = v$Q_4168_out0 == 4'h9;
assign v$5_5074_out0 = v$IR2_2660_out0[1:0];
assign v$5_5075_out0 = v$IR2_2661_out0[1:0];
assign v$STP$SAVED_5106_out0 = v$MUX6_9127_out0;
assign v$STP$SAVED_5107_out0 = v$MUX6_9128_out0;
assign v$DATA$OUT_5146_out0 = v$DATA$OUT0_8072_out0;
assign v$DATA$OUT_5147_out0 = v$DATA$OUT1_10871_out0;
assign v$_5488_out0 = v$_1213_out1[0:0];
assign v$_5488_out1 = v$_1213_out1[1:1];
assign v$_5489_out0 = v$_1214_out1[0:0];
assign v$_5489_out1 = v$_1214_out1[1:1];
assign v$S_5524_out0 = v$S_495_out0;
assign v$G61_5755_out0 = v$G62_10313_out0 && v$NQ1_7276_out0;
assign v$G61_5756_out0 = v$G62_10314_out0 && v$NQ1_7277_out0;
assign v$P_5784_out0 = v$_8872_out0;
assign v$P_5785_out0 = v$_8873_out0;
assign v$_6017_out0 = v$_807_out0[0:0];
assign v$_6017_out1 = v$_807_out0[1:1];
assign v$_6018_out0 = v$_808_out0[0:0];
assign v$_6018_out1 = v$_808_out0[1:1];
assign v$_6057_out0 = v$_3516_out1[0:0];
assign v$_6057_out1 = v$_3516_out1[1:1];
assign v$_6058_out0 = v$_3517_out1[0:0];
assign v$_6058_out1 = v$_3517_out1[1:1];
assign v$EQ5_6345_out0 = v$Q_4167_out0 == 4'ha;
assign v$EQ5_6346_out0 = v$Q_4168_out0 == 4'ha;
assign v$SEL4_6439_out0 = v$IR2_2660_out0[9:8];
assign v$SEL4_6440_out0 = v$IR2_2661_out0[9:8];
assign v$G60_6463_out0 = v$G61_11531_out0 && v$G68_12849_out0;
assign v$G60_6464_out0 = v$G61_11532_out0 && v$G68_12850_out0;
assign v$_6473_out0 = v$_6415_out0[0:0];
assign v$_6473_out1 = v$_6415_out0[1:1];
assign v$_6474_out0 = v$_6416_out0[0:0];
assign v$_6474_out1 = v$_6416_out0[1:1];
assign v$EQ4_6581_out0 = v$Q_4167_out0 == 4'hc;
assign v$EQ4_6582_out0 = v$Q_4168_out0 == 4'hc;
assign v$RXBYTE_6584_out0 = v$POut_9234_out0;
assign v$RXBYTE_6585_out0 = v$POut_9235_out0;
assign v$EQ2_7440_out0 = v$Q_8619_out0 == 4'ha;
assign v$EQ2_7441_out0 = v$Q_8620_out0 == 4'ha;
assign v$G28_7730_out0 = v$Q2_3703_out0 && v$G29_5042_out0;
assign v$G28_7731_out0 = v$Q2_3704_out0 && v$G29_5043_out0;
assign v$PARITY_7858_out0 = v$_13007_out0;
assign v$PARITY_7859_out0 = v$_13008_out0;
assign v$_7862_out0 = v$_5700_out1[0:0];
assign v$_7862_out1 = v$_5700_out1[1:1];
assign v$_7863_out0 = v$_5701_out1[0:0];
assign v$_7863_out1 = v$_5701_out1[1:1];
assign v$G35_8276_out0 = v$G36_7154_out0 && v$G37_394_out0;
assign v$G35_8277_out0 = v$G36_7155_out0 && v$G37_395_out0;
assign v$_8546_out0 = v$_11477_out0[3:0];
assign v$_8546_out1 = v$_11477_out0[11:8];
assign v$_8547_out0 = v$_11478_out0[3:0];
assign v$_8547_out1 = v$_11478_out0[11:8];
assign v$G40_9224_out0 = v$G41_13147_out0 && v$G42_6544_out0;
assign v$G40_9225_out0 = v$G41_13148_out0 && v$G42_6545_out0;
assign {v$A1_9247_out1,v$A1_9247_out0 } = v$REG1_9161_out0 + v$_12276_out0 + v$C1_4454_out0;
assign {v$A1_9248_out1,v$A1_9248_out0 } = v$REG1_9162_out0 + v$_12277_out0 + v$C1_4455_out0;
assign v$_9360_out0 = v$_4973_out1[0:0];
assign v$_9360_out1 = v$_4973_out1[1:1];
assign v$_9361_out0 = v$_4974_out1[0:0];
assign v$_9361_out1 = v$_4974_out1[1:1];
assign v$9_9550_out0 = v$IR2_2660_out0[14:12];
assign v$9_9551_out0 = v$IR2_2661_out0[14:12];
assign v$_9644_out0 = v$_807_out1[0:0];
assign v$_9644_out1 = v$_807_out1[1:1];
assign v$_9645_out0 = v$_808_out1[0:0];
assign v$_9645_out1 = v$_808_out1[1:1];
assign v$EQ1_9709_out0 = v$Q_8619_out0 == 4'h1;
assign v$EQ1_9710_out0 = v$Q_8620_out0 == 4'h1;
assign v$_9897_out0 = v$_1213_out0[0:0];
assign v$_9897_out1 = v$_1213_out0[1:1];
assign v$_9898_out0 = v$_1214_out0[0:0];
assign v$_9898_out1 = v$_1214_out0[1:1];
assign v$G25_9956_out0 = v$INTERRUPT2_857_out0 && v$G24_7868_out0;
assign v$G25_9957_out0 = v$INTERRUPT2_858_out0 && v$G24_7869_out0;
assign v$G2_10344_out0 = ! v$Write_1959_out0;
assign v$G2_10345_out0 = ! v$Write_1960_out0;
assign v$G2_10346_out0 = ! v$Write_1961_out0;
assign v$G2_10347_out0 = ! v$Write_1962_out0;
assign v$G2_10348_out0 = ! v$Write_1963_out0;
assign v$G2_10349_out0 = ! v$Write_1964_out0;
assign v$G2_10350_out0 = ! v$Write_1965_out0;
assign v$G2_10351_out0 = ! v$Write_1966_out0;
assign v$G2_10352_out0 = ! v$Write_1967_out0;
assign v$G2_10353_out0 = ! v$Write_1968_out0;
assign v$G2_10354_out0 = ! v$Write_1969_out0;
assign v$G2_10355_out0 = ! v$Write_1970_out0;
assign v$_10491_out0 = v$_8866_out0[0:0];
assign v$_10491_out1 = v$_8866_out0[1:1];
assign v$_10492_out0 = v$_8867_out0[0:0];
assign v$_10492_out1 = v$_8867_out0[1:1];
assign v$7_10649_out0 = v$IR2_2660_out0[8:8];
assign v$7_10650_out0 = v$IR2_2661_out0[8:8];
assign v$ParityEN_11013_out0 = v$_4077_out0;
assign v$ParityEN_11014_out0 = v$_4078_out0;
assign v$_11057_out0 = v$_6415_out1[0:0];
assign v$_11057_out1 = v$_6415_out1[1:1];
assign v$_11058_out0 = v$_6416_out1[0:0];
assign v$_11058_out1 = v$_6416_out1[1:1];
assign v$RXCLK_11062_out0 = v$RXCLK_507_out0;
assign v$RXCLK_11063_out0 = v$RXCLK_508_out0;
assign v$SEL11_11105_out0 = v$IR2_2660_out0[7:7];
assign v$SEL11_11106_out0 = v$IR2_2661_out0[7:7];
assign v$C_11110_out0 = v$C_2344_out0;
assign v$C_11111_out0 = v$C_2345_out0;
assign v$R_11791_out0 = v$G3_11270_out0;
assign v$_11807_out0 = v$_11477_out1[7:0];
assign v$_11807_out1 = v$_11477_out1[15:8];
assign v$_11808_out0 = v$_11478_out1[7:0];
assign v$_11808_out1 = v$_11478_out1[15:8];
assign v$G39_11939_out0 = v$Q2_3703_out0 && v$G42_13143_out0;
assign v$G39_11940_out0 = v$Q2_3704_out0 && v$G42_13144_out0;
assign v$_12039_out0 = v$_3516_out0[0:0];
assign v$_12039_out1 = v$_3516_out0[1:1];
assign v$_12040_out0 = v$_3517_out0[0:0];
assign v$_12040_out1 = v$_3517_out0[1:1];
assign v$G21_12498_out0 = v$G23_1199_out0 && v$G22_2984_out0;
assign v$G21_12499_out0 = v$G23_1200_out0 && v$G22_2985_out0;
assign v$_12741_out0 = v$_13007_out1[0:0];
assign v$_12741_out1 = v$_13007_out1[1:1];
assign v$_12742_out0 = v$_13008_out1[0:0];
assign v$_12742_out1 = v$_13008_out1[1:1];
assign v$G31_13271_out0 = v$G32_6353_out0 && v$NQ3_1759_out0;
assign v$G31_13272_out0 = v$G32_6354_out0 && v$NQ3_1760_out0;
assign v$EQ2_13294_out0 = v$Q_4167_out0 == 4'h0;
assign v$EQ2_13295_out0 = v$Q_4168_out0 == 4'h0;
assign v$G56_372_out0 = v$EQ3_1515_out0 || v$EQ4_6581_out0;
assign v$G56_373_out0 = v$EQ3_1516_out0 || v$EQ4_6582_out0;
assign v$IR2$S_463_out0 = v$7_10649_out0;
assign v$IR2$S_464_out0 = v$7_10650_out0;
assign v$G9_473_out0 = ((v$_4885_out1 && !v$_9360_out1) || (!v$_4885_out1) && v$_9360_out1);
assign v$G9_474_out0 = ((v$_4886_out1 && !v$_9361_out1) || (!v$_4886_out1) && v$_9361_out1);
assign v$DATA$OUT_538_out0 = v$DATA$OUT_5146_out0;
assign v$DATA$OUT_539_out0 = v$DATA$OUT_5147_out0;
assign v$G4_559_out0 = ((v$_7862_out1 && !v$_5488_out1) || (!v$_7862_out1) && v$_5488_out1);
assign v$G4_560_out0 = ((v$_7863_out1 && !v$_5489_out1) || (!v$_7863_out1) && v$_5489_out1);
assign v$G47_753_out0 = v$PARITY_7858_out0 && v$EQ1_5014_out0;
assign v$G47_754_out0 = v$PARITY_7859_out0 && v$EQ1_5015_out0;
assign v$R_791_out0 = v$R_11791_out0;
assign v$_863_out0 = { v$C8_4879_out0,v$_8546_out0 };
assign v$_864_out0 = { v$C8_4880_out0,v$_8547_out0 };
assign v$IR2$FPU$OP_881_out0 = v$SEL4_6439_out0;
assign v$IR2$FPU$OP_882_out0 = v$SEL4_6440_out0;
assign v$G12_995_out0 = ((v$_6017_out1 && !v$_6473_out1) || (!v$_6017_out1) && v$_6473_out1);
assign v$G12_996_out0 = ((v$_6018_out1 && !v$_6474_out1) || (!v$_6018_out1) && v$_6474_out1);
assign v$G15_1030_out0 = ((v$_6017_out0 && !v$_6473_out0) || (!v$_6017_out0) && v$_6473_out0);
assign v$G15_1031_out0 = ((v$_6018_out0 && !v$_6474_out0) || (!v$_6018_out0) && v$_6474_out0);
assign v$G10_1141_out0 = ((v$_9644_out1 && !v$_11057_out1) || (!v$_9644_out1) && v$_11057_out1);
assign v$G10_1142_out0 = ((v$_9645_out1 && !v$_11058_out1) || (!v$_9645_out1) && v$_11058_out1);
assign v$G25_1387_out0 = v$IR2$IS$LDST_3050_out0 && v$IR2$S$WB_12240_out0;
assign v$G25_1388_out0 = v$IR2$IS$LDST_3051_out0 && v$IR2$S$WB_12241_out0;
assign v$G30_1389_out0 = v$G31_13271_out0 && v$Q2_12285_out0;
assign v$G30_1390_out0 = v$G31_13272_out0 && v$Q2_12286_out0;
assign v$2StopBits_2191_out0 = v$_2714_out1;
assign v$2StopBits_2192_out0 = v$_2715_out1;
assign v$G16_2222_out0 = ((v$_4885_out0 && !v$_9360_out0) || (!v$_4885_out0) && v$_9360_out0);
assign v$G16_2223_out0 = ((v$_4886_out0 && !v$_9361_out0) || (!v$_4886_out0) && v$_9361_out0);
assign v$S_2742_out0 = v$_12741_out1;
assign v$S_2743_out0 = v$_12742_out1;
assign v$IR2$FPU$LOAD_2912_out0 = v$SEL11_11105_out0;
assign v$IR2$FPU$LOAD_2913_out0 = v$SEL11_11106_out0;
assign v$G8_3224_out0 = ((v$_3183_out1 && !v$_6057_out1) || (!v$_3183_out1) && v$_6057_out1);
assign v$G8_3225_out0 = ((v$_3184_out1 && !v$_6058_out1) || (!v$_3184_out1) && v$_6058_out1);
assign v$_3390_out0 = v$IR2_1985_out0[14:12];
assign v$_3391_out0 = v$IR2_1986_out0[14:12];
assign v$G55_3437_out0 = v$G56_1877_out0 || v$G48_1203_out0;
assign v$G55_3438_out0 = v$G56_1878_out0 || v$G48_1204_out0;
assign v$G2_3675_out0 = ((v$_2732_out1 && !v$_9897_out1) || (!v$_2732_out1) && v$_9897_out1);
assign v$G2_3676_out0 = ((v$_2733_out1 && !v$_9898_out1) || (!v$_2733_out1) && v$_9898_out1);
assign v$G22_3708_out0 = v$G25_9956_out0 && v$R2_2554_out0;
assign v$G22_3709_out0 = v$G25_9957_out0 && v$R2_2555_out0;
assign v$G39_4047_out0 = v$G40_9224_out0 || v$G43_319_out0;
assign v$G39_4048_out0 = v$G40_9225_out0 || v$G43_320_out0;
assign v$G6_4177_out0 = ((v$_3805_out1 && !v$_12039_out1) || (!v$_3805_out1) && v$_12039_out1);
assign v$G6_4178_out0 = ((v$_3806_out1 && !v$_12040_out1) || (!v$_3806_out1) && v$_12040_out1);
assign v$PIN_4634_out0 = v$_11807_out1;
assign v$PIN_4635_out0 = v$_11807_out0;
assign v$PIN_4638_out0 = v$_8546_out1;
assign v$PIN_4640_out0 = v$_11808_out1;
assign v$PIN_4641_out0 = v$_11808_out0;
assign v$PIN_4644_out0 = v$_8547_out1;
assign v$_4751_out0 = v$IR2_1985_out0[7:4];
assign v$_4752_out0 = v$IR2_1986_out0[7:4];
assign v$_4871_out0 = v$IR2_1985_out0[4:0];
assign v$_4872_out0 = v$IR2_1986_out0[4:0];
assign v$IR2$15_5012_out0 = v$6_1094_out0;
assign v$IR2$15_5013_out0 = v$6_1095_out0;
assign v$IR2_5306_out0 = v$IR2_1985_out0;
assign v$IR2_5307_out0 = v$IR2_1986_out0;
assign v$G64_5316_out0 = v$EQ3_2888_out0 && v$G63_6734_out0;
assign v$G64_5317_out0 = v$EQ3_2889_out0 && v$G63_6735_out0;
assign v$G11_5747_out0 = ((v$_10491_out1 && !v$_2495_out1) || (!v$_10491_out1) && v$_2495_out1);
assign v$G11_5748_out0 = ((v$_10492_out1 && !v$_2496_out1) || (!v$_10492_out1) && v$_2496_out1);
assign v$CLK4_6074_out0 = v$RXCLK_11062_out0;
assign v$CLK4_6075_out0 = v$RXCLK_11063_out0;
assign v$RXBIT_6165_out0 = v$RX_4204_out0;
assign v$RXBIT_6166_out0 = v$RX_4205_out0;
assign v$G57_6225_out0 = v$EQ2_7440_out0 && v$G58_162_out0;
assign v$G57_6226_out0 = v$EQ2_7441_out0 && v$G58_163_out0;
assign v$G23_6562_out0 = v$FF3_10341_out0 && v$G21_4790_out0;
assign v$G23_6563_out0 = v$FF3_10342_out0 && v$G21_4791_out0;
assign v$G1_6877_out0 = ((v$_2732_out0 && !v$_9897_out0) || (!v$_2732_out0) && v$_9897_out0);
assign v$G1_6878_out0 = ((v$_2733_out0 && !v$_9898_out0) || (!v$_2733_out0) && v$_9898_out0);
assign v$OddParity_7008_out0 = v$_2714_out0;
assign v$OddParity_7009_out0 = v$_2715_out0;
assign v$Q1P_7261_out0 = v$G21_12498_out0;
assign v$Q1P_7262_out0 = v$G21_12499_out0;
assign v$_7432_out0 = v$IR2_1985_out0[9:9];
assign v$_7433_out0 = v$IR2_1986_out0[9:9];
assign v$G61_7438_out0 = v$EQ4_1519_out0 && v$P_5784_out0;
assign v$G61_7439_out0 = v$EQ4_1520_out0 && v$P_5785_out0;
assign v$IR2$FPU$32BIT_7600_out0 = v$SEL10_2841_out0;
assign v$IR2$FPU$32BIT_7601_out0 = v$SEL10_2842_out0;
assign v$G14_7830_out0 = ((v$_9644_out0 && !v$_11057_out0) || (!v$_9644_out0) && v$_11057_out0);
assign v$G14_7831_out0 = ((v$_9645_out0 && !v$_11058_out0) || (!v$_9645_out0) && v$_11058_out0);
assign v$G7_8288_out0 = ((v$_3183_out0 && !v$_6057_out0) || (!v$_3183_out0) && v$_6057_out0);
assign v$G7_8289_out0 = ((v$_3184_out0 && !v$_6058_out0) || (!v$_3184_out0) && v$_6058_out0);
assign v$G53_8369_out0 = v$EQ1_9709_out0 && v$G52_11142_out0;
assign v$G53_8370_out0 = v$EQ1_9710_out0 && v$G52_11143_out0;
assign v$_8506_out0 = v$PIN_4636_out0[3:0];
assign v$_8506_out1 = v$PIN_4636_out0[7:4];
assign v$_8509_out0 = v$PIN_4639_out0[3:0];
assign v$_8509_out1 = v$PIN_4639_out0[7:4];
assign v$_8512_out0 = v$PIN_4642_out0[3:0];
assign v$_8512_out1 = v$PIN_4642_out0[7:4];
assign v$_8515_out0 = v$PIN_4645_out0[3:0];
assign v$_8515_out1 = v$PIN_4645_out0[7:4];
assign v$IR2$M_8626_out0 = v$5_5074_out0;
assign v$IR2$M_8627_out0 = v$5_5075_out0;
assign v$G13_9010_out0 = ((v$_10491_out0 && !v$_2495_out0) || (!v$_10491_out0) && v$_2495_out0);
assign v$G13_9011_out0 = ((v$_10492_out0 && !v$_2496_out0) || (!v$_10492_out0) && v$_2496_out0);
assign v$G57_9018_out0 = v$G61_5755_out0 || v$G58_4796_out0;
assign v$G57_9019_out0 = v$G61_5756_out0 || v$G58_4797_out0;
assign v$G18_9091_out0 = ! v$C_11110_out0;
assign v$G18_9092_out0 = ! v$C_11111_out0;
assign v$IR2$D_9879_out0 = v$8_481_out0;
assign v$IR2$D_9880_out0 = v$8_482_out0;
assign v$G28_10029_out0 = v$IR2$IS$FPU_4798_out0 && v$EQ14_3730_out0;
assign v$G28_10030_out0 = v$IR2$IS$FPU_4799_out0 && v$EQ14_3731_out0;
assign v$G59_10432_out0 = v$G58_1431_out0 || v$G60_6463_out0;
assign v$G59_10433_out0 = v$G58_1432_out0 || v$G60_6464_out0;
assign v$G40_10438_out0 = v$Q1_7197_out0 && v$G39_11939_out0;
assign v$G40_10439_out0 = v$Q1_7198_out0 && v$G39_11940_out0;
assign v$G5_10553_out0 = ((v$_3805_out0 && !v$_12039_out0) || (!v$_3805_out0) && v$_12039_out0);
assign v$G5_10554_out0 = ((v$_3806_out0 && !v$_12040_out0) || (!v$_3806_out0) && v$_12040_out0);
assign v$IR2$FPU$LOADA_10585_out0 = v$SEL12_581_out0;
assign v$IR2$FPU$LOADA_10586_out0 = v$SEL12_582_out0;
assign v$G22_10639_out0 = ! v$C_11110_out0;
assign v$G22_10640_out0 = ! v$C_11111_out0;
assign v$G28_10902_out0 = v$STALL$PREV$CYCLE_3798_out0 || v$STP$SAVED_5106_out0;
assign v$G28_10903_out0 = v$STALL$PREV$CYCLE_3799_out0 || v$STP$SAVED_5107_out0;
assign v$END_10986_out0 = v$A1_9247_out1;
assign v$END_10987_out0 = v$A1_9248_out1;
assign v$ODDPARITY_11132_out0 = v$_12741_out0;
assign v$ODDPARITY_11133_out0 = v$_12742_out0;
assign v$SEL3_11722_out0 = v$IR2_1985_out0[15:12];
assign v$SEL3_11723_out0 = v$IR2_1986_out0[15:12];
assign v$_11788_out0 = v$IR2_1985_out0[3:2];
assign v$_11789_out0 = v$IR2_1986_out0[3:2];
assign v$G45_11949_out0 = ! v$P_5784_out0;
assign v$G45_11950_out0 = ! v$P_5785_out0;
assign v$G3_12256_out0 = ((v$_7862_out0 && !v$_5488_out0) || (!v$_7862_out0) && v$_5488_out0);
assign v$G3_12257_out0 = ((v$_7863_out0 && !v$_5489_out0) || (!v$_7863_out0) && v$_5489_out0);
assign v$_12787_out0 = v$IR2_1985_out0[8:8];
assign v$_12788_out0 = v$IR2_1986_out0[8:8];
assign v$IR2$OP_12789_out0 = v$9_9550_out0;
assign v$IR2$OP_12790_out0 = v$9_9551_out0;
assign v$G25_12841_out0 = v$G26_2796_out0 || v$G28_7730_out0;
assign v$G25_12842_out0 = v$G26_2797_out0 || v$G28_7731_out0;
assign v$R_13054_out0 = v$R_56_out0;
assign v$R_13055_out0 = v$R_57_out0;
assign v$EQ7_13267_out0 = v$IR2_1985_out0 == 16'h7000;
assign v$EQ7_13268_out0 = v$IR2_1986_out0 == 16'h7000;
assign v$G2_13322_out0 = v$RXENABLE_2429_out0 && v$RXCLK_11062_out0;
assign v$G2_13323_out0 = v$RXENABLE_2430_out0 && v$RXCLK_11063_out0;
assign v$RX_40_out0 = v$RXBIT_6165_out0;
assign v$RX_41_out0 = v$RXBIT_6166_out0;
assign v$G27_225_out0 = v$G1_6877_out0 || v$G2_3675_out0;
assign v$G27_226_out0 = v$G1_6878_out0 || v$G2_3676_out0;
assign v$K_253_out0 = v$_4871_out0;
assign v$K_254_out0 = v$_4872_out0;
assign v$G17_291_out0 = v$S_2742_out0 && v$NQ2_13211_out0;
assign v$G17_292_out0 = v$S_2743_out0 && v$NQ2_13212_out0;
assign v$G25_540_out0 = v$G5_10553_out0 || v$G6_4177_out0;
assign v$G25_541_out0 = v$G5_10554_out0 || v$G6_4178_out0;
assign v$OP_1032_out0 = v$IR2$OP_12789_out0;
assign v$OP_1033_out0 = v$IR2$OP_12790_out0;
assign v$RX_1727_out0 = v$RXBIT_6165_out0;
assign v$RX_1728_out0 = v$RXBIT_6166_out0;
assign v$G52_1732_out0 = v$S_2742_out0 || v$NQ0_10890_out0;
assign v$G52_1733_out0 = v$S_2743_out0 || v$NQ0_10891_out0;
assign v$C_1917_out0 = v$_7432_out0;
assign v$C_1918_out0 = v$_7433_out0;
assign v$G12_2328_out0 = ! v$IR2$FPU$LOADA_10585_out0;
assign v$G12_2329_out0 = ! v$IR2$FPU$LOADA_10586_out0;
assign v$IR1_2845_out0 = v$R_13054_out0;
assign v$IR1_2846_out0 = v$R_13055_out0;
assign v$IR2$VALID_2898_out0 = v$G59_10432_out0;
assign v$IR2$VALID_2899_out0 = v$G59_10433_out0;
assign v$RX_3217_out0 = v$RXBIT_6165_out0;
assign v$RX_3218_out0 = v$RXBIT_6166_out0;
assign v$LOADA_3519_out0 = v$IR2$FPU$LOADA_10585_out0;
assign v$LOADA_3520_out0 = v$IR2$FPU$LOADA_10586_out0;
assign v$S_3770_out0 = v$_12787_out0;
assign v$S_3771_out0 = v$_12788_out0;
assign v$G9_4349_out0 = ((v$G8_8068_out0 && !v$OddParity_7008_out0) || (!v$G8_8068_out0) && v$OddParity_7008_out0);
assign v$G9_4350_out0 = ((v$G8_8069_out0 && !v$OddParity_7009_out0) || (!v$G8_8069_out0) && v$OddParity_7009_out0);
assign v$PIN_4637_out0 = v$_863_out0;
assign v$PIN_4643_out0 = v$_864_out0;
assign v$NP_4857_out0 = v$G45_11949_out0;
assign v$NP_4858_out0 = v$G45_11950_out0;
assign v$OPCODE_5408_out0 = v$_3390_out0;
assign v$OPCODE_5409_out0 = v$_3391_out0;
assign v$SHIFT_5531_out0 = v$_11788_out0;
assign v$SHIFT_5532_out0 = v$_11789_out0;
assign v$_5910_out0 = v$_8506_out1[1:0];
assign v$_5910_out1 = v$_8506_out1[3:2];
assign v$_5913_out0 = v$_8509_out1[1:0];
assign v$_5913_out1 = v$_8509_out1[3:2];
assign v$_5916_out0 = v$_8512_out1[1:0];
assign v$_5916_out1 = v$_8512_out1[3:2];
assign v$_5919_out0 = v$_8515_out1[1:0];
assign v$_5919_out1 = v$_8515_out1[3:2];
assign v$G17_6070_out0 = v$G13_9010_out0 || v$G11_5747_out0;
assign v$G17_6071_out0 = v$G13_9011_out0 || v$G11_5748_out0;
assign v$RXFlagSet_6347_out0 = v$G53_8369_out0;
assign v$RXFlagSet_6348_out0 = v$G53_8370_out0;
assign v$G24_6574_out0 = v$NQ3_721_out0 && v$G25_12841_out0;
assign v$G24_6575_out0 = v$NQ3_722_out0 && v$G25_12842_out0;
assign v$EQ10_6613_out0 = v$IR2$FPU$OP_881_out0 == 2'h3;
assign v$EQ10_6614_out0 = v$IR2$FPU$OP_882_out0 == 2'h3;
assign v$G27_6811_out0 = v$S_2742_out0 && v$NQ2_13211_out0;
assign v$G27_6812_out0 = v$S_2743_out0 && v$NQ2_13212_out0;
assign v$G18_6825_out0 = v$G16_2222_out0 || v$G9_473_out0;
assign v$G18_6826_out0 = v$G16_2223_out0 || v$G9_474_out0;
assign v$G70_6845_out0 = v$S_2742_out0 && v$EQ6_773_out0;
assign v$G70_6846_out0 = v$S_2743_out0 && v$EQ6_774_out0;
assign v$G24_6893_out0 = v$G7_8288_out0 || v$G8_3224_out0;
assign v$G24_6894_out0 = v$G7_8289_out0 || v$G8_3225_out0;
assign v$IR15_7010_out0 = v$IR2$15_5012_out0;
assign v$IR15_7011_out0 = v$IR2$15_5013_out0;
assign v$G46_7181_out0 = ! v$S_2742_out0;
assign v$G46_7182_out0 = ! v$S_2743_out0;
assign v$32BIT_7201_out0 = v$IR2$FPU$32BIT_7600_out0;
assign v$32BIT_7202_out0 = v$IR2$FPU$32BIT_7601_out0;
assign v$LOAD_7522_out0 = v$IR2$FPU$LOAD_2912_out0;
assign v$LOAD_7523_out0 = v$IR2$FPU$LOAD_2913_out0;
assign v$G20_7530_out0 = v$G23_6562_out0 && v$F2_7871_out0;
assign v$G20_7531_out0 = v$G23_6563_out0 && v$F2_7872_out0;
assign v$IR2$FULL$OP$CODE_7620_out0 = v$SEL3_11722_out0;
assign v$IR2$FULL$OP$CODE_7621_out0 = v$SEL3_11723_out0;
assign v$CLK4_7986_out0 = v$G2_13322_out0;
assign v$CLK4_7987_out0 = v$G2_13323_out0;
assign v$G20_8393_out0 = v$G15_1030_out0 || v$G12_995_out0;
assign v$G20_8394_out0 = v$G15_1031_out0 || v$G12_996_out0;
assign v$SHIFTEN_8420_out0 = v$G57_9018_out0;
assign v$SHIFTEN_8421_out0 = v$G57_9019_out0;
assign v$_8486_out0 = v$_8506_out0[1:0];
assign v$_8486_out1 = v$_8506_out0[3:2];
assign v$_8489_out0 = v$_8509_out0[1:0];
assign v$_8489_out1 = v$_8509_out0[3:2];
assign v$_8492_out0 = v$_8512_out0[1:0];
assign v$_8492_out1 = v$_8512_out0[3:2];
assign v$_8495_out0 = v$_8515_out0[1:0];
assign v$_8495_out1 = v$_8515_out0[3:2];
assign v$_8504_out0 = v$PIN_4634_out0[3:0];
assign v$_8504_out1 = v$PIN_4634_out0[7:4];
assign v$_8505_out0 = v$PIN_4635_out0[3:0];
assign v$_8505_out1 = v$PIN_4635_out0[7:4];
assign v$_8508_out0 = v$PIN_4638_out0[3:0];
assign v$_8508_out1 = v$PIN_4638_out0[7:4];
assign v$_8510_out0 = v$PIN_4640_out0[3:0];
assign v$_8510_out1 = v$PIN_4640_out0[7:4];
assign v$_8511_out0 = v$PIN_4641_out0[3:0];
assign v$_8511_out1 = v$PIN_4641_out0[7:4];
assign v$_8514_out0 = v$PIN_4644_out0[3:0];
assign v$_8514_out1 = v$PIN_4644_out0[7:4];
assign v$B_8806_out0 = v$_4751_out0;
assign v$B_8807_out0 = v$_4752_out0;
assign v$G54_9597_out0 = v$G28_10902_out0 || v$HALT$PREV_6935_out0;
assign v$G54_9598_out0 = v$G28_10903_out0 || v$HALT$PREV_6936_out0;
assign v$G21_9642_out0 = v$G14_7830_out0 || v$G10_1141_out0;
assign v$G21_9643_out0 = v$G14_7831_out0 || v$G10_1142_out0;
assign v$G26_10232_out0 = v$G3_12256_out0 || v$G4_559_out0;
assign v$G26_10233_out0 = v$G3_12257_out0 || v$G4_560_out0;
assign v$G66_10587_out0 = ((v$ODDPARITY_11132_out0 && !v$EVENPARITY_9157_out0) || (!v$ODDPARITY_11132_out0) && v$EVENPARITY_9157_out0);
assign v$G66_10588_out0 = ((v$ODDPARITY_11133_out0 && !v$EVENPARITY_9158_out0) || (!v$ODDPARITY_11133_out0) && v$EVENPARITY_9158_out0);
assign v$G46_11285_out0 = v$G55_3437_out0 || v$G47_3665_out0;
assign v$G46_11286_out0 = v$G55_3438_out0 || v$G47_3666_out0;
assign v$ParityCheck_11289_out0 = v$G57_6225_out0;
assign v$ParityCheck_11290_out0 = v$G57_6226_out0;
assign v$G32_11448_out0 = v$G35_8276_out0 || v$G40_10438_out0;
assign v$G32_11449_out0 = v$G35_8277_out0 || v$G40_10439_out0;
assign v$RXReset_11610_out0 = v$G64_5316_out0;
assign v$RXReset_11611_out0 = v$G64_5317_out0;
assign v$G55_11730_out0 = v$EQ2_13294_out0 || v$G56_372_out0;
assign v$G55_11731_out0 = v$EQ2_13295_out0 || v$G56_373_out0;
assign v$RAMDOUT_11827_out0 = v$DATA$OUT_538_out0;
assign v$RAMDOUT_11828_out0 = v$DATA$OUT_539_out0;
assign v$G63_11847_out0 = v$G57_9018_out0 && v$SERIALIN_3766_out0;
assign v$G63_11848_out0 = v$G57_9019_out0 && v$SERIALIN_3767_out0;
assign v$MUX4_12118_out0 = v$G47_753_out0 ? v$C4_1692_out0 : v$G39_4047_out0;
assign v$MUX4_12119_out0 = v$G47_754_out0 ? v$C4_1693_out0 : v$G39_4048_out0;
assign v$G3_12515_out0 = ! v$R_791_out0;
assign v$G9_12526_out0 = ! v$EQ7_13267_out0;
assign v$G9_12527_out0 = ! v$EQ7_13268_out0;
assign v$IR2_12729_out0 = v$IR2_5306_out0;
assign v$IR2_12730_out0 = v$IR2_5307_out0;
assign v$CHECKPARITY_557_out0 = v$ParityCheck_11289_out0;
assign v$CHECKPARITY_558_out0 = v$ParityCheck_11290_out0;
assign v$1_755_out0 = v$IR2_12729_out0[8:8];
assign v$1_756_out0 = v$IR2_12730_out0[8:8];
assign v$_839_out0 = v$_8486_out1[0:0];
assign v$_839_out1 = v$_8486_out1[1:1];
assign v$_842_out0 = v$_8489_out1[0:0];
assign v$_842_out1 = v$_8489_out1[1:1];
assign v$_845_out0 = v$_8492_out1[0:0];
assign v$_845_out1 = v$_8492_out1[1:1];
assign v$_848_out0 = v$_8495_out1[0:0];
assign v$_848_out1 = v$_8495_out1[1:1];
assign v$G65_1383_out0 = v$EQ5_6345_out0 && v$G66_10587_out0;
assign v$G65_1384_out0 = v$EQ5_6346_out0 && v$G66_10588_out0;
assign v$CLK4_1439_out0 = v$CLK4_7986_out0;
assign v$CLK4_1440_out0 = v$CLK4_7987_out0;
assign v$G10_1683_out0 = ((v$G9_4349_out0 && !v$RceivedParity_13191_out0) || (!v$G9_4349_out0) && v$RceivedParity_13191_out0);
assign v$G10_1684_out0 = ((v$G9_4350_out0 && !v$RceivedParity_13192_out0) || (!v$G9_4350_out0) && v$RceivedParity_13192_out0);
assign v$SEL6_1769_out0 = v$IR1_2845_out0[1:0];
assign v$SEL6_1770_out0 = v$IR1_2846_out0[1:0];
assign v$G11_1955_out0 = v$IR2$FPU$LOAD_2912_out0 && v$G12_2328_out0;
assign v$G11_1956_out0 = v$IR2$FPU$LOAD_2913_out0 && v$G12_2329_out0;
assign v$SEL2_2427_out0 = v$IR1_2845_out0[8:8];
assign v$SEL2_2428_out0 = v$IR1_2846_out0[8:8];
assign v$Q2P_2850_out0 = v$G24_6574_out0;
assign v$Q2P_2851_out0 = v$G24_6575_out0;
assign v$S_2914_out0 = v$S_3770_out0;
assign v$S_2915_out0 = v$S_3771_out0;
assign v$LOADA_3453_out0 = v$LOADA_3519_out0;
assign v$LOADA_3454_out0 = v$LOADA_3520_out0;
assign v$C_4069_out0 = v$C_1917_out0;
assign v$C_4070_out0 = v$C_1918_out0;
assign v$LOAD_4208_out0 = v$LOAD_7522_out0;
assign v$LOAD_4209_out0 = v$LOAD_7523_out0;
assign v$EQ6_4423_out0 = v$IR2$FULL$OP$CODE_7620_out0 == 4'h7;
assign v$EQ6_4424_out0 = v$IR2$FULL$OP$CODE_7621_out0 == 4'h7;
assign v$SHIFT_4778_out0 = v$SHIFT_5531_out0;
assign v$SHIFT_4779_out0 = v$SHIFT_5532_out0;
assign v$_5189_out0 = v$_8486_out0[0:0];
assign v$_5189_out1 = v$_8486_out0[1:1];
assign v$_5192_out0 = v$_8489_out0[0:0];
assign v$_5192_out1 = v$_8489_out0[1:1];
assign v$_5195_out0 = v$_8492_out0[0:0];
assign v$_5195_out1 = v$_8492_out0[1:1];
assign v$_5198_out0 = v$_8495_out0[0:0];
assign v$_5198_out1 = v$_8495_out0[1:1];
assign v$SEL9_5490_out0 = v$IR1_2845_out0[11:10];
assign v$SEL9_5491_out0 = v$IR1_2846_out0[11:10];
assign v$G54_5642_out0 = v$G55_11730_out0 || v$G63_11847_out0;
assign v$G54_5643_out0 = v$G55_11731_out0 || v$G63_11848_out0;
assign v$_5908_out0 = v$_8504_out1[1:0];
assign v$_5908_out1 = v$_8504_out1[3:2];
assign v$_5909_out0 = v$_8505_out1[1:0];
assign v$_5909_out1 = v$_8505_out1[3:2];
assign v$_5912_out0 = v$_8508_out1[1:0];
assign v$_5912_out1 = v$_8508_out1[3:2];
assign v$_5914_out0 = v$_8510_out1[1:0];
assign v$_5914_out1 = v$_8510_out1[3:2];
assign v$_5915_out0 = v$_8511_out1[1:0];
assign v$_5915_out1 = v$_8511_out1[3:2];
assign v$_5918_out0 = v$_8514_out1[1:0];
assign v$_5918_out1 = v$_8514_out1[3:2];
assign v$R_6019_out0 = v$RX_3217_out0;
assign v$R_6020_out0 = v$RX_3218_out0;
assign v$SEL1_6041_out0 = v$IR1_2845_out0[15:12];
assign v$SEL1_6042_out0 = v$IR1_2846_out0[15:12];
assign v$6_6615_out0 = v$IR2_12729_out0[7:7];
assign v$6_6616_out0 = v$IR2_12730_out0[7:7];
assign v$SHIFTEN_6847_out0 = v$SHIFTEN_8420_out0;
assign v$SHIFTEN_6848_out0 = v$SHIFTEN_8421_out0;
assign v$G26_6879_out0 = v$G22_3708_out0 || v$G20_7530_out0;
assign v$G26_6880_out0 = v$G22_3709_out0 || v$G20_7531_out0;
assign v$G28_7110_out0 = v$G27_225_out0 || v$G26_10232_out0;
assign v$G28_7111_out0 = v$G27_226_out0 || v$G26_10233_out0;
assign v$IR15_7240_out0 = v$IR15_7010_out0;
assign v$IR15_7241_out0 = v$IR15_7011_out0;
assign v$G18_7271_out0 = v$IR2$FPU$LOAD_2912_out0 && v$EQ10_6613_out0;
assign v$G18_7272_out0 = v$IR2$FPU$LOAD_2913_out0 && v$EQ10_6614_out0;
assign v$Q3P_7500_out0 = v$MUX4_12118_out0;
assign v$Q3P_7501_out0 = v$MUX4_12119_out0;
assign v$IR2$VALID_7594_out0 = v$IR2$VALID_2898_out0;
assign v$IR2$VALID_7595_out0 = v$IR2$VALID_2899_out0;
assign v$G11_7645_out0 = v$Q3_13107_out0 && v$G52_1732_out0;
assign v$G11_7646_out0 = v$Q3_13108_out0 && v$G52_1733_out0;
assign v$_7655_out0 = v$_5910_out1[0:0];
assign v$_7655_out1 = v$_5910_out1[1:1];
assign v$_7658_out0 = v$_5913_out1[0:0];
assign v$_7658_out1 = v$_5913_out1[1:1];
assign v$_7661_out0 = v$_5916_out1[0:0];
assign v$_7661_out1 = v$_5916_out1[1:1];
assign v$_7664_out0 = v$_5919_out1[0:0];
assign v$_7664_out1 = v$_5919_out1[1:1];
assign v$EQ11_7677_out0 = v$IR2$FULL$OP$CODE_7620_out0 == 4'h1;
assign v$EQ11_7678_out0 = v$IR2$FULL$OP$CODE_7621_out0 == 4'h1;
assign v$SEL11_7974_out0 = v$IR2_12729_out0[7:7];
assign v$SEL11_7975_out0 = v$IR2_12730_out0[7:7];
assign v$_8000_out0 = { v$K_253_out0,v$C1_11027_out0 };
assign v$_8001_out0 = { v$K_254_out0,v$C1_11028_out0 };
assign v$5_8062_out0 = v$IR2_12729_out0[9:9];
assign v$5_8063_out0 = v$IR2_12730_out0[9:9];
assign v$EQ4_8382_out0 = v$IR2_12729_out0 == 16'h7000;
assign v$EQ4_8383_out0 = v$IR2_12730_out0 == 16'h7000;
assign v$2_8391_out0 = v$IR2_12729_out0[11:10];
assign v$2_8392_out0 = v$IR2_12730_out0[11:10];
assign v$SEL10_8472_out0 = v$IR2_12729_out0[9:8];
assign v$SEL10_8473_out0 = v$IR2_12730_out0[9:8];
assign v$_8484_out0 = v$_8504_out0[1:0];
assign v$_8484_out1 = v$_8504_out0[3:2];
assign v$_8485_out0 = v$_8505_out0[1:0];
assign v$_8485_out1 = v$_8505_out0[3:2];
assign v$_8488_out0 = v$_8508_out0[1:0];
assign v$_8488_out1 = v$_8508_out0[3:2];
assign v$_8490_out0 = v$_8510_out0[1:0];
assign v$_8490_out1 = v$_8510_out0[3:2];
assign v$_8491_out0 = v$_8511_out0[1:0];
assign v$_8491_out1 = v$_8511_out0[3:2];
assign v$_8494_out0 = v$_8514_out0[1:0];
assign v$_8494_out1 = v$_8514_out0[3:2];
assign v$_8507_out0 = v$PIN_4637_out0[3:0];
assign v$_8507_out1 = v$PIN_4637_out0[7:4];
assign v$_8513_out0 = v$PIN_4643_out0[3:0];
assign v$_8513_out1 = v$PIN_4643_out0[7:4];
assign v$G1_8623_out0 = v$STATE_11198_out0 && v$G3_12515_out0;
assign v$EQ12_8848_out0 = v$IR2$FULL$OP$CODE_7620_out0 == 4'h1;
assign v$EQ12_8849_out0 = v$IR2$FULL$OP$CODE_7621_out0 == 4'h1;
assign v$3_8971_out0 = v$IR2_12729_out0[5:2];
assign v$3_8972_out0 = v$IR2_12730_out0[5:2];
assign v$Q3P_9332_out0 = v$G32_11448_out0;
assign v$Q3P_9333_out0 = v$G32_11449_out0;
assign v$G29_9392_out0 = v$G25_540_out0 || v$G24_6893_out0;
assign v$G29_9393_out0 = v$G25_541_out0 || v$G24_6894_out0;
assign v$7_9409_out0 = v$IR2_12729_out0[1:0];
assign v$7_9410_out0 = v$IR2_12730_out0[1:0];
assign v$9_9707_out0 = v$IR2_12729_out0[15:12];
assign v$9_9708_out0 = v$IR2_12730_out0[15:12];
assign v$G2_9887_out0 = ((v$RX_40_out0 && !v$FF3_4929_out0) || (!v$RX_40_out0) && v$FF3_4929_out0);
assign v$G2_9888_out0 = ((v$RX_41_out0 && !v$FF3_4930_out0) || (!v$RX_41_out0) && v$FF3_4930_out0);
assign v$_9901_out0 = v$_5910_out0[0:0];
assign v$_9901_out1 = v$_5910_out0[1:1];
assign v$_9904_out0 = v$_5913_out0[0:0];
assign v$_9904_out1 = v$_5913_out0[1:1];
assign v$_9907_out0 = v$_5916_out0[0:0];
assign v$_9907_out1 = v$_5916_out0[1:1];
assign v$_9910_out0 = v$_5919_out0[0:0];
assign v$_9910_out1 = v$_5919_out0[1:1];
assign v$B_9992_out0 = v$B_8806_out0;
assign v$B_9993_out0 = v$B_8807_out0;
assign v$RXSET_10048_out0 = v$RXFlagSet_6347_out0;
assign v$RXSET_10049_out0 = v$RXFlagSet_6348_out0;
assign v$RXINTERRUPT_10185_out0 = v$RXReset_11610_out0;
assign v$RXINTERRUPT_10186_out0 = v$RXReset_11611_out0;
assign v$SEL8_10430_out0 = v$IR1_2845_out0[9:8];
assign v$SEL8_10431_out0 = v$IR1_2846_out0[9:8];
assign v$4_10457_out0 = v$IR2_12729_out0[6:6];
assign v$4_10458_out0 = v$IR2_12730_out0[6:6];
assign v$MUX1_10579_out0 = v$G54_9597_out0 ? v$REG3_1589_out0 : v$R_13054_out0;
assign v$MUX1_10580_out0 = v$G54_9598_out0 ? v$REG3_1590_out0 : v$R_13055_out0;
assign v$8_10817_out0 = v$IR2_12729_out0[15:15];
assign v$8_10818_out0 = v$IR2_12730_out0[15:15];
assign v$SEL7_10884_out0 = v$IR1_2845_out0[9:9];
assign v$SEL7_10885_out0 = v$IR1_2846_out0[9:9];
assign v$G53_11048_out0 = v$G17_291_out0 || v$NQ3_1759_out0;
assign v$G53_11049_out0 = v$G17_292_out0 || v$NQ3_1760_out0;
assign v$G22_11070_out0 = v$G20_8393_out0 || v$G21_9642_out0;
assign v$G22_11071_out0 = v$G20_8394_out0 || v$G21_9643_out0;
assign v$32BIT_11086_out0 = v$32BIT_7201_out0;
assign v$32BIT_11087_out0 = v$32BIT_7202_out0;
assign v$G19_11146_out0 = v$G17_6070_out0 || v$G18_6825_out0;
assign v$G19_11147_out0 = v$G17_6071_out0 || v$G18_6826_out0;
assign v$G26_11205_out0 = v$NQ3_1759_out0 || v$G27_6811_out0;
assign v$G26_11206_out0 = v$NQ3_1760_out0 || v$G27_6812_out0;
assign v$EQ1_11291_out0 = v$OPCODE_5408_out0 == 3'h4;
assign v$EQ1_11292_out0 = v$OPCODE_5409_out0 == 3'h4;
assign v$ShiftOut_11458_out0 = v$G46_11285_out0;
assign v$ShiftOut_11459_out0 = v$G46_11286_out0;
assign v$OP_12461_out0 = v$OP_1032_out0;
assign v$OP_12462_out0 = v$OP_1033_out0;
assign v$G10_12927_out0 = v$NP_4857_out0 && v$G11_3264_out0;
assign v$G10_12928_out0 = v$NP_4858_out0 && v$G11_3265_out0;
assign v$NS_12937_out0 = v$G46_7181_out0;
assign v$NS_12938_out0 = v$G46_7182_out0;
assign v$EQ9_12993_out0 = v$IR2$FULL$OP$CODE_7620_out0 == 4'h1;
assign v$EQ9_12994_out0 = v$IR2$FULL$OP$CODE_7621_out0 == 4'h1;
assign v$EQ1_13237_out0 = v$IR2$FULL$OP$CODE_7620_out0 == 4'h1;
assign v$EQ1_13238_out0 = v$IR2$FULL$OP$CODE_7621_out0 == 4'h1;
assign v$IR1$S$WB_264_out0 = v$SEL2_2427_out0;
assign v$IR1$S$WB_265_out0 = v$SEL2_2428_out0;
assign v$RXSHIFT_388_out0 = v$ShiftOut_11458_out0;
assign v$RXSHIFT_389_out0 = v$ShiftOut_11459_out0;
assign v$G69_489_out0 = ! v$R_6019_out0;
assign v$G69_490_out0 = ! v$R_6020_out0;
assign v$_837_out0 = v$_8484_out1[0:0];
assign v$_837_out1 = v$_8484_out1[1:1];
assign v$_838_out0 = v$_8485_out1[0:0];
assign v$_838_out1 = v$_8485_out1[1:1];
assign v$_841_out0 = v$_8488_out1[0:0];
assign v$_841_out1 = v$_8488_out1[1:1];
assign v$_843_out0 = v$_8490_out1[0:0];
assign v$_843_out1 = v$_8490_out1[1:1];
assign v$_844_out0 = v$_8491_out1[0:0];
assign v$_844_out1 = v$_8491_out1[1:1];
assign v$_847_out0 = v$_8494_out1[0:0];
assign v$_847_out1 = v$_8494_out1[1:1];
assign v$EQ1_1429_out0 = v$OP_12461_out0 == 3'h4;
assign v$EQ1_1430_out0 = v$OP_12462_out0 == 3'h4;
assign v$IR2$OPCODE_1482_out0 = v$9_9707_out0;
assign v$IR2$OPCODE_1483_out0 = v$9_9708_out0;
assign v$MUX1_1491_out0 = v$G2_10346_out0 ? v$SIN_86_out0 : v$_5189_out0;
assign v$MUX1_1494_out0 = v$G2_10349_out0 ? v$SIN_89_out0 : v$_5192_out0;
assign v$MUX1_1497_out0 = v$G2_10352_out0 ? v$SIN_92_out0 : v$_5195_out0;
assign v$MUX1_1500_out0 = v$G2_10355_out0 ? v$SIN_95_out0 : v$_5198_out0;
assign v$_1554_out0 = v$OP_12461_out0[0:0];
assign v$_1555_out0 = v$OP_12462_out0[0:0];
assign v$IR2$FPU$OP_1657_out0 = v$SEL10_8472_out0;
assign v$IR2$FPU$OP_1658_out0 = v$SEL10_8473_out0;
assign v$IR2$IS$FPU_1696_out0 = v$EQ12_8848_out0;
assign v$IR2$IS$FPU_1697_out0 = v$EQ12_8849_out0;
assign v$_1743_out0 = v$OP_12461_out0[2:2];
assign v$_1744_out0 = v$OP_12462_out0[2:2];
assign v$IR2$N_1745_out0 = v$3_8971_out0;
assign v$IR2$N_1746_out0 = v$3_8972_out0;
assign v$MUX8_2318_out0 = v$G2_10346_out0 ? v$FF2_10135_out0 : v$_9901_out0;
assign v$MUX8_2321_out0 = v$G2_10349_out0 ? v$FF2_10138_out0 : v$_9904_out0;
assign v$MUX8_2324_out0 = v$G2_10352_out0 ? v$FF2_10141_out0 : v$_9907_out0;
assign v$MUX8_2327_out0 = v$G2_10355_out0 ? v$FF2_10144_out0 : v$_9910_out0;
assign v$B_2417_out0 = v$B_9992_out0;
assign v$B_2418_out0 = v$B_9993_out0;
assign v$G23_3040_out0 = v$G19_11146_out0 || v$G22_11070_out0;
assign v$G23_3041_out0 = v$G19_11147_out0 || v$G22_11071_out0;
assign v$IR2$D_3290_out0 = v$2_8391_out0;
assign v$IR2$D_3291_out0 = v$2_8392_out0;
assign v$RXset_3477_out0 = v$RXSET_10048_out0;
assign v$RXset_3478_out0 = v$RXSET_10049_out0;
assign v$EQ4_3659_out0 = v$SEL8_10430_out0 == 2'h2;
assign v$EQ4_3660_out0 = v$SEL8_10431_out0 == 2'h2;
assign v$IR1$RD_3732_out0 = v$SEL9_5490_out0;
assign v$IR1$RD_3733_out0 = v$SEL9_5491_out0;
assign v$IR2$U_3921_out0 = v$4_10457_out0;
assign v$IR2$U_3922_out0 = v$4_10458_out0;
assign v$G14_4141_out0 = v$G15_2890_out0 && v$G53_11048_out0;
assign v$G14_4142_out0 = v$G15_2891_out0 && v$G53_11049_out0;
assign v$ISMOV_4660_out0 = v$EQ1_11291_out0;
assign v$ISMOV_4661_out0 = v$EQ1_11292_out0;
assign v$SHIFTEN_4821_out0 = v$SHIFTEN_6847_out0;
assign v$SHIFTEN_4822_out0 = v$SHIFTEN_6848_out0;
assign v$G2_5117_out0 = v$G1_8623_out0 || v$S_5524_out0;
assign v$_5187_out0 = v$_8484_out0[0:0];
assign v$_5187_out1 = v$_8484_out0[1:1];
assign v$_5188_out0 = v$_8485_out0[0:0];
assign v$_5188_out1 = v$_8485_out0[1:1];
assign v$_5191_out0 = v$_8488_out0[0:0];
assign v$_5191_out1 = v$_8488_out0[1:1];
assign v$_5193_out0 = v$_8490_out0[0:0];
assign v$_5193_out1 = v$_8490_out0[1:1];
assign v$_5194_out0 = v$_8491_out0[0:0];
assign v$_5194_out1 = v$_8491_out0[1:1];
assign v$_5197_out0 = v$_8494_out0[0:0];
assign v$_5197_out1 = v$_8494_out0[1:1];
assign v$EQ2_5448_out0 = v$OP_12461_out0 == 3'h5;
assign v$EQ2_5449_out0 = v$OP_12462_out0 == 3'h5;
assign v$S_5664_out0 = v$S_2914_out0;
assign v$S_5665_out0 = v$S_2915_out0;
assign v$G69_5702_out0 = v$EQ7_201_out0 && v$NS_12937_out0;
assign v$G69_5703_out0 = v$EQ7_202_out0 && v$NS_12938_out0;
assign v$_5720_out0 = v$OP_12461_out0[1:1];
assign v$_5721_out0 = v$OP_12462_out0[1:1];
assign v$STOP$2_5722_out0 = v$EQ4_8382_out0;
assign v$STOP$2_5723_out0 = v$EQ4_8383_out0;
assign v$_5911_out0 = v$_8507_out1[1:0];
assign v$_5911_out1 = v$_8507_out1[3:2];
assign v$_5917_out0 = v$_8513_out1[1:0];
assign v$_5917_out1 = v$_8513_out1[3:2];
assign v$IR2$M_6072_out0 = v$7_9409_out0;
assign v$IR2$M_6073_out0 = v$7_9410_out0;
assign v$G8_6485_out0 = v$G9_9012_out0 && v$G11_7645_out0;
assign v$G8_6486_out0 = v$G9_9013_out0 && v$G11_7646_out0;
assign v$MUX5_6502_out0 = v$G2_10346_out0 ? v$FF5_935_out0 : v$_5189_out1;
assign v$MUX5_6505_out0 = v$G2_10349_out0 ? v$FF5_938_out0 : v$_5192_out1;
assign v$MUX5_6508_out0 = v$G2_10352_out0 ? v$FF5_941_out0 : v$_5195_out1;
assign v$MUX5_6511_out0 = v$G2_10355_out0 ? v$FF5_944_out0 : v$_5198_out1;
assign v$IR1$OPCODE_6530_out0 = v$SEL1_6041_out0;
assign v$IR1$OPCODE_6531_out0 = v$SEL1_6042_out0;
assign v$_6546_out0 = v$OP_12461_out0[2:2];
assign v$_6547_out0 = v$OP_12462_out0[2:2];
assign v$C_6570_out0 = v$C_4069_out0;
assign v$C_6571_out0 = v$C_4070_out0;
assign v$MUX3_6672_out0 = v$G2_10346_out0 ? v$FF7_5774_out0 : v$_9901_out1;
assign v$MUX3_6675_out0 = v$G2_10349_out0 ? v$FF7_5777_out0 : v$_9904_out1;
assign v$MUX3_6678_out0 = v$G2_10352_out0 ? v$FF7_5780_out0 : v$_9907_out1;
assign v$MUX3_6681_out0 = v$G2_10355_out0 ? v$FF7_5783_out0 : v$_9910_out1;
assign v$IR1$C$L_6754_out0 = v$SEL7_10884_out0;
assign v$IR1$C$L_6755_out0 = v$SEL7_10885_out0;
assign v$G10_6837_out0 = v$EQ6_4423_out0 && v$G9_12526_out0;
assign v$G10_6838_out0 = v$EQ6_4424_out0 && v$G9_12527_out0;
assign v$_6843_out0 = v$OP_12461_out0[1:1];
assign v$_6844_out0 = v$OP_12462_out0[1:1];
assign v$MUX6_6939_out0 = v$G2_10346_out0 ? v$FF1_11257_out0 : v$_839_out1;
assign v$MUX6_6942_out0 = v$G2_10349_out0 ? v$FF1_11260_out0 : v$_842_out1;
assign v$MUX6_6945_out0 = v$G2_10352_out0 ? v$FF1_11263_out0 : v$_845_out1;
assign v$MUX6_6948_out0 = v$G2_10355_out0 ? v$FF1_11266_out0 : v$_848_out1;
assign v$IR2$FPU$L_7070_out0 = v$SEL11_7974_out0;
assign v$IR2$FPU$L_7071_out0 = v$SEL11_7975_out0;
assign v$IS$32$BIT_7259_out0 = v$32BIT_11086_out0;
assign v$IS$32$BIT_7260_out0 = v$32BIT_11087_out0;
assign v$G62_7570_out0 = v$G61_7438_out0 && v$CLK4_1439_out0;
assign v$G62_7571_out0 = v$G61_7439_out0 && v$CLK4_1440_out0;
assign v$_7653_out0 = v$_5908_out1[0:0];
assign v$_7653_out1 = v$_5908_out1[1:1];
assign v$_7654_out0 = v$_5909_out1[0:0];
assign v$_7654_out1 = v$_5909_out1[1:1];
assign v$_7657_out0 = v$_5912_out1[0:0];
assign v$_7657_out1 = v$_5912_out1[1:1];
assign v$_7659_out0 = v$_5914_out1[0:0];
assign v$_7659_out1 = v$_5914_out1[1:1];
assign v$_7660_out0 = v$_5915_out1[0:0];
assign v$_7660_out1 = v$_5915_out1[1:1];
assign v$_7663_out0 = v$_5918_out1[0:0];
assign v$_7663_out1 = v$_5918_out1[1:1];
assign v$G20_8064_out0 = ! v$LOAD_4208_out0;
assign v$G20_8065_out0 = ! v$LOAD_4209_out0;
assign v$IR2$L_8105_out0 = v$5_8062_out0;
assign v$IR2$L_8106_out0 = v$5_8063_out0;
assign v$_8487_out0 = v$_8507_out0[1:0];
assign v$_8487_out1 = v$_8507_out0[3:2];
assign v$_8493_out0 = v$_8513_out0[1:0];
assign v$_8493_out1 = v$_8513_out0[3:2];
assign v$_8688_out0 = { v$Q2P_2850_out0,v$Q3P_9332_out0 };
assign v$_8689_out0 = { v$Q2P_2851_out0,v$Q3P_9333_out0 };
assign v$G11_8976_out0 = ! v$LOAD_4208_out0;
assign v$G11_8977_out0 = ! v$LOAD_4209_out0;
assign v$_9237_out0 = v$OP_12461_out0[0:0];
assign v$_9238_out0 = v$OP_12462_out0[0:0];
assign v$MUX2_9344_out0 = v$G2_10346_out0 ? v$FF8_9845_out0 : v$_7655_out1;
assign v$MUX2_9347_out0 = v$G2_10349_out0 ? v$FF8_9848_out0 : v$_7658_out1;
assign v$MUX2_9350_out0 = v$G2_10352_out0 ? v$FF8_9851_out0 : v$_7661_out1;
assign v$MUX2_9353_out0 = v$G2_10355_out0 ? v$FF8_9854_out0 : v$_7664_out1;
assign v$IS$32$BITS_9430_out0 = v$32BIT_11086_out0;
assign v$IS$32$BITS_9431_out0 = v$32BIT_11087_out0;
assign v$B$IS$RD_9476_out0 = v$G11_1955_out0;
assign v$B$IS$RD_9477_out0 = v$G11_1956_out0;
assign v$_9899_out0 = v$_5908_out0[0:0];
assign v$_9899_out1 = v$_5908_out0[1:1];
assign v$_9900_out0 = v$_5909_out0[0:0];
assign v$_9900_out1 = v$_5909_out0[1:1];
assign v$_9903_out0 = v$_5912_out0[0:0];
assign v$_9903_out1 = v$_5912_out0[1:1];
assign v$_9905_out0 = v$_5914_out0[0:0];
assign v$_9905_out1 = v$_5914_out0[1:1];
assign v$_9906_out0 = v$_5915_out0[0:0];
assign v$_9906_out1 = v$_5915_out0[1:1];
assign v$_9909_out0 = v$_5918_out0[0:0];
assign v$_9909_out1 = v$_5918_out0[1:1];
assign v$G10_9966_out0 = ! v$LOADA_3453_out0;
assign v$G10_9967_out0 = ! v$LOADA_3454_out0;
assign v$IR2$W_10422_out0 = v$1_755_out0;
assign v$IR2$W_10423_out0 = v$1_756_out0;
assign v$G64_10577_out0 = v$G54_5642_out0 || v$G65_1383_out0;
assign v$G64_10578_out0 = v$G54_5643_out0 || v$G65_1384_out0;
assign v$RXINTERRUPT_10643_out0 = v$RXINTERRUPT_10185_out0;
assign v$RXINTERRUPT_10644_out0 = v$RXINTERRUPT_10186_out0;
assign v$EQ3_10785_out0 = v$OP_12461_out0 == 3'h7;
assign v$EQ3_10786_out0 = v$OP_12462_out0 == 3'h7;
assign v$IR2$LS_11050_out0 = v$8_10817_out0;
assign v$IR2$LS_11051_out0 = v$8_10818_out0;
assign v$G19_11223_out0 = v$EQ9_12993_out0 && v$G18_7271_out0;
assign v$G19_11224_out0 = v$EQ9_12994_out0 && v$G18_7272_out0;
assign v$G12_11404_out0 = ! v$R_6019_out0;
assign v$G12_11405_out0 = ! v$R_6020_out0;
assign v$IR1_11742_out0 = v$MUX1_10579_out0;
assign v$IR1_11743_out0 = v$MUX1_10580_out0;
assign v$MUX4_11898_out0 = v$G2_10346_out0 ? v$FF6_1525_out0 : v$_7655_out0;
assign v$MUX4_11901_out0 = v$G2_10349_out0 ? v$FF6_1528_out0 : v$_7658_out0;
assign v$MUX4_11904_out0 = v$G2_10352_out0 ? v$FF6_1531_out0 : v$_7661_out0;
assign v$MUX4_11907_out0 = v$G2_10355_out0 ? v$FF6_1534_out0 : v$_7664_out0;
assign v$IR2$P_12145_out0 = v$6_6615_out0;
assign v$IR2$P_12146_out0 = v$6_6616_out0;
assign v$E_12165_out0 = v$G2_9887_out0;
assign v$E_12166_out0 = v$G2_9888_out0;
assign v$MUX7_12681_out0 = v$G2_10346_out0 ? v$FF3_6688_out0 : v$_839_out0;
assign v$MUX7_12684_out0 = v$G2_10349_out0 ? v$FF3_6691_out0 : v$_842_out0;
assign v$MUX7_12687_out0 = v$G2_10352_out0 ? v$FF3_6694_out0 : v$_845_out0;
assign v$MUX7_12690_out0 = v$G2_10355_out0 ? v$FF3_6697_out0 : v$_848_out0;
assign v$EDGE2_12853_out0 = v$G26_6879_out0;
assign v$EDGE2_12854_out0 = v$G26_6880_out0;
assign v$IR1$RM_13011_out0 = v$SEL6_1769_out0;
assign v$IR1$RM_13012_out0 = v$SEL6_1770_out0;
assign v$IR1$FPU$OP$CODE_13016_out0 = v$SEL8_10430_out0;
assign v$IR1$FPU$OP$CODE_13017_out0 = v$SEL8_10431_out0;
assign v$G24_13080_out0 = v$G25_9422_out0 && v$G26_11205_out0;
assign v$G24_13081_out0 = v$G25_9423_out0 && v$G26_11206_out0;
assign v$G37_13137_out0 = v$Q3_13107_out0 && v$NS_12937_out0;
assign v$G37_13138_out0 = v$Q3_13108_out0 && v$NS_12938_out0;
assign v$G30_13247_out0 = v$G28_7110_out0 || v$G29_9392_out0;
assign v$G30_13248_out0 = v$G28_7111_out0 || v$G29_9393_out0;
assign v$CheckParity_13308_out0 = v$CHECKPARITY_557_out0;
assign v$CheckParity_13309_out0 = v$CHECKPARITY_558_out0;
assign v$IR2$VALID_13383_out0 = v$IR2$VALID_7594_out0;
assign v$IR2$VALID_13384_out0 = v$IR2$VALID_7595_out0;
assign v$_256_out0 = v$IR1_11742_out0[15:12];
assign v$_257_out0 = v$IR1_11743_out0[15:12];
assign v$S_406_out0 = v$S_5664_out0;
assign v$S_407_out0 = v$S_5665_out0;
assign v$IS$32$BITS_527_out0 = v$IS$32$BITS_9430_out0;
assign v$IS$32$BITS_528_out0 = v$IS$32$BITS_9431_out0;
assign v$TX_534_out0 = v$G64_10577_out0;
assign v$TX_535_out0 = v$G64_10578_out0;
assign v$EQ16_785_out0 = v$IR1$FPU$OP$CODE_13016_out0 == 2'h3;
assign v$EQ16_786_out0 = v$IR1$FPU$OP$CODE_13017_out0 == 2'h3;
assign v$_840_out0 = v$_8487_out1[0:0];
assign v$_840_out1 = v$_8487_out1[1:1];
assign v$_846_out0 = v$_8493_out1[0:0];
assign v$_846_out1 = v$_8493_out1[1:1];
assign v$RXset_891_out0 = v$RXset_3477_out0;
assign v$RXset_892_out0 = v$RXset_3478_out0;
assign v$S_1371_out0 = v$S_5664_out0;
assign v$S_1372_out0 = v$S_5665_out0;
assign v$MUX1_1489_out0 = v$G2_10344_out0 ? v$SIN_84_out0 : v$_5187_out0;
assign v$MUX1_1490_out0 = v$G2_10345_out0 ? v$SIN_85_out0 : v$_5188_out0;
assign v$MUX1_1493_out0 = v$G2_10348_out0 ? v$SIN_88_out0 : v$_5191_out0;
assign v$MUX1_1495_out0 = v$G2_10350_out0 ? v$SIN_90_out0 : v$_5193_out0;
assign v$MUX1_1496_out0 = v$G2_10351_out0 ? v$SIN_91_out0 : v$_5194_out0;
assign v$MUX1_1499_out0 = v$G2_10354_out0 ? v$SIN_94_out0 : v$_5197_out0;
assign v$G6_1891_out0 = v$G8_6485_out0 || v$G14_4141_out0;
assign v$G6_1892_out0 = v$G8_6486_out0 || v$G14_4142_out0;
assign v$EQ7_2208_out0 = v$IR2$OPCODE_1482_out0 == 4'h1;
assign v$EQ7_2209_out0 = v$IR2$OPCODE_1483_out0 == 4'h1;
assign v$MUX8_2316_out0 = v$G2_10344_out0 ? v$FF2_10133_out0 : v$_9899_out0;
assign v$MUX8_2317_out0 = v$G2_10345_out0 ? v$FF2_10134_out0 : v$_9900_out0;
assign v$MUX8_2320_out0 = v$G2_10348_out0 ? v$FF2_10137_out0 : v$_9903_out0;
assign v$MUX8_2322_out0 = v$G2_10350_out0 ? v$FF2_10139_out0 : v$_9905_out0;
assign v$MUX8_2323_out0 = v$G2_10351_out0 ? v$FF2_10140_out0 : v$_9906_out0;
assign v$MUX8_2326_out0 = v$G2_10354_out0 ? v$FF2_10143_out0 : v$_9909_out0;
assign v$XOR3_2754_out0 = v$IR2$RD_11468_out0 ^ v$IR1$RM_13011_out0;
assign v$XOR3_2755_out0 = v$IR2$RD_11469_out0 ^ v$IR1$RM_13012_out0;
assign v$G20_3698_out0 = ! v$G19_11223_out0;
assign v$G20_3699_out0 = ! v$G19_11224_out0;
assign v$ShiftEN_3842_out0 = v$RXSHIFT_388_out0;
assign v$ShiftEN_3843_out0 = v$RXSHIFT_389_out0;
assign v$G6_3951_out0 = v$_6546_out0 && v$_5720_out0;
assign v$G6_3952_out0 = v$_6547_out0 && v$_5721_out0;
assign v$G9_4233_out0 = v$EQ2_5448_out0 || v$EQ3_10785_out0;
assign v$G9_4234_out0 = v$EQ2_5449_out0 || v$EQ3_10786_out0;
assign v$MUX2_4675_out0 = v$G47_753_out0 ? v$C2_11391_out0 : v$G24_13080_out0;
assign v$MUX2_4676_out0 = v$G47_754_out0 ? v$C2_11392_out0 : v$G24_13081_out0;
assign v$IR2$VALID_5003_out0 = v$IR2$VALID_13383_out0;
assign v$IR2$VALID_5004_out0 = v$IR2$VALID_13384_out0;
assign v$_5190_out0 = v$_8487_out0[0:0];
assign v$_5190_out1 = v$_8487_out0[1:1];
assign v$_5196_out0 = v$_8493_out0[0:0];
assign v$_5196_out1 = v$_8493_out0[1:1];
assign v$_5263_out0 = v$IR1_11742_out0[11:0];
assign v$_5264_out0 = v$IR1_11743_out0[11:0];
assign v$EQ9_5486_out0 = v$IR1_11742_out0 == 16'h7000;
assign v$EQ9_5487_out0 = v$IR1_11743_out0 == 16'h7000;
assign v$G19_5745_out0 = v$SHIFTEN_4821_out0 && v$CLK4_2409_out0;
assign v$G19_5746_out0 = v$SHIFTEN_4822_out0 && v$CLK4_2410_out0;
assign v$B_5789_out0 = v$B_2417_out0;
assign v$B_5790_out0 = v$B_2418_out0;
assign v$XOR1_5800_out0 = v$IR1$RM_13011_out0 ^ v$IR2$RD_11468_out0;
assign v$XOR1_5801_out0 = v$IR1$RM_13012_out0 ^ v$IR2$RD_11469_out0;
assign v$MUX1_5804_out0 = v$C_6570_out0 ? v$C1_9650_out0 : v$SHIFT_4778_out0;
assign v$MUX1_5805_out0 = v$C_6571_out0 ? v$C1_9651_out0 : v$SHIFT_4779_out0;
assign v$S_6419_out0 = v$S_5664_out0;
assign v$S_6420_out0 = v$S_5665_out0;
assign v$MUX5_6500_out0 = v$G2_10344_out0 ? v$FF5_933_out0 : v$_5187_out1;
assign v$MUX5_6501_out0 = v$G2_10345_out0 ? v$FF5_934_out0 : v$_5188_out1;
assign v$MUX5_6504_out0 = v$G2_10348_out0 ? v$FF5_937_out0 : v$_5191_out1;
assign v$MUX5_6506_out0 = v$G2_10350_out0 ? v$FF5_939_out0 : v$_5193_out1;
assign v$MUX5_6507_out0 = v$G2_10351_out0 ? v$FF5_940_out0 : v$_5194_out1;
assign v$MUX5_6510_out0 = v$G2_10354_out0 ? v$FF5_943_out0 : v$_5197_out1;
assign v$MUX3_6670_out0 = v$G2_10344_out0 ? v$FF7_5772_out0 : v$_9899_out1;
assign v$MUX3_6671_out0 = v$G2_10345_out0 ? v$FF7_5773_out0 : v$_9900_out1;
assign v$MUX3_6674_out0 = v$G2_10348_out0 ? v$FF7_5776_out0 : v$_9903_out1;
assign v$MUX3_6676_out0 = v$G2_10350_out0 ? v$FF7_5778_out0 : v$_9905_out1;
assign v$MUX3_6677_out0 = v$G2_10351_out0 ? v$FF7_5779_out0 : v$_9906_out1;
assign v$MUX3_6680_out0 = v$G2_10354_out0 ? v$FF7_5782_out0 : v$_9909_out1;
assign v$G3_6809_out0 = ! v$E_12165_out0;
assign v$G3_6810_out0 = ! v$E_12166_out0;
assign v$MUX6_6937_out0 = v$G2_10344_out0 ? v$FF1_11255_out0 : v$_837_out1;
assign v$MUX6_6938_out0 = v$G2_10345_out0 ? v$FF1_11256_out0 : v$_838_out1;
assign v$MUX6_6941_out0 = v$G2_10348_out0 ? v$FF1_11259_out0 : v$_841_out1;
assign v$MUX6_6943_out0 = v$G2_10350_out0 ? v$FF1_11261_out0 : v$_843_out1;
assign v$MUX6_6944_out0 = v$G2_10351_out0 ? v$FF1_11262_out0 : v$_844_out1;
assign v$MUX6_6947_out0 = v$G2_10354_out0 ? v$FF1_11265_out0 : v$_847_out1;
assign v$IS$32$BIT_7152_out0 = v$IS$32$BIT_7259_out0;
assign v$IS$32$BIT_7153_out0 = v$IS$32$BIT_7260_out0;
assign v$IR2$IS$FPU_7643_out0 = v$IR2$IS$FPU_1696_out0;
assign v$IR2$IS$FPU_7644_out0 = v$IR2$IS$FPU_1697_out0;
assign v$_7656_out0 = v$_5911_out1[0:0];
assign v$_7656_out1 = v$_5911_out1[1:1];
assign v$_7662_out0 = v$_5917_out1[0:0];
assign v$_7662_out1 = v$_5917_out1[1:1];
assign v$G32_7679_out0 = !(v$G30_13247_out0 || v$G23_3040_out0);
assign v$G32_7680_out0 = !(v$G30_13248_out0 || v$G23_3041_out0);
assign v$MUX5_7734_out0 = v$STP$SAVED_5106_out0 ? v$IR1_11742_out0 : v$R_13054_out0;
assign v$MUX5_7735_out0 = v$STP$SAVED_5107_out0 ? v$IR1_11743_out0 : v$R_13055_out0;
assign v$G4_7760_out0 = ! v$_1743_out0;
assign v$G4_7761_out0 = ! v$_1744_out0;
assign v$MUX2_8006_out0 = v$_6843_out0 ? v$FF1_6867_out0 : v$_9237_out0;
assign v$MUX2_8007_out0 = v$_6844_out0 ? v$FF1_6868_out0 : v$_9238_out0;
assign v$RXINT_8180_out0 = v$RXINTERRUPT_10643_out0;
assign v$RXINT_8181_out0 = v$RXINTERRUPT_10644_out0;
assign v$ISMOV_8272_out0 = v$ISMOV_4660_out0;
assign v$ISMOV_8273_out0 = v$ISMOV_4661_out0;
assign v$S_8468_out0 = v$S_5664_out0;
assign v$S_8469_out0 = v$S_5665_out0;
assign v$EQ2_8518_out0 = v$IR1$OPCODE_6530_out0 == 4'h1;
assign v$EQ2_8519_out0 = v$IR1$OPCODE_6531_out0 == 4'h1;
assign v$EQ1_8585_out0 = v$IR1$OPCODE_6530_out0 == 4'h0;
assign v$EQ1_8586_out0 = v$IR1$OPCODE_6531_out0 == 4'h0;
assign v$IR1_8963_out0 = v$IR1_11742_out0;
assign v$IR1_8964_out0 = v$IR1_11743_out0;
assign v$NEXTSTATE_9109_out0 = v$G2_5117_out0;
assign v$MUX2_9342_out0 = v$G2_10344_out0 ? v$FF8_9843_out0 : v$_7653_out1;
assign v$MUX2_9343_out0 = v$G2_10345_out0 ? v$FF8_9844_out0 : v$_7654_out1;
assign v$MUX2_9346_out0 = v$G2_10348_out0 ? v$FF8_9847_out0 : v$_7657_out1;
assign v$MUX2_9348_out0 = v$G2_10350_out0 ? v$FF8_9849_out0 : v$_7659_out1;
assign v$MUX2_9349_out0 = v$G2_10351_out0 ? v$FF8_9850_out0 : v$_7660_out1;
assign v$MUX2_9352_out0 = v$G2_10354_out0 ? v$FF8_9853_out0 : v$_7663_out1;
assign v$G36_9492_out0 = v$G37_13137_out0 && v$G38_6823_out0;
assign v$G36_9493_out0 = v$G37_13138_out0 && v$G38_6824_out0;
assign v$_9902_out0 = v$_5911_out0[0:0];
assign v$_9902_out1 = v$_5911_out0[1:1];
assign v$_9908_out0 = v$_5917_out0[0:0];
assign v$_9908_out1 = v$_5917_out0[1:1];
assign v$G68_10489_out0 = v$G69_5702_out0 || v$G70_6845_out0;
assign v$G68_10490_out0 = v$G69_5703_out0 || v$G70_6846_out0;
assign v$EQ6_11090_out0 = v$IR2$FPU$OP_1657_out0 == 2'h3;
assign v$EQ6_11091_out0 = v$IR2$FPU$OP_1658_out0 == 2'h3;
assign v$G9_11217_out0 = ! v$IR1$C$L_6754_out0;
assign v$G9_11218_out0 = ! v$IR1$C$L_6755_out0;
assign v$G10_11578_out0 = v$E_12165_out0 && v$NQ2_11764_out0;
assign v$G10_11579_out0 = v$E_12166_out0 && v$NQ2_11765_out0;
assign v$NR_11728_out0 = v$G12_11404_out0;
assign v$NR_11729_out0 = v$G12_11405_out0;
assign v$MUX4_11896_out0 = v$G2_10344_out0 ? v$FF6_1523_out0 : v$_7653_out0;
assign v$MUX4_11897_out0 = v$G2_10345_out0 ? v$FF6_1524_out0 : v$_7654_out0;
assign v$MUX4_11900_out0 = v$G2_10348_out0 ? v$FF6_1527_out0 : v$_7657_out0;
assign v$MUX4_11902_out0 = v$G2_10350_out0 ? v$FF6_1529_out0 : v$_7659_out0;
assign v$MUX4_11903_out0 = v$G2_10351_out0 ? v$FF6_1530_out0 : v$_7660_out0;
assign v$MUX4_11906_out0 = v$G2_10354_out0 ? v$FF6_1533_out0 : v$_7663_out0;
assign v$EQ15_12096_out0 = v$IR1$OPCODE_6530_out0 == 4'h1;
assign v$EQ15_12097_out0 = v$IR1$OPCODE_6531_out0 == 4'h1;
assign v$G2_12489_out0 = ! v$C_6570_out0;
assign v$G2_12490_out0 = ! v$C_6571_out0;
assign v$MUX1_12538_out0 = v$_1554_out0 ? v$C2_6724_out0 : v$C1_11442_out0;
assign v$MUX1_12539_out0 = v$_1555_out0 ? v$C2_6725_out0 : v$C1_11443_out0;
assign v$MUX7_12679_out0 = v$G2_10344_out0 ? v$FF3_6686_out0 : v$_837_out0;
assign v$MUX7_12680_out0 = v$G2_10345_out0 ? v$FF3_6687_out0 : v$_838_out0;
assign v$MUX7_12683_out0 = v$G2_10348_out0 ? v$FF3_6690_out0 : v$_841_out0;
assign v$MUX7_12685_out0 = v$G2_10350_out0 ? v$FF3_6692_out0 : v$_843_out0;
assign v$MUX7_12686_out0 = v$G2_10351_out0 ? v$FF3_6693_out0 : v$_844_out0;
assign v$MUX7_12689_out0 = v$G2_10354_out0 ? v$FF3_6696_out0 : v$_847_out0;
assign v$G11_12785_out0 = v$G10_1683_out0 && v$CheckParity_13308_out0;
assign v$G11_12786_out0 = v$G10_1684_out0 && v$CheckParity_13309_out0;
assign v$XOR2_13161_out0 = v$IR1$RD_3732_out0 ^ v$IR2$RD_11468_out0;
assign v$XOR2_13162_out0 = v$IR1$RD_3733_out0 ^ v$IR2$RD_11469_out0;
assign v$IR1_24_out0 = v$IR1_8963_out0;
assign v$IR1_25_out0 = v$IR1_8964_out0;
assign v$G29_390_out0 = ! v$EQ16_785_out0;
assign v$G29_391_out0 = ! v$EQ16_786_out0;
assign v$_398_out0 = v$B_5789_out0[2:2];
assign v$_399_out0 = v$B_5790_out0[2:2];
assign v$G34_777_out0 = v$G35_2986_out0 || v$G36_9492_out0;
assign v$G34_778_out0 = v$G35_2987_out0 || v$G36_9493_out0;
assign v$G15_1205_out0 = v$32BIT_11086_out0 && v$IR2$IS$FPU_7643_out0;
assign v$G15_1206_out0 = v$32BIT_11087_out0 && v$IR2$IS$FPU_7644_out0;
assign v$G8_1349_out0 = ! v$G9_4233_out0;
assign v$G8_1350_out0 = ! v$G9_4234_out0;
assign v$MUX1_1492_out0 = v$G2_10347_out0 ? v$SIN_87_out0 : v$_5190_out0;
assign v$MUX1_1498_out0 = v$G2_10353_out0 ? v$SIN_93_out0 : v$_5196_out0;
assign v$NE_2135_out0 = v$G3_6809_out0;
assign v$NE_2136_out0 = v$G3_6810_out0;
assign v$RXErrorSet_2187_out0 = v$G11_12785_out0;
assign v$RXErrorSet_2188_out0 = v$G11_12786_out0;
assign v$MUX8_2319_out0 = v$G2_10347_out0 ? v$FF2_10136_out0 : v$_9902_out0;
assign v$MUX8_2325_out0 = v$G2_10353_out0 ? v$FF2_10142_out0 : v$_9908_out0;
assign v$EQ6_2668_out0 = v$XOR2_13161_out0 == 2'h0;
assign v$EQ6_2669_out0 = v$XOR2_13162_out0 == 2'h0;
assign v$ISMOV_2786_out0 = v$ISMOV_8272_out0;
assign v$ISMOV_2787_out0 = v$ISMOV_8273_out0;
assign v$EQ5_3256_out0 = v$XOR3_2754_out0 == 2'h0;
assign v$EQ5_3257_out0 = v$XOR3_2755_out0 == 2'h0;
assign v$G1_3667_out0 = v$G10_11578_out0 && v$G11_5718_out0;
assign v$G1_3668_out0 = v$G10_11579_out0 && v$G11_5719_out0;
assign v$Q1P_3774_out0 = v$MUX2_4675_out0;
assign v$Q1P_3775_out0 = v$MUX2_4676_out0;
assign v$G21_5060_out0 = v$EQ6_11090_out0 && v$IR2$FPU$L_7070_out0;
assign v$G21_5061_out0 = v$EQ6_11091_out0 && v$IR2$FPU$L_7071_out0;
assign v$INTERRUPT1_5758_out0 = v$RXINT_8180_out0;
assign v$INTERRUPT1_5759_out0 = v$RXINT_8181_out0;
assign v$ISMOV_6007_out0 = v$ISMOV_8272_out0;
assign v$ISMOV_6008_out0 = v$ISMOV_8273_out0;
assign v$MUX5_6503_out0 = v$G2_10347_out0 ? v$FF5_936_out0 : v$_5190_out1;
assign v$MUX5_6509_out0 = v$G2_10353_out0 ? v$FF5_942_out0 : v$_5196_out1;
assign v$SR_6654_out0 = v$MUX1_5804_out0;
assign v$SR_6655_out0 = v$MUX1_5805_out0;
assign v$MUX3_6673_out0 = v$G2_10347_out0 ? v$FF7_5775_out0 : v$_9902_out1;
assign v$MUX3_6679_out0 = v$G2_10353_out0 ? v$FF7_5781_out0 : v$_9908_out1;
assign v$S_6897_out0 = v$S_8468_out0;
assign v$S_6898_out0 = v$S_8469_out0;
assign v$MUX6_6940_out0 = v$G2_10347_out0 ? v$FF1_11258_out0 : v$_840_out1;
assign v$MUX6_6946_out0 = v$G2_10353_out0 ? v$FF1_11264_out0 : v$_846_out1;
assign v$_7094_out0 = v$B_5789_out0[1:1];
assign v$_7095_out0 = v$B_5790_out0[1:1];
assign v$G67_7297_out0 = v$G71_10591_out0 && v$G68_10489_out0;
assign v$G67_7298_out0 = v$G71_10592_out0 && v$G68_10490_out0;
assign v$EQUAL_7464_out0 = v$G32_7679_out0;
assign v$EQUAL_7465_out0 = v$G32_7680_out0;
assign v$TX_7506_out0 = v$TX_534_out0;
assign v$TX_7507_out0 = v$TX_535_out0;
assign v$IR1$IS$LDST_8802_out0 = v$EQ1_8585_out0;
assign v$IR1$IS$LDST_8803_out0 = v$EQ1_8586_out0;
assign v$MUX2_9345_out0 = v$G2_10347_out0 ? v$FF8_9846_out0 : v$_7656_out1;
assign v$MUX2_9351_out0 = v$G2_10353_out0 ? v$FF8_9852_out0 : v$_7662_out1;
assign v$_9711_out0 = v$B_5789_out0[3:3];
assign v$_9712_out0 = v$B_5790_out0[3:3];
assign v$N_9895_out0 = v$_5263_out0;
assign v$N_9896_out0 = v$_5264_out0;
assign v$G10_9949_out0 = v$EQ2_8518_out0 && v$EQ4_3659_out0;
assign v$G10_9950_out0 = v$EQ2_8519_out0 && v$EQ4_3660_out0;
assign v$IR2$VALID_10171_out0 = v$IR2$VALID_5003_out0;
assign v$IR2$VALID_10172_out0 = v$IR2$VALID_5004_out0;
assign v$_10441_out0 = v$B_5789_out0[0:0];
assign v$_10442_out0 = v$B_5790_out0[0:0];
assign v$EQ3_10598_out0 = v$XOR1_5800_out0 == 2'h0;
assign v$EQ3_10599_out0 = v$XOR1_5801_out0 == 2'h0;
assign v$G5_11019_out0 = ! v$IS$32$BIT_7152_out0;
assign v$G5_11020_out0 = ! v$IS$32$BIT_7153_out0;
assign v$STP$DECODED_11614_out0 = v$EQ9_5486_out0;
assign v$STP$DECODED_11615_out0 = v$EQ9_5487_out0;
assign v$MUX4_11899_out0 = v$G2_10347_out0 ? v$FF6_1526_out0 : v$_7656_out0;
assign v$MUX4_11905_out0 = v$G2_10353_out0 ? v$FF6_1532_out0 : v$_7662_out0;
assign v$S_11990_out0 = v$RXset_891_out0;
assign v$S_12001_out0 = v$RXset_892_out0;
assign v$G16_12044_out0 = v$RXset_891_out0 && v$RXlast_8470_out0;
assign v$G16_12045_out0 = v$RXset_892_out0 && v$RXlast_8471_out0;
assign v$G9_12066_out0 = v$NQ2_1741_out0 && v$NR_11728_out0;
assign v$G9_12067_out0 = v$NQ2_1742_out0 && v$NR_11729_out0;
assign v$IS$32$BITS_12390_out0 = v$IS$32$BITS_527_out0;
assign v$IS$32$BITS_12391_out0 = v$IS$32$BITS_528_out0;
assign v$OP_12599_out0 = v$_256_out0;
assign v$OP_12600_out0 = v$_257_out0;
assign v$MUX7_12682_out0 = v$G2_10347_out0 ? v$FF3_6689_out0 : v$_840_out0;
assign v$MUX7_12688_out0 = v$G2_10353_out0 ? v$FF3_6695_out0 : v$_846_out0;
assign v$S_12723_out0 = v$S_6419_out0;
assign v$S_12724_out0 = v$S_6420_out0;
assign v$G20_12991_out0 = v$NR_11728_out0 || v$Q3_12999_out0;
assign v$G20_12992_out0 = v$NR_11729_out0 || v$Q3_13000_out0;
assign v$G1_13283_out0 = v$ShiftEN_3842_out0 && v$CLK4_6074_out0;
assign v$G1_13284_out0 = v$ShiftEN_3843_out0 && v$CLK4_6075_out0;
assign v$G1_160_out0 = v$S_1371_out0 && v$ISMOV_6007_out0;
assign v$G1_161_out0 = v$S_1372_out0 && v$ISMOV_6008_out0;
assign v$G1_511_out0 = v$S_406_out0 && v$ISMOV_2786_out0;
assign v$G1_512_out0 = v$S_407_out0 && v$ISMOV_2787_out0;
assign v$G30_897_out0 = v$EQ15_12096_out0 && v$G29_390_out0;
assign v$G30_898_out0 = v$EQ15_12097_out0 && v$G29_391_out0;
assign v$G2_1355_out0 = v$EQUAL_7464_out0 && v$G3_7242_out0;
assign v$G2_1356_out0 = v$EQUAL_7465_out0 && v$G3_7243_out0;
assign v$G15_1579_out0 = v$IR1$IS$LDST_8802_out0 && v$IR1$S$WB_264_out0;
assign v$G15_1580_out0 = v$IR1$IS$LDST_8803_out0 && v$IR1$S$WB_265_out0;
assign v$IS$IR1$FMUL_1725_out0 = v$G10_9949_out0;
assign v$IS$IR1$FMUL_1726_out0 = v$G10_9950_out0;
assign v$G24_2107_out0 = v$IR1$IS$LDST_8802_out0 && v$IR1$S$WB_264_out0;
assign v$G24_2108_out0 = v$IR1$IS$LDST_8803_out0 && v$IR1$S$WB_265_out0;
assign v$IS$32$BITS_2837_out0 = v$IS$32$BITS_12390_out0;
assign v$IS$32$BITS_2838_out0 = v$IS$32$BITS_12391_out0;
assign v$SR_3024_out0 = v$SR_6654_out0;
assign v$SR_3025_out0 = v$SR_6654_out0;
assign v$SR_3026_out0 = v$SR_6654_out0;
assign v$SR_3027_out0 = v$SR_6654_out0;
assign v$SR_3028_out0 = v$SR_6655_out0;
assign v$SR_3029_out0 = v$SR_6655_out0;
assign v$SR_3030_out0 = v$SR_6655_out0;
assign v$SR_3031_out0 = v$SR_6655_out0;
assign v$OP_3431_out0 = v$OP_12599_out0;
assign v$OP_3432_out0 = v$OP_12600_out0;
assign v$G33_3506_out0 = v$NQ2_13211_out0 && v$G34_777_out0;
assign v$G33_3507_out0 = v$NQ2_13212_out0 && v$G34_778_out0;
assign v$IR2$VALID_4452_out0 = v$IR2$VALID_10171_out0;
assign v$IR2$VALID_4453_out0 = v$IR2$VALID_10172_out0;
assign v$G1_4923_out0 = v$G2_12489_out0 && v$_10441_out0;
assign v$G1_4924_out0 = v$G2_12490_out0 && v$_10442_out0;
assign v$IR1_5151_out0 = v$IR1_24_out0;
assign v$IR1_5152_out0 = v$IR1_25_out0;
assign v$G18_5876_out0 = v$G20_12991_out0 && v$G19_1347_out0;
assign v$G18_5877_out0 = v$G20_12992_out0 && v$G19_1348_out0;
assign v$G11_6564_out0 = v$EQ6_2668_out0 || v$EQ5_3256_out0;
assign v$G11_6565_out0 = v$EQ6_2669_out0 || v$EQ5_3257_out0;
assign v$Shift_6566_out0 = v$G1_13283_out0;
assign v$Shift_6567_out0 = v$G1_13284_out0;
assign v$EXEC2_6611_out0 = v$IR2$VALID_10171_out0;
assign v$EXEC2_6612_out0 = v$IR2$VALID_10172_out0;
assign v$IR2$VALID_6998_out0 = v$IR2$VALID_10171_out0;
assign v$IR2$VALID_6999_out0 = v$IR2$VALID_10172_out0;
assign v$G8_7301_out0 = v$Q1_7197_out0 && v$G9_12066_out0;
assign v$G8_7302_out0 = v$Q1_7198_out0 && v$G9_12067_out0;
assign v$G13_7935_out0 = v$G14_13117_out0 && v$NE_2135_out0;
assign v$G13_7936_out0 = v$G14_13118_out0 && v$NE_2136_out0;
assign v$ERR_8428_out0 = v$RXErrorSet_2187_out0;
assign v$ERR_8429_out0 = v$RXErrorSet_2188_out0;
assign v$G15_9165_out0 = v$NE_2135_out0 && v$G16_1783_out0;
assign v$G15_9166_out0 = v$NE_2136_out0 && v$G16_1784_out0;
assign v$G25_10025_out0 = v$G21_5060_out0 && v$EQ7_2208_out0;
assign v$G25_10026_out0 = v$G21_5061_out0 && v$EQ7_2209_out0;
assign v$G4_10044_out0 = v$NE_2135_out0 && v$G5_7012_out0;
assign v$G4_10045_out0 = v$NE_2136_out0 && v$G5_7013_out0;
assign v$G17_10145_out0 = v$IR2$VALID_10171_out0 && v$G20_3698_out0;
assign v$G17_10146_out0 = v$IR2$VALID_10172_out0 && v$G20_3699_out0;
assign v$N_10183_out0 = v$N_9895_out0;
assign v$N_10184_out0 = v$N_9896_out0;
assign v$EQUAL_11046_out0 = v$EQUAL_7464_out0;
assign v$EQUAL_11047_out0 = v$EQUAL_7465_out0;
assign v$EXEC2_11098_out0 = v$IR2$VALID_10171_out0;
assign v$EXEC2_11099_out0 = v$IR2$VALID_10172_out0;
assign v$TXRST_11484_out0 = v$G67_7297_out0;
assign v$TXRST_11485_out0 = v$G67_7298_out0;
assign v$EN_11491_out0 = v$_7094_out0;
assign v$EN_11492_out0 = v$_398_out0;
assign v$EN_11493_out0 = v$_9711_out0;
assign v$EN_11495_out0 = v$_7095_out0;
assign v$EN_11496_out0 = v$_399_out0;
assign v$EN_11497_out0 = v$_9712_out0;
assign v$S_11992_out0 = v$G16_12044_out0;
assign v$S_12003_out0 = v$G16_12045_out0;
assign v$G16_12037_out0 = v$EQ3_10598_out0 && v$IR1$IS$LDST_8802_out0;
assign v$G16_12038_out0 = v$EQ3_10599_out0 && v$IR1$IS$LDST_8803_out0;
assign v$G14_12092_out0 = v$IR1$IS$LDST_8802_out0 && v$G9_11217_out0;
assign v$G14_12093_out0 = v$IR1$IS$LDST_8803_out0 && v$G9_11218_out0;
assign v$G36_12163_out0 = ! v$STP$DECODED_11614_out0;
assign v$G36_12164_out0 = ! v$STP$DECODED_11615_out0;
assign v$EDGE1_12216_out0 = v$INTERRUPT1_5758_out0;
assign v$EDGE1_12217_out0 = v$INTERRUPT1_5759_out0;
assign v$EXEC2_358_out0 = v$EXEC2_11098_out0;
assign v$EXEC2_359_out0 = v$EXEC2_11099_out0;
assign v$IR1$IS$FPU$ARITHMETIC_595_out0 = v$G30_897_out0;
assign v$IR1$IS$FPU$ARITHMETIC_596_out0 = v$G30_898_out0;
assign v$G1_1066_out0 = v$EXEC2_11098_out0 && v$IR15_7240_out0;
assign v$G1_1067_out0 = v$EXEC2_11099_out0 && v$IR15_7241_out0;
assign v$EXEC2_1091_out0 = v$EXEC2_6611_out0;
assign v$EXEC2_1092_out0 = v$EXEC2_6612_out0;
assign v$G12_1148_out0 = v$G13_7935_out0 || v$G15_9165_out0;
assign v$G12_1149_out0 = v$G13_7936_out0 || v$G15_9166_out0;
assign v$G3_1369_out0 = v$G15_1579_out0 && v$IS$IR2$DATA$PROCESSING_6664_out0;
assign v$G3_1370_out0 = v$G15_1580_out0 && v$IS$IR2$DATA$PROCESSING_6665_out0;
assign v$G29_2332_out0 = v$G30_1389_out0 || v$G33_3506_out0;
assign v$G29_2333_out0 = v$G30_1390_out0 || v$G33_3507_out0;
assign v$G3_2658_out0 = v$G8_7301_out0 || v$G10_12927_out0;
assign v$G3_2659_out0 = v$G8_7302_out0 || v$G10_12928_out0;
assign v$SEL1_3611_out0 = v$IR1_5151_out0[9:8];
assign v$SEL1_3612_out0 = v$IR1_5152_out0[9:8];
assign v$G12_4181_out0 = v$IS$IR1$FMUL_1725_out0 && v$G11_6564_out0;
assign v$G12_4182_out0 = v$IS$IR1$FMUL_1726_out0 && v$G11_6565_out0;
assign v$_4200_out0 = v$IR1_5151_out0[1:0];
assign v$_4201_out0 = v$IR1_5152_out0[1:0];
assign v$IR2$VALID$AND$NOT$FLOAD_4883_out0 = v$G17_10145_out0;
assign v$IR2$VALID$AND$NOT$FLOAD_4884_out0 = v$G17_10146_out0;
assign v$TXRST_5553_out0 = v$TXRST_11484_out0;
assign v$TXRST_5554_out0 = v$TXRST_11485_out0;
assign v$N_5753_out0 = v$N_10183_out0;
assign v$N_5754_out0 = v$N_10184_out0;
assign v$S_6988_out0 = v$G1_511_out0;
assign v$S_6989_out0 = v$G1_512_out0;
assign v$S_7016_out0 = v$G1_160_out0;
assign v$S_7017_out0 = v$G1_161_out0;
assign v$N_7740_out0 = v$N_10183_out0;
assign v$N_7741_out0 = v$N_10184_out0;
assign v$_8426_out0 = v$IR1_5151_out0[15:15];
assign v$_8427_out0 = v$IR1_5152_out0[15:15];
assign v$G26_8786_out0 = v$G24_2107_out0 && v$G25_1387_out0;
assign v$G26_8787_out0 = v$G24_2108_out0 && v$G25_1388_out0;
assign v$IR2$VALID_8838_out0 = v$IR2$VALID_4452_out0;
assign v$IR2$VALID_8839_out0 = v$IR2$VALID_4453_out0;
assign v$_9112_out0 = v$IR1_5151_out0[8:8];
assign v$_9113_out0 = v$IR1_5152_out0[8:8];
assign v$G23_9472_out0 = ! v$G25_10025_out0;
assign v$G23_9473_out0 = ! v$G25_10026_out0;
assign v$OP_10131_out0 = v$OP_3431_out0;
assign v$OP_10132_out0 = v$OP_3432_out0;
assign v$COUNTERINTERRUPT_10189_out0 = v$G2_1355_out0;
assign v$COUNTERINTERRUPT_10190_out0 = v$G2_1356_out0;
assign v$IR2$VALID_11092_out0 = v$IR2$VALID_6998_out0;
assign v$IR2$VALID_11093_out0 = v$IR2$VALID_6999_out0;
assign v$_11128_out0 = v$IR1_5151_out0[11:10];
assign v$_11129_out0 = v$IR1_5152_out0[11:10];
assign v$EN_11490_out0 = v$G1_4923_out0;
assign v$EN_11494_out0 = v$G1_4924_out0;
assign v$_11744_out0 = v$IR1_5151_out0[14:12];
assign v$_11745_out0 = v$IR1_5152_out0[14:12];
assign v$SR_11838_out0 = v$SR_3024_out0;
assign v$SR_11839_out0 = v$SR_3025_out0;
assign v$SR_11840_out0 = v$SR_3026_out0;
assign v$SR_11841_out0 = v$SR_3027_out0;
assign v$SR_11842_out0 = v$SR_3028_out0;
assign v$SR_11843_out0 = v$SR_3029_out0;
assign v$SR_11844_out0 = v$SR_3030_out0;
assign v$SR_11845_out0 = v$SR_3031_out0;
assign v$EN_12030_out0 = v$EN_11491_out0;
assign v$EN_12031_out0 = v$EN_11492_out0;
assign v$EN_12032_out0 = v$EN_11493_out0;
assign v$EN_12034_out0 = v$EN_11495_out0;
assign v$EN_12035_out0 = v$EN_11496_out0;
assign v$EN_12036_out0 = v$EN_11497_out0;
assign v$INTERRUPT1_12516_out0 = v$EDGE1_12216_out0;
assign v$INTERRUPT1_12517_out0 = v$EDGE1_12217_out0;
assign v$G15_12619_out0 = v$G17_7508_out0 || v$G18_5876_out0;
assign v$G15_12620_out0 = v$G17_7509_out0 || v$G18_5877_out0;
assign v$IR1_12803_out0 = v$IR1_5151_out0;
assign v$IR1_12804_out0 = v$IR1_5152_out0;
assign v$IR1_370_out0 = v$IR1_12803_out0;
assign v$IR1_371_out0 = v$IR1_12804_out0;
assign v$G31_997_out0 = v$G28_10029_out0 && v$IR1$IS$FPU$ARITHMETIC_595_out0;
assign v$G31_998_out0 = v$G28_10030_out0 && v$IR1$IS$FPU$ARITHMETIC_596_out0;
assign v$SEL2_1361_out0 = v$IR1_12803_out0[15:12];
assign v$SEL2_1362_out0 = v$IR1_12804_out0[15:12];
assign v$EQ1_1585_out0 = v$SR_11839_out0 == 2'h1;
assign v$EQ1_1586_out0 = v$SR_11843_out0 == 2'h1;
assign v$EQ2_1923_out0 = v$SR_11841_out0 == 2'h2;
assign v$EQ2_1924_out0 = v$SR_11845_out0 == 2'h2;
assign v$G18_2105_out0 = v$INTERRUPT1_12516_out0 && v$G17_3720_out0;
assign v$G18_2106_out0 = v$INTERRUPT1_12517_out0 && v$G17_3721_out0;
assign v$TXINTERRUPT_2342_out0 = v$TXRST_5553_out0;
assign v$TXINTERRUPT_2343_out0 = v$TXRST_5554_out0;
assign v$IR1$FPU$OP_2545_out0 = v$SEL1_3611_out0;
assign v$IR1$FPU$OP_2546_out0 = v$SEL1_3612_out0;
assign v$IR1$D_2900_out0 = v$_11128_out0;
assign v$IR1$D_2901_out0 = v$_11129_out0;
assign v$G2_3435_out0 = v$Q3_12999_out0 && v$G3_2658_out0;
assign v$G2_3436_out0 = v$Q3_13000_out0 && v$G3_2659_out0;
assign v$EQ1_3449_out0 = v$SR_11840_out0 == 2'h1;
assign v$EQ1_3450_out0 = v$SR_11844_out0 == 2'h1;
assign v$EQ1_3457_out0 = v$SR_11838_out0 == 2'h3;
assign v$EQ1_3458_out0 = v$SR_11842_out0 == 2'h3;
assign v$G14_3629_out0 = v$G16_4419_out0 || v$G15_12619_out0;
assign v$G14_3630_out0 = v$G16_4420_out0 || v$G15_12620_out0;
assign v$EQ3_3683_out0 = v$SR_11840_out0 == 2'h3;
assign v$EQ3_3684_out0 = v$SR_11844_out0 == 2'h3;
assign v$IR1$OP_3762_out0 = v$_11744_out0;
assign v$IR1$OP_3763_out0 = v$_11745_out0;
assign v$IR1$15_3786_out0 = v$_8426_out0;
assign v$IR1$15_3787_out0 = v$_8427_out0;
assign v$MUX3_4145_out0 = v$G47_753_out0 ? v$C3_13205_out0 : v$G29_2332_out0;
assign v$MUX3_4146_out0 = v$G47_754_out0 ? v$C3_13206_out0 : v$G29_2333_out0;
assign v$G4_5100_out0 = v$G3_1369_out0 || v$G16_12037_out0;
assign v$G4_5101_out0 = v$G3_1370_out0 || v$G16_12038_out0;
assign v$IR1$S_5370_out0 = v$_9112_out0;
assign v$IR1$S_5371_out0 = v$_9113_out0;
assign v$EQ3_5414_out0 = v$SR_11838_out0 == 2'h1;
assign v$EQ3_5415_out0 = v$SR_11842_out0 == 2'h1;
assign v$EQ1_6960_out0 = v$SR_11841_out0 == 2'h3;
assign v$EQ1_6961_out0 = v$SR_11845_out0 == 2'h3;
assign v$OP_7246_out0 = v$OP_10131_out0;
assign v$OP_7247_out0 = v$OP_10132_out0;
assign v$_7572_out0 = { v$N_7740_out0,v$C1_3657_out0 };
assign v$_7573_out0 = { v$N_7741_out0,v$C1_3658_out0 };
assign v$G6_7724_out0 = v$IR2$VALID_8838_out0 && v$IR2$L_8105_out0;
assign v$G6_7725_out0 = v$IR2$VALID_8839_out0 && v$IR2$L_8106_out0;
assign v$EQ3_7911_out0 = v$SR_11841_out0 == 2'h1;
assign v$EQ3_7912_out0 = v$SR_11845_out0 == 2'h1;
assign v$IR1$M_8836_out0 = v$_4200_out0;
assign v$IR1$M_8837_out0 = v$_4201_out0;
assign v$G7_9129_out0 = v$G1_1066_out0 && v$G8_1349_out0;
assign v$G7_9130_out0 = v$G1_1067_out0 && v$G8_1350_out0;
assign v$EQ2_9180_out0 = v$SR_11839_out0 == 2'h2;
assign v$EQ2_9181_out0 = v$SR_11843_out0 == 2'h2;
assign v$EQ2_9691_out0 = v$SR_11838_out0 == 2'h2;
assign v$EQ2_9692_out0 = v$SR_11842_out0 == 2'h2;
assign v$G14_10042_out0 = ! v$INTERRUPT1_12516_out0;
assign v$G14_10043_out0 = ! v$INTERRUPT1_12517_out0;
assign v$EXEC2_11473_out0 = v$EXEC2_1091_out0;
assign v$EXEC2_11474_out0 = v$EXEC2_1092_out0;
assign v$EQ2_11498_out0 = v$SR_11840_out0 == 2'h2;
assign v$EQ2_11499_out0 = v$SR_11844_out0 == 2'h2;
assign v$G32_11512_out0 = v$INTERRUPT3_2210_out0 || v$COUNTERINTERRUPT_10189_out0;
assign v$G32_11513_out0 = v$INTERRUPT3_2211_out0 || v$COUNTERINTERRUPT_10190_out0;
assign v$EQ3_11624_out0 = v$SR_11839_out0 == 2'h3;
assign v$EQ3_11625_out0 = v$SR_11843_out0 == 2'h3;
assign v$EN_12029_out0 = v$EN_11490_out0;
assign v$EN_12033_out0 = v$EN_11494_out0;
assign v$TXReset_12625_out0 = v$TXRST_5553_out0;
assign v$TXReset_12626_out0 = v$TXRST_5554_out0;
assign v$G24_12707_out0 = v$IR2$VALID_8838_out0 && v$G23_9472_out0;
assign v$G24_12708_out0 = v$IR2$VALID_8839_out0 && v$G23_9473_out0;
assign v$N_13005_out0 = v$N_5753_out0;
assign v$N_13006_out0 = v$N_5754_out0;
assign v$G21_13310_out0 = v$IR2$VALID$AND$NOT$FLOAD_4883_out0 && v$EQ11_7677_out0;
assign v$G21_13311_out0 = v$IR2$VALID$AND$NOT$FLOAD_4884_out0 && v$EQ11_7678_out0;
assign v$N_825_out0 = v$N_13005_out0;
assign v$N_826_out0 = v$N_13006_out0;
assign v$G8_1036_out0 = v$EQ1_3457_out0 && v$EN_12029_out0;
assign v$G8_1037_out0 = v$EQ3_11624_out0 && v$EN_12030_out0;
assign v$G8_1038_out0 = v$EQ3_3683_out0 && v$EN_12031_out0;
assign v$G8_1039_out0 = v$EQ1_6960_out0 && v$EN_12032_out0;
assign v$G8_1040_out0 = v$EQ1_3458_out0 && v$EN_12033_out0;
assign v$G8_1041_out0 = v$EQ3_11625_out0 && v$EN_12034_out0;
assign v$G8_1042_out0 = v$EQ3_3684_out0 && v$EN_12035_out0;
assign v$G8_1043_out0 = v$EQ1_6961_out0 && v$EN_12036_out0;
assign v$NEXTENDED_1060_out0 = v$_7572_out0;
assign v$NEXTENDED_1061_out0 = v$_7573_out0;
assign v$G3_1507_out0 = v$EQ3_5414_out0 && v$EN_12029_out0;
assign v$G3_1508_out0 = v$EQ1_1585_out0 && v$EN_12030_out0;
assign v$G3_1509_out0 = v$EQ1_3449_out0 && v$EN_12031_out0;
assign v$G3_1510_out0 = v$EQ3_7911_out0 && v$EN_12032_out0;
assign v$G3_1511_out0 = v$EQ3_5415_out0 && v$EN_12033_out0;
assign v$G3_1512_out0 = v$EQ1_1586_out0 && v$EN_12034_out0;
assign v$G3_1513_out0 = v$EQ1_3450_out0 && v$EN_12035_out0;
assign v$G3_1514_out0 = v$EQ3_7912_out0 && v$EN_12036_out0;
assign v$MUX2_1661_out0 = v$IR2$VALID$AND$NOT$FLOAD_4883_out0 ? v$IR2$D_9879_out0 : v$IR1$M_8836_out0;
assign v$MUX2_1662_out0 = v$IR2$VALID$AND$NOT$FLOAD_4884_out0 ? v$IR2$D_9880_out0 : v$IR1$M_8837_out0;
assign v$OP_2405_out0 = v$OP_7246_out0;
assign v$OP_2406_out0 = v$OP_7247_out0;
assign v$EXEC2_2720_out0 = v$EXEC2_11473_out0;
assign v$EXEC2_2721_out0 = v$EXEC2_11474_out0;
assign v$G4_2746_out0 = v$EQ2_9691_out0 && v$EN_12029_out0;
assign v$G4_2747_out0 = v$EQ2_9180_out0 && v$EN_12030_out0;
assign v$G4_2748_out0 = v$EQ2_11498_out0 && v$EN_12031_out0;
assign v$G4_2749_out0 = v$EQ2_1923_out0 && v$EN_12032_out0;
assign v$G4_2750_out0 = v$EQ2_9692_out0 && v$EN_12033_out0;
assign v$G4_2751_out0 = v$EQ2_9181_out0 && v$EN_12034_out0;
assign v$G4_2752_out0 = v$EQ2_11499_out0 && v$EN_12035_out0;
assign v$G4_2753_out0 = v$EQ2_1924_out0 && v$EN_12036_out0;
assign v$EXEC2_3042_out0 = v$EXEC2_11473_out0;
assign v$EXEC2_3043_out0 = v$EXEC2_11474_out0;
assign v$G16_3103_out0 = v$FF2_11724_out0 && v$G14_10042_out0;
assign v$G16_3104_out0 = v$FF2_11725_out0 && v$G14_10043_out0;
assign v$TXINT_3304_out0 = v$TXINTERRUPT_2342_out0;
assign v$TXINT_3305_out0 = v$TXINTERRUPT_2343_out0;
assign v$Q2P_4041_out0 = v$MUX3_4145_out0;
assign v$Q2P_4042_out0 = v$MUX3_4146_out0;
assign v$G8_4071_out0 = v$G4_5100_out0 || v$G14_12092_out0;
assign v$G8_4072_out0 = v$G4_5101_out0 || v$G14_12093_out0;
assign v$EQ3_4843_out0 = v$IR1$FPU$OP_2545_out0 == 2'h2;
assign v$EQ3_4844_out0 = v$IR1$FPU$OP_2546_out0 == 2'h2;
assign v$EXEC2_5520_out0 = v$EXEC2_11473_out0;
assign v$EXEC2_5521_out0 = v$EXEC2_11474_out0;
assign v$S_8290_out0 = v$IR1$S_5370_out0;
assign v$S_8291_out0 = v$IR1$S_5371_out0;
assign v$G15_8965_out0 = v$G18_2105_out0 && v$R1_10327_out0;
assign v$G15_8966_out0 = v$G18_2106_out0 && v$R1_10328_out0;
assign v$INT3_9426_out0 = v$G32_11512_out0;
assign v$INT3_9427_out0 = v$G32_11513_out0;
assign v$G13_10418_out0 = v$NQ0_5322_out0 && v$G14_3629_out0;
assign v$G13_10419_out0 = v$NQ0_5323_out0 && v$G14_3630_out0;
assign v$G4_11042_out0 = ! v$IR1$15_3786_out0;
assign v$G4_11043_out0 = ! v$IR1$15_3787_out0;
assign v$IR1_11186_out0 = v$IR1_370_out0;
assign v$IR1_11187_out0 = v$IR1_371_out0;
assign v$EQ4_11584_out0 = v$IR1$FPU$OP_2545_out0 == 2'h2;
assign v$EQ4_11585_out0 = v$IR1$FPU$OP_2546_out0 == 2'h2;
assign v$IR1$FULL$OP$CODE_12104_out0 = v$SEL2_1361_out0;
assign v$IR1$FULL$OP$CODE_12105_out0 = v$SEL2_1362_out0;
assign v$EXEC2_12457_out0 = v$EXEC2_11473_out0;
assign v$EXEC2_12458_out0 = v$EXEC2_11474_out0;
assign v$N_12713_out0 = v$N_13005_out0;
assign v$N_12714_out0 = v$N_13006_out0;
assign v$R_13038_out0 = v$TXReset_12625_out0;
assign v$R_13049_out0 = v$TXReset_12626_out0;
assign v$WENALU_13296_out0 = v$G7_9129_out0;
assign v$WENALU_13297_out0 = v$G7_9130_out0;
assign v$_38_out0 = v$IR1_11186_out0[8:8];
assign v$_39_out0 = v$IR1_11187_out0[8:8];
assign v$EQ8_217_out0 = v$IR1$FULL$OP$CODE_12104_out0 == 4'h0;
assign v$EQ8_218_out0 = v$IR1$FULL$OP$CODE_12105_out0 == 4'h0;
assign v$_414_out0 = v$IR1_11186_out0[11:10];
assign v$_415_out0 = v$IR1_11187_out0[11:10];
assign v$EXEC2_461_out0 = v$EXEC2_3042_out0;
assign v$EXEC2_462_out0 = v$EXEC2_3043_out0;
assign v$EXEC2_701_out0 = v$EXEC2_5520_out0;
assign v$EXEC2_702_out0 = v$EXEC2_5521_out0;
assign v$EQ5_733_out0 = v$IR1$FULL$OP$CODE_12104_out0 == 4'h1;
assign v$EQ5_734_out0 = v$IR1$FULL$OP$CODE_12105_out0 == 4'h1;
assign v$INTERRUPT0_979_out0 = v$TXINT_3304_out0;
assign v$INTERRUPT0_980_out0 = v$TXINT_3305_out0;
assign v$_1009_out0 = v$IR1_11186_out0[5:2];
assign v$_1010_out0 = v$IR1_11187_out0[5:2];
assign v$EQ5_1062_out0 = v$OP_2405_out0 == 4'h6;
assign v$EQ5_1063_out0 = v$OP_2406_out0 == 4'h6;
assign v$_1108_out0 = v$IR1_11186_out0[6:6];
assign v$_1109_out0 = v$IR1_11187_out0[6:6];
assign v$EDGE3_1168_out0 = v$INT3_9426_out0;
assign v$EDGE3_1169_out0 = v$INT3_9427_out0;
assign v$_1375_out0 = v$IR1_11186_out0[9:9];
assign v$_1376_out0 = v$IR1_11187_out0[9:9];
assign v$_1571_out0 = { v$Q2P_4041_out0,v$Q3P_7500_out0 };
assign v$_1572_out0 = { v$Q2P_4042_out0,v$Q3P_7501_out0 };
assign v$WENALU_2782_out0 = v$WENALU_13296_out0;
assign v$WENALU_2783_out0 = v$WENALU_13297_out0;
assign v$EQ1_2809_out0 = v$OP_2405_out0 == 4'h2;
assign v$EQ1_2810_out0 = v$OP_2406_out0 == 4'h2;
assign v$EQ3_3768_out0 = v$OP_2405_out0 == 4'h4;
assign v$EQ3_3769_out0 = v$OP_2406_out0 == 4'h4;
assign v$_4887_out0 = v$IR1_11186_out0[7:7];
assign v$_4888_out0 = v$IR1_11187_out0[7:7];
assign v$EXEC2_5557_out0 = v$EXEC2_12457_out0;
assign v$EXEC2_5558_out0 = v$EXEC2_12458_out0;
assign v$EQ13_6370_out0 = v$IR1$FULL$OP$CODE_12104_out0 == 4'h1;
assign v$EQ13_6371_out0 = v$IR1$FULL$OP$CODE_12105_out0 == 4'h1;
assign v$EQ4_6379_out0 = v$OP_2405_out0 == 4'h5;
assign v$EQ4_6380_out0 = v$OP_2406_out0 == 4'h5;
assign v$EXEC2_6435_out0 = v$EXEC2_2720_out0;
assign v$EXEC2_6436_out0 = v$EXEC2_2721_out0;
assign v$_7098_out0 = v$IR1_11186_out0[1:0];
assign v$_7099_out0 = v$IR1_11187_out0[1:0];
assign v$EQ2_7104_out0 = v$OP_2405_out0 == 4'h3;
assign v$EQ2_7105_out0 = v$OP_2406_out0 == 4'h3;
assign v$N_7568_out0 = v$N_12713_out0;
assign v$N_7569_out0 = v$N_12714_out0;
assign v$EQ14_7897_out0 = v$IR1$FULL$OP$CODE_12104_out0 == 4'h1;
assign v$EQ14_7898_out0 = v$IR1$FULL$OP$CODE_12105_out0 == 4'h1;
assign v$_8418_out0 = v$IR1_11186_out0[15:15];
assign v$_8419_out0 = v$IR1_11187_out0[15:15];
assign v$NEXTENDED_9754_out0 = v$NEXTENDED_1060_out0;
assign v$NEXTENDED_9755_out0 = v$NEXTENDED_1061_out0;
assign v$G13_10192_out0 = v$G8_4071_out0 || v$G12_4181_out0;
assign v$G13_10193_out0 = v$G8_4072_out0 || v$G12_4182_out0;
assign v$AD3_10447_out0 = v$MUX2_1661_out0;
assign v$AD3_10448_out0 = v$MUX2_1662_out0;
assign v$G1_10609_out0 = v$G2_3435_out0 || v$G13_10418_out0;
assign v$G1_10610_out0 = v$G2_3436_out0 || v$G13_10419_out0;
assign v$G6_10839_out0 = ! v$R_13038_out0;
assign v$G6_10850_out0 = ! v$R_13049_out0;
assign v$EQ2_11025_out0 = v$IR1_11186_out0 == 16'h7000;
assign v$EQ2_11026_out0 = v$IR1_11187_out0 == 16'h7000;
assign v$_11221_out0 = v$IR1_11186_out0[15:12];
assign v$_11222_out0 = v$IR1_11187_out0[15:12];
assign v$EQ6_11402_out0 = v$OP_2405_out0 == 4'h7;
assign v$EQ6_11403_out0 = v$OP_2406_out0 == 4'h7;
assign v$S_11488_out0 = v$S_8290_out0;
assign v$S_11489_out0 = v$S_8291_out0;
assign v$G13_11612_out0 = v$G16_3103_out0 && v$F1_2195_out0;
assign v$G13_11613_out0 = v$G16_3104_out0 && v$F1_2196_out0;
assign v$END_11670_out0 = v$N_825_out0;
assign v$END_11671_out0 = v$N_826_out0;
assign v$JMI_72_out0 = v$EQ4_6379_out0;
assign v$JMI_73_out0 = v$EQ4_6380_out0;
assign v$G5_423_out0 = v$FF2_8668_out0 && v$G6_10839_out0;
assign v$G5_428_out0 = v$FF2_8679_out0 && v$G6_10850_out0;
assign v$JMP_861_out0 = v$EQ3_3768_out0;
assign v$JMP_862_out0 = v$EQ3_3769_out0;
assign v$JLS_1096_out0 = v$EQ2_7104_out0;
assign v$JLS_1097_out0 = v$EQ2_7105_out0;
assign v$INTERRUPT3_1583_out0 = v$EDGE3_1168_out0;
assign v$INTERRUPT3_1584_out0 = v$EDGE3_1169_out0;
assign v$IR1$OPCODE_1671_out0 = v$_11221_out0;
assign v$IR1$OPCODE_1672_out0 = v$_11222_out0;
assign v$G25_2250_out0 = ! v$EQ14_7897_out0;
assign v$G25_2251_out0 = ! v$EQ14_7898_out0;
assign v$IR1$P_2407_out0 = v$_4887_out0;
assign v$IR1$P_2408_out0 = v$_4888_out0;
assign v$IR1$L_3512_out0 = v$_1375_out0;
assign v$IR1$L_3513_out0 = v$_1376_out0;
assign v$EDGE0_3772_out0 = v$INTERRUPT0_979_out0;
assign v$EDGE0_3773_out0 = v$INTERRUPT0_980_out0;
assign v$STP_4222_out0 = v$EQ6_11402_out0;
assign v$STP_4223_out0 = v$EQ6_11403_out0;
assign v$STOP$1_5336_out0 = v$EQ2_11025_out0;
assign v$STOP$1_5337_out0 = v$EQ2_11026_out0;
assign v$Q0P_7944_out0 = v$G1_10609_out0;
assign v$Q0P_7945_out0 = v$G1_10610_out0;
assign v$IR1$M_8274_out0 = v$_7098_out0;
assign v$IR1$M_8275_out0 = v$_7099_out0;
assign v$AD3_8756_out0 = v$AD3_10447_out0;
assign v$AD3_8757_out0 = v$AD3_10448_out0;
assign v$EQ10_8978_out0 = v$N_7568_out0 == 12'h2;
assign v$EQ10_8979_out0 = v$N_7569_out0 == 12'h2;
assign v$EQ11_9167_out0 = v$N_7568_out0 == 12'h4;
assign v$EQ11_9168_out0 = v$N_7569_out0 == 12'h4;
assign v$EQ8_9715_out0 = v$N_7568_out0 == 12'h0;
assign v$EQ8_9716_out0 = v$N_7569_out0 == 12'h0;
assign v$IR1$U_10127_out0 = v$_1108_out0;
assign v$IR1$U_10128_out0 = v$_1109_out0;
assign v$IR1$D_10187_out0 = v$_414_out0;
assign v$IR1$D_10188_out0 = v$_415_out0;
assign v$JLO_10309_out0 = v$EQ1_2809_out0;
assign v$JLO_10310_out0 = v$EQ1_2810_out0;
assign v$G22_10900_out0 = v$EQ4_11584_out0 && v$EQ13_6370_out0;
assign v$G22_10901_out0 = v$EQ4_11585_out0 && v$EQ13_6371_out0;
assign v$IR1$N_11003_out0 = v$_1009_out0;
assign v$IR1$N_11004_out0 = v$_1010_out0;
assign v$IR1$LS_11519_out0 = v$_8418_out0;
assign v$IR1$LS_11520_out0 = v$_8419_out0;
assign v$IR1$W_11628_out0 = v$_38_out0;
assign v$IR1$W_11629_out0 = v$_39_out0;
assign v$G5_11636_out0 = v$EQ3_4843_out0 && v$EQ5_733_out0;
assign v$G5_11637_out0 = v$EQ3_4844_out0 && v$EQ5_734_out0;
assign v$G19_11762_out0 = v$G15_8965_out0 || v$G13_11612_out0;
assign v$G19_11763_out0 = v$G15_8966_out0 || v$G13_11613_out0;
assign v$G23_11817_out0 = v$G13_10192_out0 || v$G26_8786_out0;
assign v$G23_11818_out0 = v$G13_10193_out0 || v$G26_8787_out0;
assign v$EQ7_11947_out0 = v$N_7568_out0 == 12'h1;
assign v$EQ7_11948_out0 = v$N_7569_out0 == 12'h1;
assign v$G2_12108_out0 = v$S_11488_out0 && v$EXEC2_358_out0;
assign v$G2_12109_out0 = v$S_11489_out0 && v$EXEC2_359_out0;
assign v$EQ9_12558_out0 = v$N_7568_out0 == 12'h3;
assign v$EQ9_12559_out0 = v$N_7569_out0 == 12'h3;
assign v$JEQ_12805_out0 = v$EQ5_1062_out0;
assign v$JEQ_12806_out0 = v$EQ5_1063_out0;
assign v$EQ13_13201_out0 = v$N_7568_out0 == 12'h5;
assign v$EQ13_13202_out0 = v$N_7569_out0 == 12'h5;
assign v$JEQ_869_out0 = v$JEQ_12805_out0;
assign v$JEQ_870_out0 = v$JEQ_12806_out0;
assign v$G32_1001_out0 = v$INTERRUPT3_1583_out0 && v$G31_6588_out0;
assign v$G32_1002_out0 = v$INTERRUPT3_1584_out0 && v$G31_6589_out0;
assign v$G3_1573_out0 = v$G2_12108_out0 && v$G4_7760_out0;
assign v$G3_1574_out0 = v$G2_12109_out0 && v$G4_7761_out0;
assign v$G28_1895_out0 = ! v$INTERRUPT3_1583_out0;
assign v$G28_1896_out0 = ! v$INTERRUPT3_1584_out0;
assign v$JMP_2998_out0 = v$JMP_861_out0;
assign v$JMP_2999_out0 = v$JMP_862_out0;
assign v$_3459_out0 = { v$Q0P_7944_out0,v$Q1P_7261_out0 };
assign v$_3460_out0 = { v$Q0P_7945_out0,v$Q1P_7262_out0 };
assign v$JLO_5611_out0 = v$JLO_10309_out0;
assign v$JLO_5612_out0 = v$JLO_10310_out0;
assign v$_7486_out0 = { v$IR1$N_11003_out0,v$C4_11121_out0 };
assign v$_7487_out0 = { v$IR1$N_11004_out0,v$C4_11122_out0 };
assign v$INTERRUPT0_7520_out0 = v$EDGE0_3772_out0;
assign v$INTERRUPT0_7521_out0 = v$EDGE0_3773_out0;
assign v$STP_7534_out0 = v$STP_4222_out0;
assign v$STP_7535_out0 = v$STP_4223_out0;
assign v$G16_7742_out0 = ! v$IR1$W_11628_out0;
assign v$G16_7743_out0 = ! v$IR1$W_11629_out0;
assign v$JMI_8762_out0 = v$JMI_72_out0;
assign v$JMI_8763_out0 = v$JMI_73_out0;
assign v$G24_9384_out0 = v$G25_2250_out0 && v$G4_11042_out0;
assign v$G24_9385_out0 = v$G25_2251_out0 && v$G4_11043_out0;
assign v$EQ5_9756_out0 = v$IR1$OPCODE_1671_out0 == 4'h0;
assign v$EQ5_9757_out0 = v$IR1$OPCODE_1672_out0 == 4'h0;
assign v$G10_10226_out0 = ! v$STOP$1_5336_out0;
assign v$G10_10227_out0 = ! v$STOP$1_5337_out0;
assign v$EDGE1_10589_out0 = v$G19_11762_out0;
assign v$EDGE1_10590_out0 = v$G19_11763_out0;
assign v$IS$IR1$FMUL_10613_out0 = v$G22_10900_out0;
assign v$IS$IR1$FMUL_10614_out0 = v$G22_10901_out0;
assign v$JLS_11527_out0 = v$JLS_1096_out0;
assign v$JLS_11528_out0 = v$JLS_1097_out0;
assign v$G27_11608_out0 = v$G23_11817_out0 || v$G31_997_out0;
assign v$G27_11609_out0 = v$G23_11818_out0 || v$G31_998_out0;
assign v$EQ3_12697_out0 = v$IR1$OPCODE_1671_out0 == 4'h0;
assign v$EQ3_12698_out0 = v$IR1$OPCODE_1672_out0 == 4'h0;
assign v$G2_13111_out0 = ! v$IR1$L_3512_out0;
assign v$G2_13112_out0 = ! v$IR1$L_3513_out0;
assign v$G8_13406_out0 = ! v$IR1$U_10127_out0;
assign v$G8_13407_out0 = ! v$IR1$U_10128_out0;
assign v$_500_out0 = { v$_3459_out0,v$_8688_out0 };
assign v$_501_out0 = { v$_3460_out0,v$_8689_out0 };
assign v$DIN_903_out0 = v$_7486_out0;
assign v$DIN_904_out0 = v$_7487_out0;
assign v$MUX11_3121_out0 = v$IS$IR1$FMUL_10613_out0 ? v$IR1$FPU$OP_2545_out0 : v$IR2$FPU$OP_881_out0;
assign v$MUX11_3122_out0 = v$IS$IR1$FMUL_10614_out0 ? v$IR1$FPU$OP_2546_out0 : v$IR2$FPU$OP_882_out0;
assign v$G17_3706_out0 = v$JLO_5611_out0 && v$G18_9091_out0;
assign v$G17_3707_out0 = v$JLO_5612_out0 && v$G18_9092_out0;
assign v$G29_3728_out0 = v$G32_1001_out0 && v$R3_10621_out0;
assign v$G29_3729_out0 = v$G32_1002_out0 && v$R3_10622_out0;
assign v$G9_3818_out0 = ! v$INTERRUPT0_7520_out0;
assign v$G9_3819_out0 = ! v$INTERRUPT0_7521_out0;
assign v$G5_5122_out0 = v$G3_1573_out0 && v$IR15_7240_out0;
assign v$G5_5123_out0 = v$G3_1574_out0 && v$IR15_7241_out0;
assign v$G20_7982_out0 = v$EQ5_9756_out0 && v$IR1$L_3512_out0;
assign v$G20_7983_out0 = v$EQ5_9757_out0 && v$IR1$L_3513_out0;
assign v$SUBEN_8502_out0 = v$G8_13406_out0;
assign v$SUBEN_8503_out0 = v$G8_13407_out0;
assign v$STALL_8758_out0 = v$G27_11608_out0;
assign v$STALL_8759_out0 = v$G27_11609_out0;
assign v$G3_9569_out0 = v$EQ3_12697_out0 && v$G2_13111_out0;
assign v$G3_9570_out0 = v$EQ3_12698_out0 && v$G2_13112_out0;
assign v$G7_10034_out0 = v$INTERRUPT0_7520_out0 && v$G1_9855_out0;
assign v$G7_10035_out0 = v$INTERRUPT0_7521_out0 && v$G1_9856_out0;
assign v$G30_11118_out0 = v$FF4_13119_out0 && v$G28_1895_out0;
assign v$G30_11119_out0 = v$FF4_13120_out0 && v$G28_1896_out0;
assign v$STP_12552_out0 = v$STP_7534_out0;
assign v$STP_12553_out0 = v$STP_7535_out0;
assign v$G15_13187_out0 = v$IR1$P_2407_out0 || v$G16_7742_out0;
assign v$G15_13188_out0 = v$IR1$P_2408_out0 || v$G16_7743_out0;
assign v$OP_553_out0 = v$MUX11_3121_out0;
assign v$OP_554_out0 = v$MUX11_3122_out0;
assign v$G27_1425_out0 = v$G30_11118_out0 && v$F3_5730_out0;
assign v$G27_1426_out0 = v$G30_11119_out0 && v$F3_5731_out0;
assign v$G8_4049_out0 = v$G7_10034_out0 && v$R0_10497_out0;
assign v$G8_4050_out0 = v$G7_10035_out0 && v$R0_10498_out0;
assign v$G43_4800_out0 = v$STALL_8758_out0 && v$IR2$VALID_2898_out0;
assign v$G43_4801_out0 = v$STALL_8759_out0 && v$IR2$VALID_2899_out0;
assign v$STP_7120_out0 = v$STP_12552_out0;
assign v$STP_7121_out0 = v$STP_12553_out0;
assign v$MUX1_7566_out0 = v$SUBEN_8502_out0 ? v$C2_7980_out0 : v$C1_12939_out0;
assign v$MUX1_7567_out0 = v$SUBEN_8503_out0 ? v$C2_7981_out0 : v$C1_12940_out0;
assign v$G10_8887_out0 = v$FF1_4029_out0 && v$G9_3818_out0;
assign v$G10_8888_out0 = v$FF1_4030_out0 && v$G9_3819_out0;
assign v$QP_13189_out0 = v$_500_out0;
assign v$QP_13190_out0 = v$_501_out0;
assign v$G10_471_out0 = v$EQ11_9167_out0 && v$STP_7120_out0;
assign v$G10_472_out0 = v$EQ11_9168_out0 && v$STP_7121_out0;
assign v$G33_502_out0 = v$G29_3728_out0 || v$G27_1425_out0;
assign v$G33_503_out0 = v$G29_3729_out0 || v$G27_1426_out0;
assign v$G11_823_out0 = v$G10_8887_out0 && v$F0_11052_out0;
assign v$G11_824_out0 = v$G10_8888_out0 && v$F0_11053_out0;
assign v$G8_1170_out0 = v$EQ9_12558_out0 && v$STP_7120_out0;
assign v$G8_1171_out0 = v$EQ9_12559_out0 && v$STP_7121_out0;
assign v$G7_1889_out0 = v$EQ10_8978_out0 && v$STP_7120_out0;
assign v$G7_1890_out0 = v$EQ10_8979_out0 && v$STP_7121_out0;
assign v$G12_3238_out0 = v$G43_4800_out0 && v$INITIAL$FETCH$OCCURRED_759_out0;
assign v$G12_3239_out0 = v$G43_4801_out0 && v$INITIAL$FETCH$OCCURRED_760_out0;
assign v$XOR1_3455_out0 = v$MUX1_7566_out0 ^ v$DIN_903_out0;
assign v$XOR1_3456_out0 = v$MUX1_7567_out0 ^ v$DIN_904_out0;
assign v$G6_3710_out0 = v$EQ7_11947_out0 && v$STP_7120_out0;
assign v$G6_3711_out0 = v$EQ7_11948_out0 && v$STP_7121_out0;
assign v$G14_4440_out0 = v$EQ13_13201_out0 && v$STP_7120_out0;
assign v$G14_4441_out0 = v$EQ13_13202_out0 && v$STP_7121_out0;
assign v$EQ5_6738_out0 = v$QP_13189_out0 == 4'hb;
assign v$EQ5_6739_out0 = v$QP_13190_out0 == 4'hb;
assign v$FPU$OP_9460_out0 = v$OP_553_out0;
assign v$FPU$OP_9461_out0 = v$OP_554_out0;
assign v$G9_10434_out0 = v$EQ8_9715_out0 && v$STP_7120_out0;
assign v$G9_10435_out0 = v$EQ8_9716_out0 && v$STP_7121_out0;
assign v$G37_585_out0 = v$G12_3238_out0 && v$G48_3270_out0;
assign v$G37_586_out0 = v$G12_3239_out0 && v$G48_3271_out0;
assign v$EQ5_1729_out0 = v$FPU$OP_9460_out0 == 2'h3;
assign v$EQ5_1730_out0 = v$FPU$OP_9461_out0 == 2'h3;
assign v$EQ2_2910_out0 = v$FPU$OP_9460_out0 == 2'h0;
assign v$EQ2_2911_out0 = v$FPU$OP_9461_out0 == 2'h0;
assign v$INTDISABLE_3392_out0 = v$G7_1889_out0;
assign v$INTDISABLE_3393_out0 = v$G7_1890_out0;
assign v$NEXTINT_4763_out0 = v$G10_471_out0;
assign v$NEXTINT_4764_out0 = v$G10_472_out0;
assign v$INTCLEAR_5308_out0 = v$G8_1170_out0;
assign v$INTCLEAR_5309_out0 = v$G8_1171_out0;
assign v$EDGE3_7278_out0 = v$G33_502_out0;
assign v$EDGE3_7279_out0 = v$G33_503_out0;
assign v$FPU$OP_8416_out0 = v$FPU$OP_9460_out0;
assign v$FPU$OP_8417_out0 = v$FPU$OP_9461_out0;
assign v$LDMAINPC_9191_out0 = v$G14_4440_out0;
assign v$LDMAINPC_9192_out0 = v$G14_4441_out0;
assign v$EQ3_9316_out0 = v$FPU$OP_9460_out0 == 2'h2;
assign v$EQ3_9317_out0 = v$FPU$OP_9461_out0 == 2'h2;
assign v$G12_10062_out0 = v$G8_4049_out0 || v$G11_823_out0;
assign v$G12_10063_out0 = v$G8_4050_out0 || v$G11_824_out0;
assign v$EQ1_10605_out0 = v$FPU$OP_9460_out0 == 2'h1;
assign v$EQ1_10606_out0 = v$FPU$OP_9461_out0 == 2'h1;
assign v$EQ6_11337_out0 = v$FPU$OP_9460_out0 == 2'h3;
assign v$EQ6_11338_out0 = v$FPU$OP_9461_out0 == 2'h3;
assign v$EQ4_11767_out0 = v$FPU$OP_9460_out0 == 2'h3;
assign v$EQ4_11768_out0 = v$FPU$OP_9461_out0 == 2'h3;
assign v$G66_11892_out0 = !(v$G69_489_out0 && v$EQ5_6738_out0);
assign v$G66_11893_out0 = !(v$G69_490_out0 && v$EQ5_6739_out0);
assign v$NEXTINTERRUPT_13199_out0 = v$G10_471_out0;
assign v$NEXTINTERRUPT_13200_out0 = v$G10_472_out0;
assign v$INTCLR_194_out0 = v$INTCLEAR_5308_out0;
assign v$INTCLR_195_out0 = v$INTCLEAR_5309_out0;
assign v$G35_445_out0 = v$G37_585_out0 && v$G36_12163_out0;
assign v$G35_446_out0 = v$G37_586_out0 && v$G36_12164_out0;
assign v$G8_509_out0 = v$EQ4_11767_out0 && v$LOADA_3453_out0;
assign v$G8_510_out0 = v$EQ4_11768_out0 && v$LOADA_3454_out0;
assign v$INTDISABLE_1581_out0 = v$INTDISABLE_3392_out0;
assign v$INTDISABLE_1582_out0 = v$INTDISABLE_3393_out0;
assign v$G16_2547_out0 = ! v$EQ6_11337_out0;
assign v$G16_2548_out0 = ! v$EQ6_11338_out0;
assign v$EDGE0_2712_out0 = v$G12_10062_out0;
assign v$EDGE0_2713_out0 = v$G12_10063_out0;
assign v$G34_3310_out0 = v$NEXTINTERRUPT_13199_out0 || v$FF2_469_out0;
assign v$G34_3311_out0 = v$NEXTINTERRUPT_13200_out0 || v$FF2_470_out0;
assign v$ADD_5712_out0 = v$EQ2_2910_out0;
assign v$ADD_5713_out0 = v$EQ2_2911_out0;
assign v$FPU$LOAD$STORE_7238_out0 = v$EQ4_11767_out0;
assign v$FPU$LOAD$STORE_7239_out0 = v$EQ4_11768_out0;
assign v$G12_7750_out0 = v$G11_8976_out0 && v$EQ5_1729_out0;
assign v$G12_7751_out0 = v$G11_8977_out0 && v$EQ5_1730_out0;
assign v$G15_8990_out0 = v$G6_3710_out0 || v$NEXTINT_4763_out0;
assign v$G15_8991_out0 = v$G6_3711_out0 || v$NEXTINT_4764_out0;
assign v$SUB_9314_out0 = v$EQ1_10605_out0;
assign v$SUB_9315_out0 = v$EQ1_10606_out0;
assign v$LDMAIN_9330_out0 = v$LDMAINPC_9191_out0;
assign v$LDMAIN_9331_out0 = v$LDMAINPC_9192_out0;
assign v$G65_9509_out0 = v$G66_11892_out0 && v$CLK4_1439_out0;
assign v$G65_9510_out0 = v$G66_11893_out0 && v$CLK4_1440_out0;
assign v$EQ1_11375_out0 = v$FPU$OP_8416_out0 == 2'h1;
assign v$EQ1_11376_out0 = v$FPU$OP_8417_out0 == 2'h1;
assign v$G9_12027_out0 = v$EQ4_11767_out0 && v$G10_9966_out0;
assign v$G9_12028_out0 = v$EQ4_11768_out0 && v$G10_9967_out0;
assign v$MUL_12088_out0 = v$EQ3_9316_out0;
assign v$MUL_12089_out0 = v$EQ3_9317_out0;
assign v$CLRINTERRUPTS_276_out0 = v$INTCLR_194_out0;
assign v$CLRINTERRUPTS_277_out0 = v$INTCLR_195_out0;
assign v$INTENABLE_1705_out0 = v$G15_8990_out0;
assign v$INTENABLE_1706_out0 = v$G15_8991_out0;
assign v$G2_2437_out0 = v$ADD_5712_out0 || v$SUB_9314_out0;
assign v$G2_2438_out0 = v$ADD_5713_out0 || v$SUB_9315_out0;
assign v$G17_3764_out0 = v$G15_1205_out0 && v$G16_2547_out0;
assign v$G17_3765_out0 = v$G15_1206_out0 && v$G16_2548_out0;
assign v$G13_5410_out0 = v$G9_12027_out0 && v$IR2$IS$FPU_7643_out0;
assign v$G13_5411_out0 = v$G9_12028_out0 && v$IR2$IS$FPU_7644_out0;
assign v$G6_5440_out0 = v$ADD_5712_out0 || v$SUB_9314_out0;
assign v$G6_5441_out0 = v$ADD_5713_out0 || v$SUB_9315_out0;
assign v$G35_6881_out0 = v$INTDISABLE_1581_out0 || v$AUTODISABLE_12944_out0;
assign v$G35_6882_out0 = v$INTDISABLE_1582_out0 || v$AUTODISABLE_12945_out0;
assign v$STOPBITERROR_7542_out0 = v$G65_9509_out0;
assign v$STOPBITERROR_7543_out0 = v$G65_9510_out0;
assign v$G21_10066_out0 = v$G20_8064_out0 && v$FPU$LOAD$STORE_7238_out0;
assign v$G21_10067_out0 = v$G20_8065_out0 && v$FPU$LOAD$STORE_7239_out0;
assign v$G14_11038_out0 = v$G8_509_out0 && v$IR2$IS$FPU_7643_out0;
assign v$G14_11039_out0 = v$G8_510_out0 && v$IR2$IS$FPU_7644_out0;
assign v$STALL_12672_out0 = v$G35_445_out0;
assign v$STALL_12673_out0 = v$G35_446_out0;
assign v$NEXTINTERRUPT_13115_out0 = v$G34_3310_out0;
assign v$NEXTINTERRUPT_13116_out0 = v$G34_3311_out0;
assign v$STOPERROR_246_out0 = v$STOPBITERROR_7542_out0;
assign v$STOPERROR_247_out0 = v$STOPBITERROR_7543_out0;
assign v$CLR_3083_out0 = v$CLRINTERRUPTS_276_out0;
assign v$CLR_3084_out0 = v$CLRINTERRUPTS_277_out0;
assign v$G49_3615_out0 = ! v$STALL_12672_out0;
assign v$G49_3616_out0 = ! v$STALL_12673_out0;
assign v$G18_5076_out0 = v$G17_3764_out0 && v$IR2$VALID_11092_out0;
assign v$G18_5077_out0 = v$G17_3765_out0 && v$IR2$VALID_11093_out0;
assign v$G3_6377_out0 = v$MUL_12088_out0 || v$G6_5440_out0;
assign v$G3_6378_out0 = v$MUL_12089_out0 || v$G6_5441_out0;
assign v$NEXTINTERRUPT_8406_out0 = v$NEXTINTERRUPT_13115_out0;
assign v$NEXTINTERRUPT_8407_out0 = v$NEXTINTERRUPT_13116_out0;
assign v$DISABLEINTERRUPTS_10305_out0 = v$G35_6881_out0;
assign v$DISABLEINTERRUPTS_10306_out0 = v$G35_6882_out0;
assign v$STALL_10775_out0 = v$STALL_12672_out0;
assign v$STALL_10776_out0 = v$STALL_12673_out0;
assign v$INTENABLE_12210_out0 = v$INTENABLE_1705_out0;
assign v$INTENABLE_12211_out0 = v$INTENABLE_1706_out0;
assign v$G4_3292_out0 = v$ERR_8428_out0 || v$STOPERROR_246_out0;
assign v$G4_3293_out0 = v$ERR_8429_out0 || v$STOPERROR_247_out0;
assign v$G27_7528_out0 = v$STP$DECODED_11614_out0 || v$G49_3615_out0;
assign v$G27_7529_out0 = v$STP$DECODED_11615_out0 || v$G49_3616_out0;
assign v$STALL_8002_out0 = v$STALL_10775_out0;
assign v$STALL_8003_out0 = v$STALL_10776_out0;
assign v$ENABLEINTERRUPTS_8182_out0 = v$INTENABLE_12210_out0;
assign v$ENABLEINTERRUPTS_8183_out0 = v$INTENABLE_12211_out0;
assign v$G19_11088_out0 = v$G21_10066_out0 || v$G3_6377_out0;
assign v$G19_11089_out0 = v$G21_10067_out0 || v$G3_6378_out0;
assign v$NEXTINTERRUPT_11825_out0 = v$NEXTINTERRUPT_8406_out0;
assign v$NEXTINTERRUPT_11826_out0 = v$NEXTINTERRUPT_8407_out0;
assign v$R_13033_out0 = v$DISABLEINTERRUPTS_10305_out0;
assign v$R_13036_out0 = v$CLR_3083_out0;
assign v$R_13044_out0 = v$DISABLEINTERRUPTS_10306_out0;
assign v$R_13047_out0 = v$CLR_3084_out0;
assign v$G7_727_out0 = v$G19_11088_out0 && v$IR2$VALID_11092_out0;
assign v$G7_728_out0 = v$G19_11089_out0 && v$IR2$VALID_11093_out0;
assign v$G3_2802_out0 = v$I0P_3002_out0 && v$NEXTINTERRUPT_11825_out0;
assign v$G3_2803_out0 = v$I0P_3003_out0 && v$NEXTINTERRUPT_11826_out0;
assign v$G1_4832_out0 = v$I2P_5068_out0 && v$NEXTINTERRUPT_11825_out0;
assign v$G1_4833_out0 = v$I2P_5069_out0 && v$NEXTINTERRUPT_11826_out0;
assign v$G2_5802_out0 = v$I3P_7124_out0 && v$NEXTINTERRUPT_11825_out0;
assign v$G2_5803_out0 = v$I3P_7125_out0 && v$NEXTINTERRUPT_11826_out0;
assign v$G3_6660_out0 = v$INITIAL$FETCH$OCCURRED_759_out0 && v$G27_7528_out0;
assign v$G3_6661_out0 = v$INITIAL$FETCH$OCCURRED_760_out0 && v$G27_7529_out0;
assign v$PIPELINEHALT_10164_out0 = v$STALL_8002_out0;
assign v$PIPELINEHALT_10165_out0 = v$STALL_8003_out0;
assign v$G4_10750_out0 = v$I1P_1427_out0 && v$NEXTINTERRUPT_11825_out0;
assign v$G4_10751_out0 = v$I1P_1428_out0 && v$NEXTINTERRUPT_11826_out0;
assign v$G6_10834_out0 = ! v$R_13033_out0;
assign v$G6_10837_out0 = ! v$R_13036_out0;
assign v$G6_10845_out0 = ! v$R_13044_out0;
assign v$G6_10848_out0 = ! v$R_13047_out0;
assign v$S_11984_out0 = v$ENABLEINTERRUPTS_8182_out0;
assign v$S_11995_out0 = v$ENABLEINTERRUPTS_8183_out0;
assign v$SetError_12380_out0 = v$G4_3292_out0;
assign v$SetError_12381_out0 = v$G4_3293_out0;
assign v$G9_1435_out0 = v$CLR_3083_out0 || v$G4_10750_out0;
assign v$G9_1436_out0 = v$CLR_3084_out0 || v$G4_10751_out0;
assign v$G11_1773_out0 = v$CLR_3083_out0 || v$G2_5802_out0;
assign v$G11_1774_out0 = v$CLR_3084_out0 || v$G2_5803_out0;
assign v$G10_4679_out0 = v$CLR_3083_out0 || v$G1_4832_out0;
assign v$G10_4680_out0 = v$CLR_3084_out0 || v$G1_4833_out0;
assign v$WENFPU_9279_out0 = v$G7_727_out0;
assign v$WENFPU_9280_out0 = v$G7_728_out0;
assign v$G8_9653_out0 = v$FF2_8663_out0 || v$S_11984_out0;
assign v$G8_9659_out0 = v$FF2_8674_out0 || v$S_11995_out0;
assign v$G8_10770_out0 = v$CLR_3083_out0 || v$G3_2802_out0;
assign v$G8_10771_out0 = v$CLR_3084_out0 || v$G3_2803_out0;
assign v$G50_11471_out0 = v$G51_9413_out0 && v$G3_6660_out0;
assign v$G50_11472_out0 = v$G51_9414_out0 && v$G3_6661_out0;
assign v$S_11993_out0 = v$SetError_12380_out0;
assign v$S_12004_out0 = v$SetError_12381_out0;
assign v$WENFPU_2200_out0 = v$WENFPU_9279_out0;
assign v$WENFPU_2201_out0 = v$WENFPU_9280_out0;
assign v$G7_9512_out0 = v$G8_9653_out0 && v$G6_10834_out0;
assign v$G7_9518_out0 = v$G8_9659_out0 && v$G6_10845_out0;
assign v$IR1$VALID_12593_out0 = v$G50_11471_out0;
assign v$IR1$VALID_12594_out0 = v$G50_11472_out0;
assign v$R_13032_out0 = v$G8_10770_out0;
assign v$R_13034_out0 = v$G10_4679_out0;
assign v$R_13035_out0 = v$G11_1773_out0;
assign v$R_13037_out0 = v$G9_1435_out0;
assign v$R_13043_out0 = v$G8_10771_out0;
assign v$R_13045_out0 = v$G10_4680_out0;
assign v$R_13046_out0 = v$G11_1774_out0;
assign v$R_13048_out0 = v$G9_1436_out0;
assign v$IR1$VALID_6451_out0 = v$IR1$VALID_12593_out0;
assign v$IR1$VALID_6452_out0 = v$IR1$VALID_12594_out0;
assign v$Q_9529_out0 = v$G7_9512_out0;
assign v$Q_9540_out0 = v$G7_9518_out0;
assign v$G6_10833_out0 = ! v$R_13032_out0;
assign v$G6_10835_out0 = ! v$R_13034_out0;
assign v$G6_10836_out0 = ! v$R_13035_out0;
assign v$G6_10838_out0 = ! v$R_13037_out0;
assign v$G6_10844_out0 = ! v$R_13043_out0;
assign v$G6_10846_out0 = ! v$R_13045_out0;
assign v$G6_10847_out0 = ! v$R_13046_out0;
assign v$G6_10849_out0 = ! v$R_13048_out0;
assign v$IR1$VALID_3778_out0 = v$IR1$VALID_6451_out0;
assign v$IR1$VALID_3779_out0 = v$IR1$VALID_6452_out0;
assign v$ENABLEINTERRUPTS_12084_out0 = v$Q_9529_out0;
assign v$ENABLEINTERRUPTS_12085_out0 = v$Q_9540_out0;
assign v$G19_272_out0 = v$EDGE0_2712_out0 && v$ENABLEINTERRUPTS_12084_out0;
assign v$G19_273_out0 = v$EDGE0_2713_out0 && v$ENABLEINTERRUPTS_12085_out0;
assign v$G22_3274_out0 = v$EDGE3_7278_out0 && v$ENABLEINTERRUPTS_12084_out0;
assign v$G22_3275_out0 = v$EDGE3_7279_out0 && v$ENABLEINTERRUPTS_12085_out0;
assign v$IR1$VALID_9411_out0 = v$IR1$VALID_3778_out0;
assign v$IR1$VALID_9412_out0 = v$IR1$VALID_3779_out0;
assign v$G21_11040_out0 = v$EDGE2_12853_out0 && v$ENABLEINTERRUPTS_12084_out0;
assign v$G21_11041_out0 = v$EDGE2_12854_out0 && v$ENABLEINTERRUPTS_12085_out0;
assign v$G20_11140_out0 = v$EDGE1_10589_out0 && v$ENABLEINTERRUPTS_12084_out0;
assign v$G20_11141_out0 = v$EDGE1_10590_out0 && v$ENABLEINTERRUPTS_12085_out0;
assign v$G13_3006_out0 = v$G21_11040_out0 || v$G22_3274_out0;
assign v$G13_3007_out0 = v$G21_11041_out0 || v$G22_3275_out0;
assign v$G24_5412_out0 = v$LASTQ_7875_out0 && v$G21_11040_out0;
assign v$G24_5413_out0 = v$LASTQ_7886_out0 && v$G21_11041_out0;
assign v$G12_7686_out0 = v$G19_272_out0 || v$G20_11140_out0;
assign v$G12_7687_out0 = v$G19_273_out0 || v$G20_11141_out0;
assign v$G26_8296_out0 = v$LASTQ_7873_out0 && v$G19_272_out0;
assign v$G26_8297_out0 = v$LASTQ_7884_out0 && v$G19_273_out0;
assign v$G25_8634_out0 = v$LASTQ_7878_out0 && v$G20_11140_out0;
assign v$G25_8635_out0 = v$LASTQ_7889_out0 && v$G20_11141_out0;
assign v$S_11983_out0 = v$G19_272_out0;
assign v$S_11985_out0 = v$G21_11040_out0;
assign v$S_11986_out0 = v$G22_3274_out0;
assign v$S_11988_out0 = v$G20_11140_out0;
assign v$S_11994_out0 = v$G19_273_out0;
assign v$S_11996_out0 = v$G21_11041_out0;
assign v$S_11997_out0 = v$G22_3275_out0;
assign v$S_11999_out0 = v$G20_11141_out0;
assign v$IR1$VALID_13109_out0 = v$IR1$VALID_9411_out0;
assign v$IR1$VALID_13110_out0 = v$IR1$VALID_9412_out0;
assign v$G23_13291_out0 = v$LASTQ_7876_out0 && v$G22_3274_out0;
assign v$G23_13292_out0 = v$LASTQ_7887_out0 && v$G22_3275_out0;
assign v$G6_231_out0 = v$G5_11636_out0 && v$IR1$VALID_13109_out0;
assign v$G6_232_out0 = v$G5_11637_out0 && v$IR1$VALID_13110_out0;
assign v$IR1$VALID_2556_out0 = v$IR1$VALID_13109_out0;
assign v$IR1$VALID_2557_out0 = v$IR1$VALID_13110_out0;
assign v$G23_4753_out0 = v$EQ8_217_out0 && v$IR1$VALID_13109_out0;
assign v$G23_4754_out0 = v$EQ8_218_out0 && v$IR1$VALID_13110_out0;
assign v$G7_6658_out0 = v$IR1$VALID_13109_out0 && v$IS$IR1$FMUL_10613_out0;
assign v$G7_6659_out0 = v$IR1$VALID_13110_out0 && v$IS$IR1$FMUL_10614_out0;
assign v$G8_9652_out0 = v$FF2_8662_out0 || v$S_11983_out0;
assign v$G8_9654_out0 = v$FF2_8664_out0 || v$S_11985_out0;
assign v$G8_9655_out0 = v$FF2_8665_out0 || v$S_11986_out0;
assign v$G8_9657_out0 = v$FF2_8667_out0 || v$S_11988_out0;
assign v$G8_9658_out0 = v$FF2_8673_out0 || v$S_11994_out0;
assign v$G8_9660_out0 = v$FF2_8675_out0 || v$S_11996_out0;
assign v$G8_9661_out0 = v$FF2_8676_out0 || v$S_11997_out0;
assign v$G8_9663_out0 = v$FF2_8678_out0 || v$S_11999_out0;
assign v$G14_10607_out0 = v$G12_7686_out0 || v$G13_3006_out0;
assign v$G14_10608_out0 = v$G12_7687_out0 || v$G13_3007_out0;
assign v$G28_10676_out0 = v$G24_5412_out0 || v$G23_13291_out0;
assign v$G28_10677_out0 = v$G24_5413_out0 || v$G23_13292_out0;
assign v$G27_13157_out0 = v$G26_8296_out0 || v$G25_8634_out0;
assign v$G27_13158_out0 = v$G26_8297_out0 || v$G25_8635_out0;
assign v$IR1$VALID_58_out0 = v$IR1$VALID_2556_out0;
assign v$IR1$VALID_59_out0 = v$IR1$VALID_2557_out0;
assign v$INCOMINGINTERRUPT_1054_out0 = v$G14_10607_out0;
assign v$INCOMINGINTERRUPT_1055_out0 = v$G14_10608_out0;
assign v$MUX9_5181_out0 = v$G6_231_out0 ? v$IR1$D_2900_out0 : v$IR2$D_9879_out0;
assign v$MUX9_5182_out0 = v$G6_232_out0 ? v$IR1$D_2901_out0 : v$IR2$D_9880_out0;
assign v$G8_8123_out0 = v$G10_6837_out0 || v$G6_231_out0;
assign v$G8_8124_out0 = v$G10_6838_out0 || v$G6_232_out0;
assign v$EXEC1$FPU_9221_out0 = v$G7_6658_out0;
assign v$EXEC1$FPU_9222_out0 = v$G7_6659_out0;
assign v$G7_9511_out0 = v$G8_9652_out0 && v$G6_10833_out0;
assign v$G7_9513_out0 = v$G8_9654_out0 && v$G6_10835_out0;
assign v$G7_9514_out0 = v$G8_9655_out0 && v$G6_10836_out0;
assign v$G7_9516_out0 = v$G8_9657_out0 && v$G6_10838_out0;
assign v$G7_9517_out0 = v$G8_9658_out0 && v$G6_10844_out0;
assign v$G7_9519_out0 = v$G8_9660_out0 && v$G6_10846_out0;
assign v$G7_9520_out0 = v$G8_9661_out0 && v$G6_10847_out0;
assign v$G7_9522_out0 = v$G8_9663_out0 && v$G6_10849_out0;
assign v$G29_11007_out0 = v$G27_13157_out0 || v$G28_10676_out0;
assign v$G29_11008_out0 = v$G27_13158_out0 || v$G28_10677_out0;
assign v$INTERRUPTOVERFLOW_1160_out0 = v$G29_11007_out0;
assign v$INTERRUPTOVERFLOW_1161_out0 = v$G29_11008_out0;
assign v$G19_1593_out0 = v$G20_7982_out0 && v$IR1$VALID_58_out0;
assign v$G19_1594_out0 = v$G20_7983_out0 && v$IR1$VALID_59_out0;
assign v$AD1_4656_out0 = v$MUX9_5181_out0;
assign v$AD1_4657_out0 = v$MUX9_5182_out0;
assign v$G13_6807_out0 = v$G8_8123_out0 || v$G23_4753_out0;
assign v$G13_6808_out0 = v$G8_8124_out0 || v$G23_4754_out0;
assign v$EXEC1_6827_out0 = v$EXEC1$FPU_9221_out0;
assign v$EXEC1_6828_out0 = v$EXEC1$FPU_9222_out0;
assign v$G17_7915_out0 = v$INCOMINGINTERRUPT_1054_out0 && v$G18_1749_out0;
assign v$G17_7916_out0 = v$INCOMINGINTERRUPT_1055_out0 && v$G18_1750_out0;
assign v$Q_9528_out0 = v$G7_9511_out0;
assign v$Q_9530_out0 = v$G7_9513_out0;
assign v$Q_9531_out0 = v$G7_9514_out0;
assign v$Q_9533_out0 = v$G7_9516_out0;
assign v$Q_9539_out0 = v$G7_9517_out0;
assign v$Q_9541_out0 = v$G7_9519_out0;
assign v$Q_9542_out0 = v$G7_9520_out0;
assign v$Q_9544_out0 = v$G7_9522_out0;
assign v$G5_10018_out0 = v$IR1$VALID_58_out0 && v$IR1$W_11628_out0;
assign v$G5_10019_out0 = v$IR1$VALID_59_out0 && v$IR1$W_11629_out0;
assign v$G4_10821_out0 = v$G3_9569_out0 && v$IR1$VALID_58_out0;
assign v$G4_10822_out0 = v$G3_9570_out0 && v$IR1$VALID_59_out0;
assign v$MUX10_2334_out0 = v$G13_6807_out0 ? v$IR1$M_8836_out0 : v$IR2$M_8626_out0;
assign v$MUX10_2335_out0 = v$G13_6808_out0 ? v$IR1$M_8837_out0 : v$IR2$M_8627_out0;
assign v$I3_3228_out0 = v$Q_9531_out0;
assign v$I3_3229_out0 = v$Q_9542_out0;
assign v$I1_3282_out0 = v$Q_9533_out0;
assign v$I1_3283_out0 = v$Q_9544_out0;
assign v$NEWINTERRUPT_3679_out0 = v$G17_7915_out0;
assign v$NEWINTERRUPT_3680_out0 = v$G17_7916_out0;
assign v$G16_4405_out0 = v$NEXTINTERRUPT_11825_out0 || v$G17_7915_out0;
assign v$G16_4406_out0 = v$NEXTINTERRUPT_11826_out0 || v$G17_7916_out0;
assign v$G6_5056_out0 = v$Q_9530_out0 || v$Q_9531_out0;
assign v$G6_5057_out0 = v$Q_9541_out0 || v$Q_9542_out0;
assign v$G7_7596_out0 = v$G5_10018_out0 || v$G6_7724_out0;
assign v$G7_7597_out0 = v$G5_10019_out0 || v$G6_7725_out0;
assign v$READ$REQUEST_9841_out0 = v$G19_1593_out0;
assign v$READ$REQUEST_9842_out0 = v$G19_1594_out0;
assign v$I2_9881_out0 = v$Q_9530_out0;
assign v$I2_9882_out0 = v$Q_9541_out0;
assign v$G11_9962_out0 = v$G4_10821_out0 && v$G10_10226_out0;
assign v$G11_9963_out0 = v$G4_10822_out0 && v$G10_10227_out0;
assign v$G5_11287_out0 = v$Q_9528_out0 || v$Q_9533_out0;
assign v$G5_11288_out0 = v$Q_9539_out0 || v$Q_9544_out0;
assign v$S_11987_out0 = v$INTERRUPTOVERFLOW_1160_out0;
assign v$S_11998_out0 = v$INTERRUPTOVERFLOW_1161_out0;
assign v$I0_13167_out0 = v$Q_9528_out0;
assign v$I0_13168_out0 = v$Q_9539_out0;
assign v$AD1_13302_out0 = v$AD1_4656_out0;
assign v$AD1_13303_out0 = v$AD1_4657_out0;
assign v$EXEC1_13347_out0 = v$EXEC1_6827_out0;
assign v$EXEC1_13348_out0 = v$EXEC1_6828_out0;
assign v$CAPTURE_207_out0 = v$G16_4405_out0;
assign v$CAPTURE_208_out0 = v$G16_4406_out0;
assign v$G7_1007_out0 = v$G5_11287_out0 || v$G6_5056_out0;
assign v$G7_1008_out0 = v$G5_11288_out0 || v$G6_5057_out0;
assign v$AD1_1011_out0 = v$AD1_13302_out0;
assign v$AD1_1012_out0 = v$AD1_13303_out0;
assign v$NEWINTERRUPT_4784_out0 = v$NEWINTERRUPT_3679_out0;
assign v$NEWINTERRUPT_4785_out0 = v$NEWINTERRUPT_3680_out0;
assign v$G4_5283_out0 = ! v$I1_3282_out0;
assign v$G4_5284_out0 = ! v$I1_3283_out0;
assign v$RAMWEN_5302_out0 = v$G11_9962_out0;
assign v$RAMWEN_5303_out0 = v$G11_9963_out0;
assign v$G2_5310_out0 = ! v$I3_3228_out0;
assign v$G2_5311_out0 = ! v$I3_3229_out0;
assign v$G3_6067_out0 = ! v$I2_9881_out0;
assign v$G3_6068_out0 = ! v$I2_9882_out0;
assign v$AD2_6334_out0 = v$MUX10_2334_out0;
assign v$AD2_6335_out0 = v$MUX10_2335_out0;
assign v$WENLDST_8125_out0 = v$G7_7596_out0;
assign v$WENLDST_8126_out0 = v$G7_7597_out0;
assign v$I3P_9176_out0 = v$I3_3228_out0;
assign v$I3P_9177_out0 = v$I3_3229_out0;
assign v$G8_9656_out0 = v$FF2_8666_out0 || v$S_11987_out0;
assign v$G8_9662_out0 = v$FF2_8677_out0 || v$S_11998_out0;
assign v$READ$REQUEST_11632_out0 = v$READ$REQUEST_9841_out0;
assign v$READ$REQUEST_11633_out0 = v$READ$REQUEST_9842_out0;
assign v$EXEC1_12950_out0 = v$EXEC1_13347_out0;
assign v$EXEC1_12951_out0 = v$EXEC1_13348_out0;
assign v$EXEC1_2564_out0 = v$EXEC1_12950_out0;
assign v$EXEC1_2565_out0 = v$EXEC1_12951_out0;
assign v$NEWINTERRUPT_3080_out0 = v$NEWINTERRUPT_4784_out0;
assign v$NEWINTERRUPT_3081_out0 = v$NEWINTERRUPT_4785_out0;
assign v$MUX1_3405_out0 = v$G16_4405_out0 ? v$G7_1007_out0 : v$FF1_8718_out0;
assign v$MUX1_3406_out0 = v$G16_4406_out0 ? v$G7_1008_out0 : v$FF1_8719_out0;
assign v$READ$REQUEST_5332_out0 = v$READ$REQUEST_11632_out0;
assign v$READ$REQUEST_5333_out0 = v$READ$REQUEST_11633_out0;
assign v$G7_7231_out0 = v$I0_13167_out0 && v$G4_5283_out0;
assign v$G7_7232_out0 = v$I0_13168_out0 && v$G4_5284_out0;
assign v$_7866_out0 = v$AD1_1011_out0[0:0];
assign v$_7866_out1 = v$AD1_1011_out0[1:1];
assign v$_7867_out0 = v$AD1_1012_out0[0:0];
assign v$_7867_out1 = v$AD1_1012_out0[1:1];
assign v$G1_9116_out0 = v$I2_9881_out0 && v$G2_5310_out0;
assign v$G1_9117_out0 = v$I2_9882_out0 && v$G2_5311_out0;
assign v$G7_9515_out0 = v$G8_9656_out0 && v$G6_10837_out0;
assign v$G7_9521_out0 = v$G8_9662_out0 && v$G6_10848_out0;
assign v$AD2_10930_out0 = v$AD2_6334_out0;
assign v$AD2_10931_out0 = v$AD2_6335_out0;
assign v$RAMWEN_10932_out0 = v$RAMWEN_5302_out0;
assign v$RAMWEN_10933_out0 = v$RAMWEN_5303_out0;
assign v$G8_12674_out0 = v$G3_6067_out0 && v$G2_5310_out0;
assign v$G8_12675_out0 = v$G3_6068_out0 && v$G2_5311_out0;
assign v$WENLDST_13265_out0 = v$WENLDST_8125_out0;
assign v$WENLDST_13266_out0 = v$WENLDST_8126_out0;
assign v$WENRAM_3362_out0 = v$RAMWEN_10932_out0;
assign v$WENRAM_3363_out0 = v$RAMWEN_10933_out0;
assign v$MUX1_3839_out0 = v$_7866_out0 ? v$REG1_3286_out0 : v$REG0_11406_out0;
assign v$MUX1_3840_out0 = v$_7867_out0 ? v$REG1_3287_out0 : v$REG0_11407_out0;
assign v$AD2_4413_out0 = v$AD2_10930_out0;
assign v$AD2_4414_out0 = v$AD2_10931_out0;
assign v$I2P_4445_out0 = v$G1_9116_out0;
assign v$I2P_4446_out0 = v$G1_9117_out0;
assign v$WENLDST_4677_out0 = v$WENLDST_13265_out0;
assign v$WENLDST_4678_out0 = v$WENLDST_13266_out0;
assign v$G12_6662_out0 = !(v$NEWINTERRUPT_3080_out0 || v$FF1_601_out0);
assign v$G12_6663_out0 = !(v$NEWINTERRUPT_3081_out0 || v$FF1_602_out0);
assign v$MUX2_7000_out0 = v$_7866_out0 ? v$REG3_7255_out0 : v$REG2_12278_out0;
assign v$MUX2_7001_out0 = v$_7867_out0 ? v$REG3_7256_out0 : v$REG2_12279_out0;
assign v$ISINTERRUPTED_7745_out0 = v$MUX1_3405_out0;
assign v$ISINTERRUPTED_7746_out0 = v$MUX1_3406_out0;
assign v$G6_7901_out0 = v$G7_7231_out0 && v$G8_12674_out0;
assign v$G6_7902_out0 = v$G7_7232_out0 && v$G8_12675_out0;
assign v$Q_9532_out0 = v$G7_9515_out0;
assign v$Q_9543_out0 = v$G7_9521_out0;
assign v$G9_10813_out0 = v$I1_3282_out0 && v$G8_12674_out0;
assign v$G9_10814_out0 = v$I1_3283_out0 && v$G8_12675_out0;
assign v$READ$REQUEST1_11877_out0 = v$READ$REQUEST_5333_out0;
assign v$READ$REQUEST0_13146_out0 = v$READ$REQUEST_5332_out0;
assign v$EXEC1_13169_out0 = v$EXEC1_2564_out0;
assign v$EXEC1_13170_out0 = v$EXEC1_2565_out0;
assign v$ININTERRUPT_433_out0 = v$ISINTERRUPTED_7745_out0;
assign v$ININTERRUPT_434_out0 = v$ISINTERRUPTED_7746_out0;
assign v$MUX3_787_out0 = v$_7866_out1 ? v$MUX2_7000_out0 : v$MUX1_3839_out0;
assign v$MUX3_788_out0 = v$_7867_out1 ? v$MUX2_7001_out0 : v$MUX1_3840_out0;
assign v$G11_1211_out0 = v$G9_10434_out0 && v$G12_6662_out0;
assign v$G11_1212_out0 = v$G9_10435_out0 && v$G12_6663_out0;
assign v$I0P_1365_out0 = v$G6_7901_out0;
assign v$I0P_1366_out0 = v$G6_7902_out0;
assign v$G11_1739_out0 = v$I2P_4445_out0 || v$I3P_9176_out0;
assign v$G11_1740_out0 = v$I2P_4446_out0 || v$I3P_9177_out0;
assign v$G2_2792_out0 = v$G24_9384_out0 && v$WENLDST_4677_out0;
assign v$G2_2793_out0 = v$G24_9385_out0 && v$WENLDST_4678_out0;
assign v$MUX8_3004_out0 = v$IR2$15_5012_out0 ? v$WENALU_2782_out0 : v$WENLDST_4677_out0;
assign v$MUX8_3005_out0 = v$IR2$15_5013_out0 ? v$WENALU_2783_out0 : v$WENLDST_4678_out0;
assign v$XOR1_3401_out0 = v$AD3_8756_out0 ^ v$AD2_4413_out0;
assign v$XOR1_3402_out0 = v$AD3_8757_out0 ^ v$AD2_4414_out0;
assign v$READ$REQUEST1_4462_out0 = v$READ$REQUEST1_11877_out0;
assign v$_4849_out0 = v$AD2_4413_out0[0:0];
assign v$_4849_out1 = v$AD2_4413_out0[1:1];
assign v$_4850_out0 = v$AD2_4414_out0[0:0];
assign v$_4850_out1 = v$AD2_4414_out0[1:1];
assign v$EXEC1_5456_out0 = v$EXEC1_13169_out0;
assign v$EXEC1_5457_out0 = v$EXEC1_13169_out0;
assign v$EXEC1_5458_out0 = v$EXEC1_13169_out0;
assign v$EXEC1_5459_out0 = v$EXEC1_13169_out0;
assign v$EXEC1_5460_out0 = v$EXEC1_13169_out0;
assign v$EXEC1_5461_out0 = v$EXEC1_13169_out0;
assign v$EXEC1_5462_out0 = v$EXEC1_13169_out0;
assign v$EXEC1_5463_out0 = v$EXEC1_13169_out0;
assign v$EXEC1_5464_out0 = v$EXEC1_13169_out0;
assign v$EXEC1_5465_out0 = v$EXEC1_13169_out0;
assign v$EXEC1_5466_out0 = v$EXEC1_13169_out0;
assign v$EXEC1_5467_out0 = v$EXEC1_13170_out0;
assign v$EXEC1_5468_out0 = v$EXEC1_13170_out0;
assign v$EXEC1_5469_out0 = v$EXEC1_13170_out0;
assign v$EXEC1_5470_out0 = v$EXEC1_13170_out0;
assign v$EXEC1_5471_out0 = v$EXEC1_13170_out0;
assign v$EXEC1_5472_out0 = v$EXEC1_13170_out0;
assign v$EXEC1_5473_out0 = v$EXEC1_13170_out0;
assign v$EXEC1_5474_out0 = v$EXEC1_13170_out0;
assign v$EXEC1_5475_out0 = v$EXEC1_13170_out0;
assign v$EXEC1_5476_out0 = v$EXEC1_13170_out0;
assign v$EXEC1_5477_out0 = v$EXEC1_13170_out0;
assign v$READ$REQUEST0_7434_out0 = v$READ$REQUEST0_13146_out0;
assign v$I1P_10166_out0 = v$G9_10813_out0;
assign v$I1P_10167_out0 = v$G9_10814_out0;
assign v$INTERRUPTOVERFLOW_10426_out0 = v$Q_9532_out0;
assign v$INTERRUPTOVERFLOW_10427_out0 = v$Q_9543_out0;
assign v$WENRAM_12116_out0 = v$WENRAM_3362_out0;
assign v$WENRAM_12117_out0 = v$WENRAM_3363_out0;
assign v$G3_0_out0 = v$G2_2792_out0 && v$IR1$VALID_13109_out0;
assign v$G3_1_out0 = v$G2_2793_out0 && v$IR1$VALID_13110_out0;
assign v$MUX4_849_out0 = v$_4849_out0 ? v$R1_9296_out0 : v$R0_1977_out0;
assign v$MUX4_850_out0 = v$_4850_out0 ? v$R1_9297_out0 : v$R0_1978_out0;
assign v$WENRAM_1277_out0 = v$WENRAM_12116_out0;
assign v$WENRAM_1278_out0 = v$WENRAM_12117_out0;
assign v$DOUT1_1887_out0 = v$MUX3_787_out0;
assign v$DOUT1_1888_out0 = v$MUX3_788_out0;
assign v$EQ1_1925_out0 = v$XOR1_3401_out0 == 2'h0;
assign v$EQ1_1926_out0 = v$XOR1_3402_out0 == 2'h0;
assign v$G10_2511_out0 = v$I1P_10166_out0 || v$I3P_9176_out0;
assign v$G10_2512_out0 = v$I1P_10167_out0 || v$I3P_9177_out0;
assign v$G14_3504_out0 = ! v$ININTERRUPT_433_out0;
assign v$G14_3505_out0 = ! v$ININTERRUPT_434_out0;
assign v$G52_5403_out0 = v$READ$REQUEST0_7434_out0 || v$FF2_9024_out0;
assign v$G44_5734_out0 = v$READ$REQUEST1_4462_out0 || v$FF1_3695_out0;
assign v$ARR1_6305_out0 = v$READ$REQUEST1_4462_out0;
assign v$ENCODED1_6496_out0 = v$G11_1739_out0;
assign v$ENCODED1_6497_out0 = v$G11_1740_out0;
assign v$G31_7100_out0 = v$NEXTINTERRUPT_13115_out0 && v$ININTERRUPT_433_out0;
assign v$G31_7101_out0 = v$NEXTINTERRUPT_13116_out0 && v$ININTERRUPT_434_out0;
assign v$ARR0_7237_out0 = v$READ$REQUEST0_7434_out0;
assign v$MUX5_7647_out0 = v$EQ1_13237_out0 ? v$WENFPU_2200_out0 : v$MUX8_3004_out0;
assign v$MUX5_7648_out0 = v$EQ1_13238_out0 ? v$WENFPU_2201_out0 : v$MUX8_3005_out0;
assign v$WEN_7946_out0 = v$WENRAM_12116_out0;
assign v$WEN_7947_out0 = v$WENRAM_12117_out0;
assign v$MUX5_9474_out0 = v$_4849_out0 ? v$R3_7072_out0 : v$R2_5454_out0;
assign v$MUX5_9475_out0 = v$_4850_out0 ? v$R3_7073_out0 : v$R2_5455_out0;
assign v$WEN_9615_out0 = v$WENRAM_12116_out0;
assign v$WEN_9616_out0 = v$WENRAM_12117_out0;
assign v$INTOVERFLOW_11219_out0 = v$INTERRUPTOVERFLOW_10426_out0;
assign v$INTOVERFLOW_11220_out0 = v$INTERRUPTOVERFLOW_10427_out0;
assign v$STPHALT_12859_out0 = v$G11_1211_out0;
assign v$STPHALT_12860_out0 = v$G11_1212_out0;
assign v$WENRAM1_899_out0 = v$WENRAM_1278_out0;
assign v$RR1_1093_out0 = v$G44_5734_out0;
assign v$RD_1154_out0 = v$DOUT1_1887_out0;
assign v$RD_1155_out0 = v$DOUT1_1888_out0;
assign v$WEN_2398_out0 = v$WEN_9615_out0;
assign v$WEN_2399_out0 = v$WEN_9616_out0;
assign v$WEN_2509_out0 = v$WEN_7946_out0;
assign v$WEN_2510_out0 = v$WEN_7947_out0;
assign v$STPHALT_2988_out0 = v$STPHALT_12859_out0;
assign v$STPHALT_2989_out0 = v$STPHALT_12860_out0;
assign v$MUX6_3439_out0 = v$_4849_out1 ? v$MUX5_9474_out0 : v$MUX4_849_out0;
assign v$MUX6_3440_out0 = v$_4850_out1 ? v$MUX5_9475_out0 : v$MUX4_850_out0;
assign v$G29_5378_out0 = v$NEWINTERRUPT_4784_out0 || v$G31_7100_out0;
assign v$G29_5379_out0 = v$NEWINTERRUPT_4785_out0 || v$G31_7101_out0;
assign v$RR0_5596_out0 = v$G52_5403_out0;
assign v$WENRAM0_6651_out0 = v$WENRAM_1277_out0;
assign v$G33_7075_out0 = v$LDMAIN_9330_out0 || v$G14_3504_out0;
assign v$G33_7076_out0 = v$LDMAIN_9331_out0 || v$G14_3505_out0;
assign v$MUX7_7229_out0 = v$IR2$VALID$AND$NOT$FLOAD_4883_out0 ? v$MUX5_7647_out0 : v$G3_0_out0;
assign v$MUX7_7230_out0 = v$IR2$VALID$AND$NOT$FLOAD_4884_out0 ? v$MUX5_7648_out0 : v$G3_1_out0;
assign v$ENCODED0_9415_out0 = v$G10_2511_out0;
assign v$ENCODED0_9416_out0 = v$G10_2512_out0;
assign v$AD3$EQUALS$AD2_9945_out0 = v$EQ1_1925_out0;
assign v$AD3$EQUALS$AD2_9946_out0 = v$EQ1_1926_out0;
assign v$OP1_10521_out0 = v$DOUT1_1887_out0;
assign v$OP1_10522_out0 = v$DOUT1_1888_out0;
assign v$WEN3_1983_out0 = v$MUX7_7229_out0;
assign v$WEN3_1984_out0 = v$MUX7_7230_out0;
assign v$DOUT2_2214_out0 = v$MUX6_3439_out0;
assign v$DOUT2_2215_out0 = v$MUX6_3440_out0;
assign v$OP1_3661_out0 = v$OP1_10521_out0;
assign v$OP1_3662_out0 = v$OP1_10522_out0;
assign v$A_5932_out0 = v$RD_1154_out0;
assign v$A_5933_out0 = v$RD_1155_out0;
assign v$RDOUT_6895_out0 = v$RD_1154_out0;
assign v$RDOUT_6896_out0 = v$RD_1155_out0;
assign v$RAMWEN1_7089_out0 = v$WENRAM1_899_out0;
assign v$WEN_8101_out0 = v$WEN_2509_out0;
assign v$WEN_8102_out0 = v$WEN_2510_out0;
assign v$_9984_out0 = { v$ENCODED0_9415_out0,v$ENCODED1_6496_out0 };
assign v$_9985_out0 = { v$ENCODED0_9416_out0,v$ENCODED1_6497_out0 };
assign v$RAMWEN0_11645_out0 = v$WENRAM0_6651_out0;
assign v$INTERRUPTNUMBER_36_out0 = v$_9984_out0;
assign v$INTERRUPTNUMBER_37_out0 = v$_9985_out0;
assign v$AWR0_972_out0 = v$RAMWEN0_11645_out0;
assign v$DATA$IN_4809_out0 = v$RDOUT_6895_out0;
assign v$DATA$IN_4810_out0 = v$RDOUT_6896_out0;
assign v$A_7280_out0 = v$A_5932_out0;
assign v$A_7281_out0 = v$A_5933_out0;
assign v$G55_9243_out0 = v$RAMWEN0_11645_out0 || v$FF3_2072_out0;
assign v$D1_9486_out0 = (v$AD3_8756_out0 == 2'b00) ? v$WEN3_1983_out0 : 1'h0;
assign v$D1_9486_out1 = (v$AD3_8756_out0 == 2'b01) ? v$WEN3_1983_out0 : 1'h0;
assign v$D1_9486_out2 = (v$AD3_8756_out0 == 2'b10) ? v$WEN3_1983_out0 : 1'h0;
assign v$D1_9486_out3 = (v$AD3_8756_out0 == 2'b11) ? v$WEN3_1983_out0 : 1'h0;
assign v$D1_9487_out0 = (v$AD3_8757_out0 == 2'b00) ? v$WEN3_1984_out0 : 1'h0;
assign v$D1_9487_out1 = (v$AD3_8757_out0 == 2'b01) ? v$WEN3_1984_out0 : 1'h0;
assign v$D1_9487_out2 = (v$AD3_8757_out0 == 2'b10) ? v$WEN3_1984_out0 : 1'h0;
assign v$D1_9487_out3 = (v$AD3_8757_out0 == 2'b11) ? v$WEN3_1984_out0 : 1'h0;
assign v$AWR1_11104_out0 = v$RAMWEN1_7089_out0;
assign v$RM_11349_out0 = v$DOUT2_2214_out0;
assign v$RM_11350_out0 = v$DOUT2_2215_out0;
assign v$A_11516_out0 = v$OP1_3661_out0;
assign v$A_11517_out0 = v$OP1_3662_out0;
assign v$G56_12500_out0 = v$RAMWEN1_7089_out0 || v$FF4_9118_out0;
assign v$WEN_13084_out0 = v$WEN_8101_out0;
assign v$WEN_13085_out0 = v$WEN_8102_out0;
assign v$RM_13239_out0 = v$DOUT2_2214_out0;
assign v$RM_13240_out0 = v$DOUT2_2215_out0;
assign v$WR1_255_out0 = v$G56_12500_out0;
assign v$G6_382_out0 = ! v$WEN_13084_out0;
assign v$G6_383_out0 = ! v$WEN_13085_out0;
assign v$G84_504_out0 = v$AWR1_11104_out0 || v$ARR1_6305_out0;
assign v$NINTERRUPT_798_out0 = v$INTERRUPTNUMBER_36_out0;
assign v$NINTERRUPT_799_out0 = v$INTERRUPTNUMBER_37_out0;
assign v$DATA$IN_811_out0 = v$DATA$IN_4809_out0;
assign v$DATA$IN_812_out0 = v$DATA$IN_4810_out0;
assign v$MUX1_985_out0 = v$C_4069_out0 ? v$_8000_out0 : v$RM_11349_out0;
assign v$MUX1_986_out0 = v$C_4070_out0 ? v$_8001_out0 : v$RM_11350_out0;
assign v$A_1456_out0 = v$A_11516_out0;
assign v$A_1457_out0 = v$A_11517_out0;
assign v$MUX13_1458_out0 = v$B$IS$RD_9476_out0 ? v$RD_1154_out0 : v$RM_13239_out0;
assign v$MUX13_1459_out0 = v$B$IS$RD_9477_out0 ? v$RD_1155_out0 : v$RM_13240_out0;
assign v$A_2886_out0 = v$A_7280_out0;
assign v$A_2887_out0 = v$A_7281_out0;
assign v$RAMDIN_4792_out0 = v$DATA$IN_4809_out0;
assign v$RAMDIN_4793_out0 = v$DATA$IN_4810_out0;
assign v$G88_4994_out0 = v$ARR0_7237_out0 || v$AWR0_972_out0;
assign v$RM_6813_out0 = v$RM_13239_out0;
assign v$RM_6814_out0 = v$RM_13240_out0;
assign v$G8_8973_out0 = ! v$WEN_13084_out0;
assign v$G8_8974_out0 = ! v$WEN_13085_out0;
assign v$DATA_9478_out0 = v$DATA$IN_4809_out0;
assign v$DATA_9479_out0 = v$DATA$IN_4810_out0;
assign v$WR0_9664_out0 = v$G55_9243_out0;
assign v$A_13003_out0 = v$A_7280_out0;
assign v$A_13004_out0 = v$A_7281_out0;
assign v$IN_180_out0 = v$MUX1_985_out0;
assign v$IN_181_out0 = v$MUX1_986_out0;
assign v$_392_out0 = v$A_1456_out0[7:4];
assign v$_393_out0 = v$A_1457_out0[7:4];
assign v$WR0_546_out0 = v$WR0_9664_out0;
assign v$DIN_977_out0 = v$RAMDIN_4792_out0;
assign v$DIN_978_out0 = v$RAMDIN_4793_out0;
assign v$A_1951_out0 = v$A_13003_out0;
assign v$A_1952_out0 = v$A_13004_out0;
assign v$_2507_out0 = v$A_1456_out0[15:12];
assign v$_2508_out0 = v$A_1457_out0[15:12];
assign v$_2854_out0 = v$A_1456_out0[3:0];
assign v$_2855_out0 = v$A_1457_out0[3:0];
assign v$DATA_3010_out0 = v$DATA_9478_out0;
assign v$DATA_3011_out0 = v$DATA_9479_out0;
assign v$_5930_out0 = v$A_1456_out0[11:8];
assign v$_5931_out0 = v$A_1457_out0[11:8];
assign v$SEL2_6423_out0 = v$NINTERRUPT_798_out0[0:0];
assign v$SEL2_6424_out0 = v$NINTERRUPT_799_out0[0:0];
assign v$DATA$IN0_6953_out0 = v$DATA$IN_811_out0;
assign v$G79_8390_out0 = v$RR0_5596_out0 || v$WR0_9664_out0;
assign v$B_9458_out0 = v$MUX13_1458_out0;
assign v$B_9459_out0 = v$MUX13_1459_out0;
assign v$WR1_9723_out0 = v$WR1_255_out0;
assign v$DATA$IN1_10600_out0 = v$DATA$IN_812_out0;
assign v$A_11271_out0 = v$A_2886_out0;
assign v$A_11272_out0 = v$A_2887_out0;
assign v$G36_11766_out0 = v$RR1_1093_out0 || v$WR1_255_out0;
assign v$SEL3_12208_out0 = v$NINTERRUPT_798_out0[1:1];
assign v$SEL3_12209_out0 = v$NINTERRUPT_799_out0[1:1];
assign v$RM_12933_out0 = v$RM_6813_out0;
assign v$RM_12934_out0 = v$RM_6814_out0;
assign v$SEL5_260_out0 = v$A_1951_out0[15:15];
assign v$SEL5_261_out0 = v$A_1952_out0[15:15];
assign v$MUX7_435_out0 = v$SEL2_6423_out0 ? v$INT3_233_out0 : v$INT2_221_out0;
assign v$MUX7_436_out0 = v$SEL2_6424_out0 ? v$INT3_234_out0 : v$INT2_222_out0;
assign v$_1024_out0 = { v$A$SAVED_6682_out0,v$A_11271_out0 };
assign v$_1025_out0 = { v$A$SAVED_6683_out0,v$A_11272_out0 };
assign v$R0_1143_out0 = v$G79_8390_out0;
assign v$PIN_1702_out0 = v$DIN_977_out0;
assign v$PIN_1703_out0 = v$DIN_978_out0;
assign v$B_2056_out0 = v$B_9458_out0;
assign v$B_2057_out0 = v$B_9459_out0;
assign v$_2415_out0 = v$_392_out0[1:0];
assign v$_2415_out1 = v$_392_out0[3:2];
assign v$_2416_out0 = v$_393_out0[1:0];
assign v$_2416_out1 = v$_393_out0[3:2];
assign v$SEL1_2433_out0 = v$A_11271_out0[15:15];
assign v$SEL1_2434_out0 = v$A_11272_out0[15:15];
assign v$IN_3016_out0 = v$IN_180_out0;
assign v$IN_3020_out0 = v$IN_181_out0;
assign v$A_6399_out0 = v$RM_12933_out0;
assign v$A_6400_out0 = v$RM_12934_out0;
assign v$DATAIN1_6590_out0 = v$DATA$IN1_10600_out0;
assign v$SEL9_6684_out0 = v$A_1951_out0[9:0];
assign v$SEL9_6685_out0 = v$A_1952_out0[9:0];
assign v$DATAIN0_7296_out0 = v$DATA$IN0_6953_out0;
assign v$SEL4_7649_out0 = v$DATA_3010_out0[7:0];
assign v$SEL4_7650_out0 = v$DATA_3011_out0[7:0];
assign v$SEL1_7748_out0 = v$DATA_3010_out0[11:0];
assign v$SEL1_7749_out0 = v$DATA_3011_out0[11:0];
assign v$SEL7_8117_out0 = v$A_11271_out0[9:0];
assign v$SEL7_8118_out0 = v$A_11272_out0[9:0];
assign v$_8844_out0 = v$_5930_out0[1:0];
assign v$_8844_out1 = v$_5930_out0[3:2];
assign v$_8845_out0 = v$_5931_out0[1:0];
assign v$_8845_out1 = v$_5931_out0[3:2];
assign v$A_9334_out0 = v$A_11271_out0;
assign v$A_9336_out0 = v$A_1951_out0;
assign v$A_9338_out0 = v$A_11272_out0;
assign v$A_9340_out0 = v$A_1952_out0;
assign v$MUX6_9803_out0 = v$SEL2_6423_out0 ? v$INT1_13185_out0 : v$INT0_11100_out0;
assign v$MUX6_9804_out0 = v$SEL2_6424_out0 ? v$INT1_13186_out0 : v$INT0_11101_out0;
assign v$_10329_out0 = v$_2854_out0[1:0];
assign v$_10329_out1 = v$_2854_out0[3:2];
assign v$_10330_out0 = v$_2855_out0[1:0];
assign v$_10330_out1 = v$_2855_out0[3:2];
assign v$THRESHOLD_10815_out0 = v$DATA_3010_out0;
assign v$THRESHOLD_10816_out0 = v$DATA_3011_out0;
assign v$SEL11_10831_out0 = v$A_1951_out0[15:15];
assign v$SEL11_10832_out0 = v$A_1952_out0[15:15];
assign v$_11044_out0 = { v$A$SAVED_10000_out0,v$A_1951_out0 };
assign v$_11045_out0 = { v$A$SAVED_10001_out0,v$A_1952_out0 };
assign v$_11387_out0 = v$_2507_out0[1:0];
assign v$_11387_out1 = v$_2507_out0[3:2];
assign v$_11388_out0 = v$_2508_out0[1:0];
assign v$_11388_out1 = v$_2508_out0[3:2];
assign v$SEL13_12388_out0 = v$A_1951_out0[15:15];
assign v$SEL13_12389_out0 = v$A_1952_out0[15:15];
assign v$R1_12676_out0 = v$G36_11766_out0;
assign v$SEL1_12970_out0 = v$DIN_977_out0[3:0];
assign v$SEL1_12971_out0 = v$DIN_978_out0[3:0];
assign v$MODE_44_out0 = v$SEL4_7649_out0;
assign v$MODE_45_out0 = v$SEL4_7650_out0;
assign v$_266_out0 = v$_8844_out0[0:0];
assign v$_266_out1 = v$_8844_out0[1:1];
assign v$_267_out0 = v$_8845_out0[0:0];
assign v$_267_out1 = v$_8845_out0[1:1];
assign v$_879_out0 = { v$C6_757_out0,v$SEL7_8117_out0 };
assign v$_880_out0 = { v$C6_758_out0,v$SEL7_8118_out0 };
assign v$_1158_out0 = { v$C8_5698_out0,v$SEL9_6684_out0 };
assign v$_1159_out0 = { v$C8_5699_out0,v$SEL9_6685_out0 };
assign v$G59_1484_out0 = v$PHALT_10440_out0 && v$R1_12676_out0;
assign v$A$32BIT_1751_out0 = v$_11044_out0;
assign v$A$32BIT_1752_out0 = v$_11045_out0;
assign v$_1868_out0 = v$_11387_out1[0:0];
assign v$_1868_out1 = v$_11387_out1[1:1];
assign v$_1869_out0 = v$_11388_out1[0:0];
assign v$_1869_out1 = v$_11388_out1[1:1];
assign v$MUX4_2551_out0 = v$G68_10170_out0 ? v$REG10_11541_out0 : v$DATAIN0_7296_out0;
assign v$_2736_out0 = v$_2415_out0[0:0];
assign v$_2736_out1 = v$_2415_out0[1:1];
assign v$_2737_out0 = v$_2416_out0[0:0];
assign v$_2737_out1 = v$_2416_out0[1:1];
assign v$_3284_out0 = v$_8844_out1[0:0];
assign v$_3284_out1 = v$_8844_out1[1:1];
assign v$_3285_out0 = v$_8845_out1[0:0];
assign v$_3285_out1 = v$_8845_out1[1:1];
assign v$_3651_out0 = v$_10329_out1[0:0];
assign v$_3651_out1 = v$_10329_out1[1:1];
assign v$_3652_out0 = v$_10330_out1[0:0];
assign v$_3652_out1 = v$_10330_out1[1:1];
assign {v$A1_4421_out1,v$A1_4421_out0 } = v$XOR1_3455_out0 + v$A_6399_out0 + v$SUBEN_8502_out0;
assign {v$A1_4422_out1,v$A1_4422_out0 } = v$XOR1_3456_out0 + v$A_6400_out0 + v$SUBEN_8503_out0;
assign v$R0_4666_out0 = v$R0_1143_out0;
assign v$SEL1_5086_out0 = v$A_9334_out0[14:10];
assign v$SEL1_5088_out0 = v$A_9336_out0[14:10];
assign v$SEL1_5090_out0 = v$A_9338_out0[14:10];
assign v$SEL1_5092_out0 = v$A_9340_out0[14:10];
assign v$_5418_out0 = v$PIN_1702_out0[7:0];
assign v$_5418_out1 = v$PIN_1702_out0[15:8];
assign v$_5419_out0 = v$PIN_1703_out0[7:0];
assign v$_5419_out1 = v$PIN_1703_out0[15:8];
assign v$IN_6532_out0 = v$IN_3016_out0;
assign v$IN_6536_out0 = v$IN_3020_out0;
assign v$_6815_out0 = v$_2415_out1[0:0];
assign v$_6815_out1 = v$_2415_out1[1:1];
assign v$_6816_out0 = v$_2416_out1[0:0];
assign v$_6816_out1 = v$_2416_out1[1:1];
assign v$MUX5_7180_out0 = v$G69_11035_out0 ? v$REG11_6578_out0 : v$DATAIN1_6590_out0;
assign v$_7294_out0 = v$_10329_out0[0:0];
assign v$_7294_out1 = v$_10329_out0[1:1];
assign v$_7295_out0 = v$_10330_out0[0:0];
assign v$_7295_out1 = v$_10330_out0[1:1];
assign v$R1_7681_out0 = v$R1_12676_out0;
assign v$G1_10445_out0 = ! v$SEL5_260_out0;
assign v$G1_10446_out0 = ! v$SEL5_261_out0;
assign v$_11630_out0 = v$_11387_out0[0:0];
assign v$_11630_out1 = v$_11387_out0[1:1];
assign v$_11631_out0 = v$_11388_out0[0:0];
assign v$_11631_out1 = v$_11388_out0[1:1];
assign v$MUX5_12042_out0 = v$SEL3_12208_out0 ? v$MUX7_435_out0 : v$MUX6_9803_out0;
assign v$MUX5_12043_out0 = v$SEL3_12209_out0 ? v$MUX7_436_out0 : v$MUX6_9804_out0;
assign v$B_12100_out0 = v$B_2056_out0;
assign v$B_12101_out0 = v$B_2057_out0;
assign v$B_12845_out0 = v$B_2056_out0;
assign v$B_12846_out0 = v$B_2057_out0;
assign v$A$32$BIT_13121_out0 = v$_1024_out0;
assign v$A$32$BIT_13122_out0 = v$_1025_out0;
assign v$A$EXP_236_out0 = v$SEL1_5086_out0;
assign v$A$EXP_238_out0 = v$SEL1_5088_out0;
assign v$A$EXP_240_out0 = v$SEL1_5090_out0;
assign v$A$EXP_242_out0 = v$SEL1_5092_out0;
assign v$_485_out0 = v$IN_6532_out0[0:0];
assign v$_486_out0 = v$IN_6536_out0[0:0];
assign v$G6_2205_out0 = v$R0_4666_out0 && v$R1_7681_out0;
assign v$_3209_out0 = v$IN_6532_out0[14:0];
assign v$_3213_out0 = v$IN_6536_out0[14:0];
assign v$SEL2_4179_out0 = v$B_12100_out0[14:0];
assign v$SEL2_4180_out0 = v$B_12101_out0[14:0];
assign v$_5001_out0 = { v$_1158_out0,v$C2_465_out0 };
assign v$_5002_out0 = { v$_1159_out0,v$C2_466_out0 };
assign v$8LSB_5144_out0 = v$_5418_out0;
assign v$8LSB_5145_out0 = v$_5419_out0;
assign v$COUT_5766_out0 = v$A1_4421_out1;
assign v$COUT_5767_out0 = v$A1_4422_out1;
assign v$SUM_6865_out0 = v$A1_4421_out0;
assign v$SUM_6866_out0 = v$A1_4422_out0;
assign v$_6962_out0 = v$IN_6532_out0[15:15];
assign v$_6963_out0 = v$IN_6536_out0[15:15];
assign v$EQ1_7467_out0 = v$A$32$BIT_13121_out0 == 32'h0;
assign v$EQ1_7468_out0 = v$A$32$BIT_13122_out0 == 32'h0;
assign v$G62_7744_out0 = v$G59_1484_out0 && v$PCHALT_11644_out0;
assign v$B_7913_out0 = v$B_12845_out0;
assign v$B_7914_out0 = v$B_12846_out0;
assign v$END_8367_out0 = v$_5418_out1;
assign v$END_8368_out0 = v$_5419_out1;
assign v$SEL4_8615_out0 = v$A$32BIT_1751_out0[22:0];
assign v$SEL4_8616_out0 = v$A$32BIT_1752_out0[22:0];
assign v$_8852_out0 = v$IN_6532_out0[0:0];
assign v$_8855_out0 = v$IN_6536_out0[0:0];
assign v$A_9335_out0 = v$A$32$BIT_13121_out0;
assign v$A_9337_out0 = v$A$32BIT_1751_out0;
assign v$A_9339_out0 = v$A$32$BIT_13122_out0;
assign v$A_9341_out0 = v$A$32BIT_1752_out0;
assign v$EQ3_9693_out0 = v$A$32$BIT_13121_out0 == 32'h0;
assign v$EQ3_9694_out0 = v$A$32$BIT_13122_out0 == 32'h0;
assign v$SEL6_9839_out0 = v$B_12100_out0[15:15];
assign v$SEL6_9840_out0 = v$B_12101_out0[15:15];
assign v$_9976_out0 = v$IN_6532_out0[15:1];
assign v$_9980_out0 = v$IN_6536_out0[15:1];
assign v$_10002_out0 = v$IN_6532_out0[15:1];
assign v$_10006_out0 = v$IN_6536_out0[15:1];
assign v$_11794_out0 = v$IN_6532_out0[15:1];
assign v$_11798_out0 = v$IN_6536_out0[15:1];
assign v$SEL8_12288_out0 = v$A$32$BIT_13121_out0[22:0];
assign v$SEL8_12289_out0 = v$A$32$BIT_13122_out0[22:0];
assign v$MODE_12630_out0 = v$MODE_44_out0;
assign v$MODE_12631_out0 = v$MODE_45_out0;
assign v$_709_out0 = { v$C1_5478_out0,v$_3209_out0 };
assign v$_713_out0 = { v$C1_5482_out0,v$_3213_out0 };
assign v$G3_2662_out0 = ! v$SEL6_9839_out0;
assign v$G3_2663_out0 = ! v$SEL6_9840_out0;
assign v$B_3230_out0 = v$B_7913_out0;
assign v$B_3234_out0 = v$B_7914_out0;
assign v$RMN_4169_out0 = v$SUM_6865_out0;
assign v$RMN_4170_out0 = v$SUM_6866_out0;
assign v$MUX8_4811_out0 = v$IS$32$BITS_527_out0 ? v$SEL8_12288_out0 : v$_879_out0;
assign v$MUX8_4812_out0 = v$IS$32$BITS_528_out0 ? v$SEL8_12289_out0 : v$_880_out0;
assign v$SEL1_5087_out0 = v$A_9335_out0[30:23];
assign v$SEL1_5089_out0 = v$A_9337_out0[30:23];
assign v$SEL1_5091_out0 = v$A_9339_out0[30:23];
assign v$SEL1_5093_out0 = v$A_9341_out0[30:23];
assign v$SEL5_5338_out0 = v$B_7913_out0[9:0];
assign v$SEL5_5339_out0 = v$B_7914_out0[9:0];
assign v$_5706_out0 = v$8LSB_5144_out0[3:0];
assign v$_5706_out1 = v$8LSB_5144_out0[7:4];
assign v$_5707_out0 = v$8LSB_5145_out0[3:0];
assign v$_5707_out1 = v$8LSB_5145_out0[7:4];
assign v$_6441_out0 = { v$_11794_out0,v$LSB_5342_out0 };
assign v$_6445_out0 = { v$_11798_out0,v$LSB_5343_out0 };
assign v$MODE_7108_out0 = v$MODE_12630_out0;
assign v$MODE_7109_out0 = v$MODE_12631_out0;
assign v$A_7350_out0 = v$A$EXP_236_out0;
assign v$A_7362_out0 = v$A$EXP_238_out0;
assign v$A_7366_out0 = v$A$EXP_240_out0;
assign v$A_7378_out0 = v$A$EXP_242_out0;
assign v$_8159_out0 = { v$B$SAVED_2592_out0,v$B_7913_out0 };
assign v$_8160_out0 = { v$B$SAVED_2593_out0,v$B_7914_out0 };
assign v$HALTVALID_8869_out0 = v$G6_2205_out0;
assign v$_8877_out0 = { v$_9976_out0,v$_8852_out0 };
assign v$_8881_out0 = { v$_9980_out0,v$_8855_out0 };
assign v$SEL2_9004_out0 = v$B_7913_out0[15:15];
assign v$SEL2_9005_out0 = v$B_7914_out0[15:15];
assign v$MUX6_9277_out0 = v$S$FF_7118_out0 ? v$LSB_5342_out0 : v$_6962_out0;
assign v$MUX6_9278_out0 = v$S$FF_7119_out0 ? v$LSB_5343_out0 : v$_6963_out0;
assign v$DM1_11395_out0 = v$HALTSEL_10098_out0 ? 1'h0 : v$G6_2205_out0;
assign v$DM1_11395_out1 = v$HALTSEL_10098_out0 ? v$G6_2205_out0 : 1'h0;
assign v$HALT_11481_out0 = v$G6_2205_out0;
assign v$MUX5_12110_out0 = v$S_7016_out0 ? v$_485_out0 : v$C2_1568_out0;
assign v$MUX5_12111_out0 = v$S_7017_out0 ? v$_486_out0 : v$C2_1569_out0;
assign v$_12560_out0 = { v$SEL4_8615_out0,v$C3_3631_out0 };
assign v$_12561_out0 = { v$SEL4_8616_out0,v$C3_3632_out0 };
assign v$A$EXP_237_out0 = v$SEL1_5087_out0;
assign v$A$EXP_239_out0 = v$SEL1_5089_out0;
assign v$A$EXP_241_out0 = v$SEL1_5091_out0;
assign v$A$EXP_243_out0 = v$SEL1_5093_out0;
assign v$_885_out0 = v$_5706_out0[1:0];
assign v$_885_out1 = v$_5706_out0[3:2];
assign v$_886_out0 = v$_5707_out0[1:0];
assign v$_886_out1 = v$_5707_out0[3:2];
assign v$B$32$BIT_1046_out0 = v$_8159_out0;
assign v$B$32$BIT_1047_out0 = v$_8160_out0;
assign v$MUX1_1505_out0 = v$G15_13187_out0 ? v$RMN_4169_out0 : v$RM_12933_out0;
assign v$MUX1_1506_out0 = v$G15_13188_out0 ? v$RMN_4170_out0 : v$RM_12934_out0;
assign v$MUX8_3643_out0 = v$IS$32$BIT_7152_out0 ? v$_12560_out0 : v$_5001_out0;
assign v$MUX8_3644_out0 = v$IS$32$BIT_7153_out0 ? v$_12561_out0 : v$_5002_out0;
assign v$SEL2_4733_out0 = v$B_3230_out0[14:10];
assign v$SEL2_4737_out0 = v$B_3234_out0[14:10];
assign v$HALT1_4838_out0 = v$DM1_11395_out1;
assign v$SEL4_4932_out0 = v$A_7350_out0[1:1];
assign v$SEL4_4941_out0 = v$A_7362_out0[1:1];
assign v$SEL4_4944_out0 = v$A_7366_out0[1:1];
assign v$SEL4_4953_out0 = v$A_7378_out0[1:1];
assign v$HALTVALID_5289_out0 = v$HALTVALID_8869_out0;
assign v$SEL3_5880_out0 = v$A_7350_out0[2:2];
assign v$SEL3_5889_out0 = v$A_7362_out0[2:2];
assign v$SEL3_5892_out0 = v$A_7366_out0[2:2];
assign v$SEL3_5901_out0 = v$A_7378_out0[2:2];
assign v$G7_6617_out0 = ! v$DM1_11395_out0;
assign v$HALT0_7510_out0 = v$DM1_11395_out0;
assign v$_7608_out0 = { v$_10002_out0,v$MUX6_9277_out0 };
assign v$_7612_out0 = { v$_10006_out0,v$MUX6_9278_out0 };
assign v$A$MANTISA_7625_out0 = v$MUX8_4811_out0;
assign v$A$MANTISA_7626_out0 = v$MUX8_4812_out0;
assign v$SEL5_8430_out0 = v$A_7350_out0[0:0];
assign v$SEL5_8439_out0 = v$A_7362_out0[0:0];
assign v$SEL5_8442_out0 = v$A_7366_out0[0:0];
assign v$SEL5_8451_out0 = v$A_7378_out0[0:0];
assign v$_8764_out0 = v$_5706_out1[1:0];
assign v$_8764_out1 = v$_5706_out1[3:2];
assign v$_8765_out0 = v$_5707_out1[1:0];
assign v$_8765_out1 = v$_5707_out1[3:2];
assign v$MUX4_11178_out0 = v$EN_12029_out0 ? v$_709_out0 : v$IN_6532_out0;
assign v$MUX4_11182_out0 = v$EN_12033_out0 ? v$_713_out0 : v$IN_6536_out0;
assign v$MUX10_11502_out0 = v$EQ1_11375_out0 ? v$G3_2662_out0 : v$SEL6_9839_out0;
assign v$MUX10_11503_out0 = v$EQ1_11376_out0 ? v$G3_2663_out0 : v$SEL6_9840_out0;
assign v$SEL2_11672_out0 = v$A_7350_out0[3:3];
assign v$SEL2_11681_out0 = v$A_7362_out0[3:3];
assign v$SEL2_11684_out0 = v$A_7366_out0[3:3];
assign v$SEL2_11693_out0 = v$A_7378_out0[3:3];
assign v$G1_12670_out0 = ((v$SEL1_2433_out0 && !v$SEL2_9004_out0) || (!v$SEL1_2433_out0) && v$SEL2_9004_out0);
assign v$G1_12671_out0 = ((v$SEL1_2434_out0 && !v$SEL2_9005_out0) || (!v$SEL1_2434_out0) && v$SEL2_9005_out0);
assign v$SEL1_12809_out0 = v$A_7350_out0[4:4];
assign v$SEL1_12810_out0 = v$A_7362_out0[4:4];
assign v$SEL1_12811_out0 = v$A_7366_out0[4:4];
assign v$SEL1_12812_out0 = v$A_7378_out0[4:4];
assign v$_12839_out0 = { v$C7_4039_out0,v$SEL5_5338_out0 };
assign v$_12840_out0 = { v$C7_4040_out0,v$SEL5_5339_out0 };
assign v$HALT0_290_out0 = v$HALT0_7510_out0;
assign v$_723_out0 = { v$SEL2_4179_out0,v$MUX10_11502_out0 };
assign v$_724_out0 = { v$SEL2_4180_out0,v$MUX10_11503_out0 };
assign v$A0_905_out0 = v$SEL5_8430_out0;
assign v$A0_914_out0 = v$SEL5_8439_out0;
assign v$A0_917_out0 = v$SEL5_8442_out0;
assign v$A0_926_out0 = v$SEL5_8451_out0;
assign v$EQ4_1767_out0 = v$B$32$BIT_1046_out0 == 32'h0;
assign v$EQ4_1768_out0 = v$B$32$BIT_1047_out0 == 32'h0;
assign v$_2193_out0 = v$_885_out0[0:0];
assign v$_2193_out1 = v$_885_out0[1:1];
assign v$_2194_out0 = v$_886_out0[0:0];
assign v$_2194_out1 = v$_886_out0[1:1];
assign v$A$MANTISA_2469_out0 = v$MUX8_3643_out0;
assign v$A$MANTISA_2470_out0 = v$MUX8_3644_out0;
assign v$HALT1_2849_out0 = v$HALT1_4838_out0;
assign v$SEL6_3085_out0 = v$B$32$BIT_1046_out0[22:0];
assign v$SEL6_3086_out0 = v$B$32$BIT_1047_out0[22:0];
assign v$B_3231_out0 = v$B$32$BIT_1046_out0;
assign v$B_3235_out0 = v$B$32$BIT_1047_out0;
assign v$A2_5564_out0 = v$SEL3_5880_out0;
assign v$A2_5573_out0 = v$SEL3_5889_out0;
assign v$A2_5576_out0 = v$SEL3_5892_out0;
assign v$A2_5585_out0 = v$SEL3_5901_out0;
assign v$_5597_out0 = v$_8764_out0[0:0];
assign v$_5597_out1 = v$_8764_out0[1:1];
assign v$_5598_out0 = v$_8765_out0[0:0];
assign v$_5598_out1 = v$_8765_out0[1:1];
assign v$_6383_out0 = v$_8764_out1[0:0];
assign v$_6383_out1 = v$_8764_out1[1:1];
assign v$_6384_out0 = v$_8765_out1[0:0];
assign v$_6384_out1 = v$_8765_out1[1:1];
assign v$A3_7018_out0 = v$SEL2_11672_out0;
assign v$A3_7027_out0 = v$SEL2_11681_out0;
assign v$A3_7030_out0 = v$SEL2_11684_out0;
assign v$A3_7039_out0 = v$SEL2_11693_out0;
assign v$A_7351_out0 = v$A$EXP_237_out0;
assign v$A_7363_out0 = v$A$EXP_239_out0;
assign v$A_7367_out0 = v$A$EXP_241_out0;
assign v$A_7379_out0 = v$A$EXP_243_out0;
assign v$MUX2_7822_out0 = v$G3_1507_out0 ? v$_6441_out0 : v$MUX4_11178_out0;
assign v$MUX2_7826_out0 = v$G3_1511_out0 ? v$_6445_out0 : v$MUX4_11182_out0;
assign v$SIGN_8414_out0 = v$G1_12670_out0;
assign v$SIGN_8415_out0 = v$G1_12671_out0;
assign v$_9417_out0 = v$MUX1_1505_out0[11:0];
assign v$_9417_out1 = v$MUX1_1505_out0[15:4];
assign v$_9418_out0 = v$MUX1_1506_out0[11:0];
assign v$_9418_out1 = v$MUX1_1506_out0[15:4];
assign v$_9470_out0 = v$_885_out1[0:0];
assign v$_9470_out1 = v$_885_out1[1:1];
assign v$_9471_out0 = v$_886_out1[0:0];
assign v$_9471_out1 = v$_886_out1[1:1];
assign v$A1_9726_out0 = v$SEL4_4932_out0;
assign v$A1_9735_out0 = v$SEL4_4941_out0;
assign v$A1_9738_out0 = v$SEL4_4944_out0;
assign v$A1_9747_out0 = v$SEL4_4953_out0;
assign v$A4_10323_out0 = v$SEL1_12809_out0;
assign v$A4_10324_out0 = v$SEL1_12810_out0;
assign v$A4_10325_out0 = v$SEL1_12811_out0;
assign v$A4_10326_out0 = v$SEL1_12812_out0;
assign v$G8_10979_out0 = v$G7_6617_out0 && v$DM1_11395_out1;
assign v$EQ2_11320_out0 = v$B$32$BIT_1046_out0 == 32'h0;
assign v$EQ2_11321_out0 = v$B$32$BIT_1047_out0 == 32'h0;
assign v$B$EXP_11734_out0 = v$SEL2_4733_out0;
assign v$B$EXP_11738_out0 = v$SEL2_4737_out0;
assign v$A$MANTISA_12691_out0 = v$A$MANTISA_7625_out0;
assign v$A$MANTISA_12692_out0 = v$A$MANTISA_7626_out0;
assign v$SIGN_591_out0 = v$SIGN_8414_out0;
assign v$SIGN_592_out0 = v$SIGN_8414_out0;
assign v$SIGN_593_out0 = v$SIGN_8415_out0;
assign v$SIGN_594_out0 = v$SIGN_8415_out0;
assign v$HALT1_1859_out0 = v$HALT1_2849_out0;
assign v$HALT0_3824_out0 = v$HALT0_290_out0;
assign v$G72_3918_out0 = ! v$HALT0_290_out0;
assign v$G5_4215_out0 = v$EQ3_9693_out0 || v$EQ4_1767_out0;
assign v$G5_4216_out0 = v$EQ3_9694_out0 || v$EQ4_1768_out0;
assign v$MUX1_4667_out0 = v$G4_2746_out0 ? v$_7608_out0 : v$MUX2_7822_out0;
assign v$MUX1_4671_out0 = v$G4_2750_out0 ? v$_7612_out0 : v$MUX2_7826_out0;
assign v$SEL2_4734_out0 = v$B_3231_out0[30:23];
assign v$SEL2_4738_out0 = v$B_3235_out0[30:23];
assign v$G78_4825_out0 = ! v$HALT1_2849_out0;
assign v$SEL1_6851_out0 = v$A_7351_out0[3:0];
assign v$SEL1_6854_out0 = v$A_7363_out0[3:0];
assign v$SEL1_6855_out0 = v$A_7367_out0[3:0];
assign v$SEL1_6858_out0 = v$A_7379_out0[3:0];
assign v$MUX7_8395_out0 = v$IS$32$BITS_527_out0 ? v$SEL6_3085_out0 : v$_12839_out0;
assign v$MUX7_8396_out0 = v$IS$32$BITS_528_out0 ? v$SEL6_3086_out0 : v$_12840_out0;
assign v$A$MANTISSA_8789_out0 = v$A$MANTISA_2469_out0;
assign v$A$MANTISSA_8790_out0 = v$A$MANTISA_2470_out0;
assign v$G54_8868_out0 = v$RAMWEN1_7089_out0 && v$HALT1_2849_out0;
assign v$G50_8876_out0 = ! v$HALT1_2849_out0;
assign v$G63_9223_out0 = v$HALT0_290_out0 || v$HALT1_2849_out0;
assign v$HALT0_9525_out0 = v$HALT0_290_out0;
assign v$RAMADDRMUX_9758_out0 = v$_9417_out0;
assign v$RAMADDRMUX_9759_out0 = v$_9418_out0;
assign v$B_9807_out0 = v$B$EXP_11734_out0;
assign v$B_9823_out0 = v$B$EXP_11738_out0;
assign v$A$MANTISA_9937_out0 = v$A$MANTISA_12691_out0;
assign v$A$MANTISA_9938_out0 = v$A$MANTISA_12692_out0;
assign v$ADDRMSB_10339_out0 = v$_9417_out1;
assign v$ADDRMSB_10340_out0 = v$_9418_out1;
assign v$G45_10651_out0 = v$READ$REQUEST1_4462_out0 && v$HALT1_2849_out0;
assign v$G3_11192_out0 = v$EQ1_7467_out0 || v$EQ2_11320_out0;
assign v$G3_11193_out0 = v$EQ1_7468_out0 || v$EQ2_11321_out0;
assign v$SEL4_12149_out0 = v$A_7351_out0[7:4];
assign v$SEL4_12152_out0 = v$A_7363_out0[7:4];
assign v$SEL4_12153_out0 = v$A_7367_out0[7:4];
assign v$SEL4_12156_out0 = v$A_7379_out0[7:4];
assign v$G53_12287_out0 = v$RAMWEN0_11645_out0 && v$HALT0_290_out0;
assign v$B_12546_out0 = v$_723_out0;
assign v$B_12547_out0 = v$_724_out0;
assign v$HALT1_13013_out0 = v$HALT1_2849_out0;
assign v$G51_13389_out0 = v$READ$REQUEST0_7434_out0 && v$HALT0_290_out0;
assign v$SEL12_18_out0 = v$B_12546_out0[9:0];
assign v$SEL12_19_out0 = v$B_12547_out0[9:0];
assign v$SEL3_513_out0 = v$A$MANTISSA_8789_out0[23:12];
assign v$SEL3_514_out0 = v$A$MANTISSA_8790_out0[23:12];
assign v$HALT_531_out0 = v$G63_9223_out0;
assign v$MUX3_1098_out0 = v$G8_1036_out0 ? v$_8877_out0 : v$MUX1_4667_out0;
assign v$MUX3_1102_out0 = v$G8_1040_out0 ? v$_8881_out0 : v$MUX1_4671_out0;
assign v$ARBHALT0_1685_out0 = v$HALT0_3824_out0;
assign v$B$MANTISA_1763_out0 = v$MUX7_8395_out0;
assign v$B$MANTISA_1764_out0 = v$MUX7_8396_out0;
assign v$SEL1_1953_out0 = v$A$MANTISSA_8789_out0[11:0];
assign v$SEL1_1954_out0 = v$A$MANTISSA_8790_out0[11:0];
assign v$SEL7_2856_out0 = v$B_9807_out0[3:3];
assign v$SEL7_2868_out0 = v$B_9823_out0[3:3];
assign v$RAMADDRMUX_3221_out0 = v$RAMADDRMUX_9758_out0;
assign v$RAMADDRMUX_3222_out0 = v$RAMADDRMUX_9759_out0;
assign v$B_3232_out0 = v$B_12546_out0;
assign v$B_3236_out0 = v$B_12547_out0;
assign v$ARBHALT1_3700_out0 = v$HALT1_1859_out0;
assign v$SEL6_3825_out0 = v$B_9807_out0[4:4];
assign v$SEL6_3827_out0 = v$B_9823_out0[4:4];
assign v$G64_4444_out0 = v$G50_8876_out0 && v$R1_12676_out0;
assign v$G1_4931_out0 = ! v$HALT1_13013_out0;
assign v$G2_5639_out0 = ! v$HALT0_9525_out0;
assign v$SEL9_7128_out0 = v$B_9807_out0[1:1];
assign v$SEL9_7140_out0 = v$B_9823_out0[1:1];
assign v$A_7352_out0 = v$SEL4_12149_out0;
assign v$A_7353_out0 = v$SEL1_6851_out0;
assign v$A_7364_out0 = v$SEL4_12152_out0;
assign v$A_7365_out0 = v$SEL1_6854_out0;
assign v$A_7368_out0 = v$SEL4_12153_out0;
assign v$A_7369_out0 = v$SEL1_6855_out0;
assign v$A_7380_out0 = v$SEL4_12156_out0;
assign v$A_7381_out0 = v$SEL1_6858_out0;
assign v$SEL3_7684_out0 = v$A$MANTISA_9937_out0[22:0];
assign v$SEL3_7685_out0 = v$A$MANTISA_9938_out0[22:0];
assign v$SEL10_8248_out0 = v$B_9807_out0[0:0];
assign v$SEL10_8260_out0 = v$B_9823_out0[0:0];
assign v$SEL8_8559_out0 = v$B_9807_out0[2:2];
assign v$SEL8_8571_out0 = v$B_9823_out0[2:2];
assign v$SEL15_9174_out0 = v$B_12546_out0[15:15];
assign v$SEL15_9175_out0 = v$B_12547_out0[15:15];
assign v$G74_10988_out0 = v$REG4_7248_out0 && v$G72_3918_out0;
assign v$SEL1_10991_out0 = v$A$MANTISA_9937_out0[22:0];
assign v$SEL1_10992_out0 = v$A$MANTISA_9938_out0[22:0];
assign v$B$EXP_11735_out0 = v$SEL2_4734_out0;
assign v$B$EXP_11739_out0 = v$SEL2_4738_out0;
assign v$G77_12941_out0 = v$REG7_4199_out0 && v$G78_4825_out0;
assign v$_12980_out0 = { v$B$SAVED_3014_out0,v$B_12546_out0 };
assign v$_12981_out0 = { v$B$SAVED_3015_out0,v$B_12547_out0 };
assign v$RAMADDRMUX_347_out0 = v$RAMADDRMUX_3221_out0;
assign v$RAMADDRMUX_348_out0 = v$RAMADDRMUX_3222_out0;
assign v$G83_357_out0 = v$G74_10988_out0 && v$G87_3518_out0;
assign v$A_1452_out0 = v$SEL3_513_out0;
assign v$A_1453_out0 = v$SEL1_1953_out0;
assign v$A_1454_out0 = v$SEL3_514_out0;
assign v$A_1455_out0 = v$SEL1_1954_out0;
assign v$G3_1738_out0 = v$G1_4931_out0 && v$WR1_9723_out0;
assign v$OUT_1899_out0 = v$MUX3_1098_out0;
assign v$OUT_1903_out0 = v$MUX3_1102_out0;
assign v$B0_2348_out0 = v$SEL10_8248_out0;
assign v$B0_2360_out0 = v$SEL10_8260_out0;
assign v$B$MANTISA_2780_out0 = v$B$MANTISA_1763_out0;
assign v$B$MANTISA_2781_out0 = v$B$MANTISA_1764_out0;
assign v$G85_4217_out0 = v$G77_12941_out0 && v$G86_9099_out0;
assign v$SEL2_4735_out0 = v$B_3232_out0[14:10];
assign v$SEL2_4739_out0 = v$B_3236_out0[14:10];
assign v$SEL4_4933_out0 = v$A_7352_out0[1:1];
assign v$SEL4_4934_out0 = v$A_7353_out0[1:1];
assign v$SEL4_4942_out0 = v$A_7364_out0[1:1];
assign v$SEL4_4943_out0 = v$A_7365_out0[1:1];
assign v$SEL4_4945_out0 = v$A_7368_out0[1:1];
assign v$SEL4_4946_out0 = v$A_7369_out0[1:1];
assign v$SEL4_4954_out0 = v$A_7380_out0[1:1];
assign v$SEL4_4955_out0 = v$A_7381_out0[1:1];
assign v$HALT_5113_out0 = v$ARBHALT0_1685_out0;
assign v$HALT_5114_out0 = v$ARBHALT1_3700_out0;
assign v$SEL3_5881_out0 = v$A_7352_out0[2:2];
assign v$SEL3_5882_out0 = v$A_7353_out0[2:2];
assign v$SEL3_5890_out0 = v$A_7364_out0[2:2];
assign v$SEL3_5891_out0 = v$A_7365_out0[2:2];
assign v$SEL3_5893_out0 = v$A_7368_out0[2:2];
assign v$SEL3_5894_out0 = v$A_7369_out0[2:2];
assign v$SEL3_5902_out0 = v$A_7380_out0[2:2];
assign v$SEL3_5903_out0 = v$A_7381_out0[2:2];
assign v$SEL5_8431_out0 = v$A_7352_out0[0:0];
assign v$SEL5_8432_out0 = v$A_7353_out0[0:0];
assign v$SEL5_8440_out0 = v$A_7364_out0[0:0];
assign v$SEL5_8441_out0 = v$A_7365_out0[0:0];
assign v$SEL5_8443_out0 = v$A_7368_out0[0:0];
assign v$SEL5_8444_out0 = v$A_7369_out0[0:0];
assign v$SEL5_8452_out0 = v$A_7380_out0[0:0];
assign v$SEL5_8453_out0 = v$A_7381_out0[0:0];
assign v$G4_8791_out0 = v$G2_5639_out0 && v$WR0_546_out0;
assign v$G6_9184_out0 = ((v$SEL11_10831_out0 && !v$SEL15_9174_out0) || (!v$SEL11_10831_out0) && v$SEL15_9174_out0);
assign v$G6_9185_out0 = ((v$SEL11_10832_out0 && !v$SEL15_9175_out0) || (!v$SEL11_10832_out0) && v$SEL15_9175_out0);
assign v$B1_9617_out0 = v$SEL9_7128_out0;
assign v$B1_9629_out0 = v$SEL9_7140_out0;
assign v$B_9808_out0 = v$B$EXP_11735_out0;
assign v$B_9824_out0 = v$B$EXP_11739_out0;
assign v$_11393_out0 = { v$C10_6197_out0,v$SEL12_18_out0 };
assign v$_11394_out0 = { v$C10_6198_out0,v$SEL12_19_out0 };
assign v$SEL2_11673_out0 = v$A_7352_out0[3:3];
assign v$SEL2_11674_out0 = v$A_7353_out0[3:3];
assign v$SEL2_11682_out0 = v$A_7364_out0[3:3];
assign v$SEL2_11683_out0 = v$A_7365_out0[3:3];
assign v$SEL2_11685_out0 = v$A_7368_out0[3:3];
assign v$SEL2_11686_out0 = v$A_7369_out0[3:3];
assign v$SEL2_11694_out0 = v$A_7380_out0[3:3];
assign v$SEL2_11695_out0 = v$A_7381_out0[3:3];
assign v$B2_11696_out0 = v$SEL8_8559_out0;
assign v$B2_11708_out0 = v$SEL8_8571_out0;
assign v$B4_11979_out0 = v$SEL6_3825_out0;
assign v$B4_11981_out0 = v$SEL6_3827_out0;
assign v$B3_12638_out0 = v$SEL7_2856_out0;
assign v$B3_12650_out0 = v$SEL7_2868_out0;
assign v$G57_12731_out0 = v$G62_7744_out0 || v$G64_4444_out0;
assign v$B$32BIT_13139_out0 = v$_12980_out0;
assign v$B$32BIT_13140_out0 = v$_12981_out0;
assign v$G37_743_out0 = !((v$B4_11979_out0 && !v$A4_10323_out0) || (!v$B4_11979_out0) && v$A4_10323_out0);
assign v$G37_745_out0 = !((v$B4_11981_out0 && !v$A4_10325_out0) || (!v$B4_11981_out0) && v$A4_10325_out0);
assign v$A0_906_out0 = v$SEL5_8431_out0;
assign v$A0_907_out0 = v$SEL5_8432_out0;
assign v$A0_915_out0 = v$SEL5_8440_out0;
assign v$A0_916_out0 = v$SEL5_8441_out0;
assign v$A0_918_out0 = v$SEL5_8443_out0;
assign v$A0_919_out0 = v$SEL5_8444_out0;
assign v$A0_927_out0 = v$SEL5_8452_out0;
assign v$A0_928_out0 = v$SEL5_8453_out0;
assign v$G5_1570_out0 = v$G4_8791_out0 || v$G3_1738_out0;
assign v$HALT_1675_out0 = v$HALT_5113_out0;
assign v$HALT_1676_out0 = v$HALT_5114_out0;
assign v$G21_2224_out0 = ! v$B1_9617_out0;
assign v$G21_2236_out0 = ! v$B1_9629_out0;
assign v$G8_2439_out0 = !((v$A3_7018_out0 && !v$B3_12638_out0) || (!v$A3_7018_out0) && v$B3_12638_out0);
assign v$G8_2451_out0 = !((v$A3_7030_out0 && !v$B3_12650_out0) || (!v$A3_7030_out0) && v$B3_12650_out0);
assign v$IN_3017_out0 = v$OUT_1899_out0;
assign v$IN_3021_out0 = v$OUT_1903_out0;
assign v$IS$SUB_3087_out0 = v$G6_9184_out0;
assign v$IS$SUB_3088_out0 = v$G6_9185_out0;
assign v$B_3233_out0 = v$B$32BIT_13139_out0;
assign v$B_3237_out0 = v$B$32BIT_13140_out0;
assign v$B$MANTISA_3300_out0 = v$B$MANTISA_2780_out0;
assign v$B$MANTISA_3301_out0 = v$B$MANTISA_2781_out0;
assign v$G36_3923_out0 = !((v$B3_12638_out0 && !v$A3_7018_out0) || (!v$B3_12638_out0) && v$A3_7018_out0);
assign v$G36_3935_out0 = !((v$B3_12650_out0 && !v$A3_7030_out0) || (!v$B3_12650_out0) && v$A3_7030_out0);
assign v$G6_4554_out0 = ! v$B3_12638_out0;
assign v$G6_4566_out0 = ! v$B3_12650_out0;
assign v$SEL8_4873_out0 = v$B$32BIT_13139_out0[22:0];
assign v$SEL8_4874_out0 = v$B$32BIT_13140_out0[22:0];
assign v$G3_5062_out0 = !((v$A4_10323_out0 && !v$B4_11979_out0) || (!v$A4_10323_out0) && v$B4_11979_out0);
assign v$G3_5064_out0 = !((v$A4_10325_out0 && !v$B4_11981_out0) || (!v$A4_10325_out0) && v$B4_11981_out0);
assign v$G90_5561_out0 = v$PHALT0$PREV_5150_out0 || v$G83_357_out0;
assign v$A2_5565_out0 = v$SEL3_5881_out0;
assign v$A2_5566_out0 = v$SEL3_5882_out0;
assign v$A2_5574_out0 = v$SEL3_5890_out0;
assign v$A2_5575_out0 = v$SEL3_5891_out0;
assign v$A2_5577_out0 = v$SEL3_5893_out0;
assign v$A2_5578_out0 = v$SEL3_5894_out0;
assign v$A2_5586_out0 = v$SEL3_5902_out0;
assign v$A2_5587_out0 = v$SEL3_5903_out0;
assign v$SEL1_5590_out0 = v$A_1452_out0[7:0];
assign v$SEL1_5591_out0 = v$A_1453_out0[7:0];
assign v$SEL1_5592_out0 = v$A_1454_out0[7:0];
assign v$SEL1_5593_out0 = v$A_1455_out0[7:0];
assign v$G17_5670_out0 = !((v$A0_905_out0 && !v$B0_2348_out0) || (!v$A0_905_out0) && v$B0_2348_out0);
assign v$G17_5682_out0 = !((v$A0_917_out0 && !v$B0_2360_out0) || (!v$A0_917_out0) && v$B0_2360_out0);
assign v$SEL3_6295_out0 = v$B_9808_out0[7:4];
assign v$SEL3_6299_out0 = v$B_9824_out0[7:4];
assign v$A3_7019_out0 = v$SEL2_11673_out0;
assign v$A3_7020_out0 = v$SEL2_11674_out0;
assign v$A3_7028_out0 = v$SEL2_11682_out0;
assign v$A3_7029_out0 = v$SEL2_11683_out0;
assign v$A3_7031_out0 = v$SEL2_11685_out0;
assign v$A3_7032_out0 = v$SEL2_11686_out0;
assign v$A3_7040_out0 = v$SEL2_11694_out0;
assign v$A3_7041_out0 = v$SEL2_11695_out0;
assign v$G23_7948_out0 = ! v$B0_2348_out0;
assign v$G23_7960_out0 = ! v$B0_2360_out0;
assign v$G33_8722_out0 = !((v$A0_905_out0 && !v$B0_2348_out0) || (!v$A0_905_out0) && v$B0_2348_out0);
assign v$G33_8734_out0 = !((v$A0_917_out0 && !v$B0_2360_out0) || (!v$A0_917_out0) && v$B0_2360_out0);
assign v$G1_8792_out0 = ! v$B4_11979_out0;
assign v$G1_8794_out0 = ! v$B4_11981_out0;
assign v$G15_9195_out0 = !((v$A2_5564_out0 && !v$B2_11696_out0) || (!v$A2_5564_out0) && v$B2_11696_out0);
assign v$G15_9207_out0 = !((v$A2_5576_out0 && !v$B2_11708_out0) || (!v$A2_5576_out0) && v$B2_11708_out0);
assign v$A1_9727_out0 = v$SEL4_4933_out0;
assign v$A1_9728_out0 = v$SEL4_4934_out0;
assign v$A1_9736_out0 = v$SEL4_4942_out0;
assign v$A1_9737_out0 = v$SEL4_4943_out0;
assign v$A1_9739_out0 = v$SEL4_4945_out0;
assign v$A1_9740_out0 = v$SEL4_4946_out0;
assign v$A1_9748_out0 = v$SEL4_4954_out0;
assign v$A1_9749_out0 = v$SEL4_4955_out0;
assign v$G35_9911_out0 = !((v$A2_5564_out0 && !v$B2_11696_out0) || (!v$A2_5564_out0) && v$B2_11696_out0);
assign v$G35_9923_out0 = !((v$A2_5576_out0 && !v$B2_11708_out0) || (!v$A2_5576_out0) && v$B2_11708_out0);
assign v$RAM$ADDR_10549_out0 = v$RAMADDRMUX_347_out0;
assign v$RAM$ADDR_10550_out0 = v$RAMADDRMUX_348_out0;
assign v$_10645_out0 = { v$_11393_out0,v$C1_11126_out0 };
assign v$_10646_out0 = { v$_11394_out0,v$C1_11127_out0 };
assign v$G12_11546_out0 = ! v$B2_11696_out0;
assign v$G12_11558_out0 = ! v$B2_11708_out0;
assign v$B$EXP_11736_out0 = v$SEL2_4735_out0;
assign v$B$EXP_11740_out0 = v$SEL2_4739_out0;
assign v$G16_11911_out0 = !((v$A1_9726_out0 && !v$B1_9617_out0) || (!v$A1_9726_out0) && v$B1_9617_out0);
assign v$G16_11923_out0 = !((v$A1_9738_out0 && !v$B1_9629_out0) || (!v$A1_9738_out0) && v$B1_9629_out0);
assign v$G34_12121_out0 = !((v$A1_9726_out0 && !v$B1_9617_out0) || (!v$A1_9726_out0) && v$B1_9617_out0);
assign v$G34_12133_out0 = !((v$A1_9738_out0 && !v$B1_9629_out0) || (!v$A1_9738_out0) && v$B1_9629_out0);
assign v$SEL2_12242_out0 = v$B_9808_out0[3:0];
assign v$SEL2_12246_out0 = v$B_9824_out0[3:0];
assign v$G89_12562_out0 = v$G85_4217_out0 || v$PHALT1$PREV_4956_out0;
assign v$SELIN_12946_out0 = v$G57_12731_out0;
assign v$SEL3_13253_out0 = v$A_1452_out0[11:8];
assign v$SEL3_13254_out0 = v$A_1453_out0[11:8];
assign v$SEL3_13255_out0 = v$A_1454_out0[11:8];
assign v$SEL3_13256_out0 = v$A_1455_out0[11:8];
assign v$A4XNORB4_597_out0 = v$G3_5062_out0;
assign v$A4XNORB4_599_out0 = v$G3_5064_out0;
assign v$A0XNORB0_669_out0 = v$G17_5670_out0;
assign v$A0XNORB0_681_out0 = v$G17_5682_out0;
assign v$SEL4_1201_out0 = v$B$MANTISA_3300_out0[22:0];
assign v$SEL4_1202_out0 = v$B$MANTISA_3301_out0[22:0];
assign v$A2XNORB2_3125_out0 = v$G15_9195_out0;
assign v$A2XNORB2_3137_out0 = v$G15_9207_out0;
assign v$RAM$ADDR_4425_out0 = v$RAM$ADDR_10549_out0;
assign v$RAM$ADDR_4426_out0 = v$RAM$ADDR_10550_out0;
assign v$G5_4704_out0 = v$A3_7018_out0 && v$G6_4554_out0;
assign v$G5_4716_out0 = v$A3_7030_out0 && v$G6_4566_out0;
assign v$SEL2_4736_out0 = v$B_3233_out0[30:23];
assign v$SEL2_4740_out0 = v$B_3237_out0[30:23];
assign v$RAMADDRESS_4749_out0 = v$RAM$ADDR_10549_out0;
assign v$RAMADDRESS_4750_out0 = v$RAM$ADDR_10550_out0;
assign v$G38_4889_out0 = v$G33_8722_out0 && v$G34_12121_out0;
assign v$G38_4901_out0 = v$G33_8734_out0 && v$G34_12133_out0;
assign v$V0_5005_out0 = v$G90_5561_out0;
assign v$_5153_out0 = { v$SEL8_4873_out0,v$C6_775_out0 };
assign v$_5154_out0 = { v$SEL8_4874_out0,v$C6_776_out0 };
assign v$IN_6533_out0 = v$IN_3017_out0;
assign v$IN_6537_out0 = v$IN_3021_out0;
assign v$G20_6619_out0 = v$A1_9726_out0 && v$G21_2224_out0;
assign v$G20_6631_out0 = v$A1_9738_out0 && v$G21_2236_out0;
assign v$G2_6949_out0 = v$A4_10323_out0 && v$G1_8792_out0;
assign v$G2_6951_out0 = v$A4_10325_out0 && v$G1_8794_out0;
assign v$G25_7203_out0 = v$A0_905_out0 && v$G23_7948_out0;
assign v$G25_7215_out0 = v$A0_917_out0 && v$G23_7960_out0;
assign v$SEL2_7265_out0 = v$B$MANTISA_3300_out0[22:0];
assign v$SEL2_7266_out0 = v$B$MANTISA_3301_out0[22:0];
assign v$A_7354_out0 = v$SEL3_13253_out0;
assign v$A_7355_out0 = v$SEL1_5590_out0;
assign v$A_7358_out0 = v$SEL3_13254_out0;
assign v$A_7359_out0 = v$SEL1_5591_out0;
assign v$A_7370_out0 = v$SEL3_13255_out0;
assign v$A_7371_out0 = v$SEL1_5592_out0;
assign v$A_7374_out0 = v$SEL3_13256_out0;
assign v$A_7375_out0 = v$SEL1_5593_out0;
assign v$B_9809_out0 = v$SEL3_6295_out0;
assign v$B_9810_out0 = v$SEL2_12242_out0;
assign v$B_9819_out0 = v$B$EXP_11736_out0;
assign v$B_9825_out0 = v$SEL3_6299_out0;
assign v$B_9826_out0 = v$SEL2_12246_out0;
assign v$B_9835_out0 = v$B$EXP_11740_out0;
assign v$A3XNORB3_10072_out0 = v$G8_2439_out0;
assign v$A3XNORB3_10084_out0 = v$G8_2451_out0;
assign v$IS$SUB_10742_out0 = v$IS$SUB_3087_out0;
assign v$IS$SUB_10743_out0 = v$IS$SUB_3088_out0;
assign v$G11_10906_out0 = v$A2_5564_out0 && v$G12_11546_out0;
assign v$G11_10918_out0 = v$A2_5576_out0 && v$G12_11558_out0;
assign v$MUX2_11061_out0 = v$SELIN_12946_out0 ? v$MUX5_7180_out0 : v$MUX4_2551_out0;
assign v$ADDRESS_11116_out0 = v$RAM$ADDR_10549_out0;
assign v$ADDRESS_11117_out0 = v$RAM$ADDR_10550_out0;
assign v$A1XNORB1_11225_out0 = v$G16_11911_out0;
assign v$A1XNORB1_11237_out0 = v$G16_11923_out0;
assign v$V1_11769_out0 = v$G89_12562_out0;
assign v$G39_12167_out0 = v$G36_3923_out0 && v$G37_743_out0;
assign v$G39_12169_out0 = v$G36_3935_out0 && v$G37_745_out0;
assign v$HALT_12505_out0 = v$HALT_1675_out0;
assign v$HALT_12506_out0 = v$HALT_1676_out0;
assign v$MEMHALT_12595_out0 = v$HALT_1675_out0;
assign v$MEMHALT_12596_out0 = v$HALT_1676_out0;
assign v$MUX5_815_out0 = v$IS$32$BIT_7152_out0 ? v$_5153_out0 : v$_10645_out0;
assign v$MUX5_816_out0 = v$IS$32$BIT_7153_out0 ? v$_5154_out0 : v$_10646_out0;
assign v$G7_1164_out0 = v$A4XNORB4_597_out0 && v$G5_4704_out0;
assign v$G7_1166_out0 = v$A4XNORB4_599_out0 && v$G5_4716_out0;
assign v$SEL7_2857_out0 = v$B_9809_out0[3:3];
assign v$SEL7_2858_out0 = v$B_9810_out0[3:3];
assign v$SEL7_2865_out0 = v$B_9819_out0[3:3];
assign v$SEL7_2869_out0 = v$B_9825_out0[3:3];
assign v$SEL7_2870_out0 = v$B_9826_out0[3:3];
assign v$SEL7_2877_out0 = v$B_9835_out0[3:3];
assign v$G13_3054_out0 = v$A3XNORB3_10072_out0 && v$G11_10906_out0;
assign v$G13_3066_out0 = v$A3XNORB3_10084_out0 && v$G11_10918_out0;
assign v$_3210_out0 = v$IN_6533_out0[13:0];
assign v$_3214_out0 = v$IN_6537_out0[13:0];
assign v$SEL6_3826_out0 = v$B_9819_out0[4:4];
assign v$SEL6_3828_out0 = v$B_9835_out0[4:4];
assign v$ADDRESS_3831_out0 = v$ADDRESS_11116_out0;
assign v$ADDRESS_3832_out0 = v$ADDRESS_11117_out0;
assign v$RAM$ADDR1_4451_out0 = v$RAM$ADDR_4426_out0;
assign v$SEL4_4935_out0 = v$A_7354_out0[1:1];
assign v$SEL4_4938_out0 = v$A_7358_out0[1:1];
assign v$SEL4_4947_out0 = v$A_7370_out0[1:1];
assign v$SEL4_4950_out0 = v$A_7374_out0[1:1];
assign v$A4$COMP$B4_4997_out0 = v$G2_6949_out0;
assign v$A4$COMP$B4_4999_out0 = v$G2_6951_out0;
assign v$SEL3_5883_out0 = v$A_7354_out0[2:2];
assign v$SEL3_5886_out0 = v$A_7358_out0[2:2];
assign v$SEL3_5895_out0 = v$A_7370_out0[2:2];
assign v$SEL3_5898_out0 = v$A_7374_out0[2:2];
assign v$VALID1_6051_out0 = v$V1_11769_out0;
assign v$SEL1_6852_out0 = v$A_7355_out0[3:0];
assign v$SEL1_6853_out0 = v$A_7359_out0[3:0];
assign v$SEL1_6856_out0 = v$A_7371_out0[3:0];
assign v$SEL1_6857_out0 = v$A_7375_out0[3:0];
assign v$SEL9_7129_out0 = v$B_9809_out0[1:1];
assign v$SEL9_7130_out0 = v$B_9810_out0[1:1];
assign v$SEL9_7137_out0 = v$B_9819_out0[1:1];
assign v$SEL9_7141_out0 = v$B_9825_out0[1:1];
assign v$SEL9_7142_out0 = v$B_9826_out0[1:1];
assign v$SEL9_7149_out0 = v$B_9835_out0[1:1];
assign v$_7576_out0 = v$IN_6533_out0[15:15];
assign v$_7577_out0 = v$IN_6537_out0[15:15];
assign v$RAM$ADDR0_8161_out0 = v$RAM$ADDR_4425_out0;
assign v$SEL10_8249_out0 = v$B_9809_out0[0:0];
assign v$SEL10_8250_out0 = v$B_9810_out0[0:0];
assign v$SEL10_8257_out0 = v$B_9819_out0[0:0];
assign v$SEL10_8261_out0 = v$B_9825_out0[0:0];
assign v$SEL10_8262_out0 = v$B_9826_out0[0:0];
assign v$SEL10_8269_out0 = v$B_9835_out0[0:0];
assign v$RAMADDRESS_8378_out0 = v$RAMADDRESS_4749_out0;
assign v$RAMADDRESS_8379_out0 = v$RAMADDRESS_4750_out0;
assign v$SEL5_8433_out0 = v$A_7354_out0[0:0];
assign v$SEL5_8436_out0 = v$A_7358_out0[0:0];
assign v$SEL5_8445_out0 = v$A_7370_out0[0:0];
assign v$SEL5_8448_out0 = v$A_7374_out0[0:0];
assign v$HALT_8544_out0 = v$HALT_12505_out0;
assign v$HALT_8545_out0 = v$HALT_12506_out0;
assign v$SEL8_8560_out0 = v$B_9809_out0[2:2];
assign v$SEL8_8561_out0 = v$B_9810_out0[2:2];
assign v$SEL8_8568_out0 = v$B_9819_out0[2:2];
assign v$SEL8_8572_out0 = v$B_9825_out0[2:2];
assign v$SEL8_8573_out0 = v$B_9826_out0[2:2];
assign v$SEL8_8580_out0 = v$B_9835_out0[2:2];
assign v$G28_8638_out0 = v$A1XNORB1_11225_out0 && v$G25_7203_out0;
assign v$G28_8650_out0 = v$A1XNORB1_11237_out0 && v$G25_7215_out0;
assign v$IS$SUB_8690_out0 = v$IS$SUB_10742_out0;
assign v$IS$SUB_8691_out0 = v$IS$SUB_10743_out0;
assign v$G22_8901_out0 = v$A2XNORB2_3125_out0 && v$G20_6619_out0;
assign v$G22_8913_out0 = v$A2XNORB2_3137_out0 && v$G20_6631_out0;
assign v$G40_8934_out0 = v$G35_9911_out0 && v$G39_12167_out0;
assign v$G40_8946_out0 = v$G35_9923_out0 && v$G39_12169_out0;
assign v$VALID0_8975_out0 = v$V0_5005_out0;
assign v$_9552_out0 = v$IN_6533_out0[1:0];
assign v$_9553_out0 = v$IN_6537_out0[1:0];
assign v$_9977_out0 = v$IN_6533_out0[15:2];
assign v$_9981_out0 = v$IN_6537_out0[15:2];
assign v$_10003_out0 = v$IN_6533_out0[15:2];
assign v$_10007_out0 = v$IN_6537_out0[15:2];
assign v$SEL2_11675_out0 = v$A_7354_out0[3:3];
assign v$SEL2_11678_out0 = v$A_7358_out0[3:3];
assign v$SEL2_11687_out0 = v$A_7370_out0[3:3];
assign v$SEL2_11690_out0 = v$A_7374_out0[3:3];
assign v$B$EXP_11737_out0 = v$SEL2_4736_out0;
assign v$B$EXP_11741_out0 = v$SEL2_4740_out0;
assign v$_11795_out0 = v$IN_6533_out0[15:2];
assign v$_11799_out0 = v$IN_6537_out0[15:2];
assign v$_12106_out0 = v$IN_6533_out0[1:0];
assign v$_12107_out0 = v$IN_6537_out0[1:0];
assign v$SEL4_12150_out0 = v$A_7355_out0[7:4];
assign v$SEL4_12151_out0 = v$A_7359_out0[7:4];
assign v$SEL4_12154_out0 = v$A_7371_out0[7:4];
assign v$SEL4_12155_out0 = v$A_7375_out0[7:4];
assign v$G28_13203_out0 = v$MEMHALT_12595_out0 || v$PIPELINEHALT_10164_out0;
assign v$G28_13204_out0 = v$MEMHALT_12596_out0 || v$PIPELINEHALT_10165_out0;
assign v$_710_out0 = { v$C1_5479_out0,v$_3210_out0 };
assign v$_714_out0 = { v$C1_5483_out0,v$_3214_out0 };
assign v$A0_908_out0 = v$SEL5_8433_out0;
assign v$A0_911_out0 = v$SEL5_8436_out0;
assign v$A0_920_out0 = v$SEL5_8445_out0;
assign v$A0_923_out0 = v$SEL5_8448_out0;
assign v$RAMAddress_1183_out0 = v$RAMADDRESS_8378_out0;
assign v$RAMAddress_1184_out0 = v$RAMADDRESS_8379_out0;
assign v$EQ1_1719_out0 = v$ADDRESS_3831_out0 == 12'hff8;
assign v$EQ1_1720_out0 = v$ADDRESS_3832_out0 == 12'hff8;
assign v$EQ5_2252_out0 = v$ADDRESS_3831_out0 == 12'hff7;
assign v$EQ5_2253_out0 = v$ADDRESS_3832_out0 == 12'hff7;
assign v$B0_2349_out0 = v$SEL10_8249_out0;
assign v$B0_2350_out0 = v$SEL10_8250_out0;
assign v$B0_2357_out0 = v$SEL10_8257_out0;
assign v$B0_2361_out0 = v$SEL10_8261_out0;
assign v$B0_2362_out0 = v$SEL10_8262_out0;
assign v$B0_2369_out0 = v$SEL10_8269_out0;
assign v$MUX3_2479_out0 = v$IS$SUB_8690_out0 ? v$C8_9178_out0 : v$C1_11389_out0;
assign v$MUX3_2480_out0 = v$IS$SUB_8691_out0 ? v$C8_9179_out0 : v$C1_11390_out0;
assign v$G27_3185_out0 = v$A2XNORB2_3125_out0 && v$G28_8638_out0;
assign v$G27_3197_out0 = v$A2XNORB2_3137_out0 && v$G28_8650_out0;
assign v$A3$COMP$B3_3338_out0 = v$G7_1164_out0;
assign v$A3$COMP$B3_3350_out0 = v$G7_1166_out0;
assign v$G18_3366_out0 = v$A3XNORB3_10072_out0 && v$G22_8901_out0;
assign v$G18_3378_out0 = v$A3XNORB3_10084_out0 && v$G22_8913_out0;
assign v$EXTHALT_4456_out0 = v$G28_13203_out0;
assign v$EXTHALT_4457_out0 = v$G28_13204_out0;
assign v$MUX5_5450_out0 = v$S_6988_out0 ? v$_9552_out0 : v$C1_1779_out0;
assign v$MUX5_5451_out0 = v$S_6989_out0 ? v$_9553_out0 : v$C1_1780_out0;
assign v$A2_5567_out0 = v$SEL3_5883_out0;
assign v$A2_5570_out0 = v$SEL3_5886_out0;
assign v$A2_5579_out0 = v$SEL3_5895_out0;
assign v$A2_5582_out0 = v$SEL3_5898_out0;
assign v$V0_6376_out0 = v$VALID0_8975_out0;
assign v$_6442_out0 = { v$_11795_out0,v$S$REG_2143_out0 };
assign v$_6446_out0 = { v$_11799_out0,v$S$REG_2144_out0 };
assign v$A3_7021_out0 = v$SEL2_11675_out0;
assign v$A3_7024_out0 = v$SEL2_11678_out0;
assign v$A3_7033_out0 = v$SEL2_11687_out0;
assign v$A3_7036_out0 = v$SEL2_11690_out0;
assign v$G41_7156_out0 = v$G38_4889_out0 && v$G40_8934_out0;
assign v$G41_7168_out0 = v$G38_4901_out0 && v$G40_8946_out0;
assign v$A_7356_out0 = v$SEL4_12150_out0;
assign v$A_7357_out0 = v$SEL1_6852_out0;
assign v$A_7360_out0 = v$SEL4_12151_out0;
assign v$A_7361_out0 = v$SEL1_6853_out0;
assign v$A_7372_out0 = v$SEL4_12154_out0;
assign v$A_7373_out0 = v$SEL1_6856_out0;
assign v$A_7376_out0 = v$SEL4_12155_out0;
assign v$A_7377_out0 = v$SEL1_6857_out0;
assign v$EQ3_7532_out0 = v$ADDRESS_3831_out0 == 12'hffa;
assign v$EQ3_7533_out0 = v$ADDRESS_3832_out0 == 12'hffa;
assign v$G14_8284_out0 = v$A4XNORB4_597_out0 && v$G13_3054_out0;
assign v$G14_8286_out0 = v$A4XNORB4_599_out0 && v$G13_3066_out0;
assign v$RAMADDR1_8300_out0 = v$RAM$ADDR1_4451_out0;
assign v$_8810_out0 = { v$_7576_out0,v$_7576_out0 };
assign v$_8811_out0 = { v$_7577_out0,v$_7577_out0 };
assign v$_8878_out0 = { v$_9977_out0,v$_12106_out0 };
assign v$_8882_out0 = { v$_9981_out0,v$_12107_out0 };
assign v$B1_9618_out0 = v$SEL9_7129_out0;
assign v$B1_9619_out0 = v$SEL9_7130_out0;
assign v$B1_9626_out0 = v$SEL9_7137_out0;
assign v$B1_9630_out0 = v$SEL9_7141_out0;
assign v$B1_9631_out0 = v$SEL9_7142_out0;
assign v$B1_9638_out0 = v$SEL9_7149_out0;
assign v$A1_9729_out0 = v$SEL4_4935_out0;
assign v$A1_9732_out0 = v$SEL4_4938_out0;
assign v$A1_9741_out0 = v$SEL4_4947_out0;
assign v$A1_9744_out0 = v$SEL4_4950_out0;
assign v$B_9820_out0 = v$B$EXP_11737_out0;
assign v$B_9836_out0 = v$B$EXP_11741_out0;
assign v$EQ12_10420_out0 = v$ADDRESS_3831_out0 == 12'hff6;
assign v$EQ12_10421_out0 = v$ADDRESS_3832_out0 == 12'hff6;
assign v$S_10768_out0 = v$HALT_8544_out0;
assign v$S_10769_out0 = v$HALT_8545_out0;
assign v$B$MANTISA_10857_out0 = v$MUX5_815_out0;
assign v$B$MANTISA_10858_out0 = v$MUX5_816_out0;
assign v$EQ4_11654_out0 = v$ADDRESS_3831_out0 == 12'hffb;
assign v$EQ4_11655_out0 = v$ADDRESS_3832_out0 == 12'hffb;
assign v$B2_11697_out0 = v$SEL8_8560_out0;
assign v$B2_11698_out0 = v$SEL8_8561_out0;
assign v$B2_11705_out0 = v$SEL8_8568_out0;
assign v$B2_11709_out0 = v$SEL8_8572_out0;
assign v$B2_11710_out0 = v$SEL8_8573_out0;
assign v$B2_11717_out0 = v$SEL8_8580_out0;
assign v$EQ2_11951_out0 = v$ADDRESS_3831_out0 == 12'hff9;
assign v$EQ2_11952_out0 = v$ADDRESS_3832_out0 == 12'hff9;
assign v$B4_11980_out0 = v$SEL6_3826_out0;
assign v$B4_11982_out0 = v$SEL6_3828_out0;
assign v$RAMADDR0_12041_out0 = v$RAM$ADDR0_8161_out0;
assign v$V1_12627_out0 = v$VALID1_6051_out0;
assign v$B3_12639_out0 = v$SEL7_2857_out0;
assign v$B3_12640_out0 = v$SEL7_2858_out0;
assign v$B3_12647_out0 = v$SEL7_2865_out0;
assign v$B3_12651_out0 = v$SEL7_2869_out0;
assign v$B3_12652_out0 = v$SEL7_2870_out0;
assign v$B3_12659_out0 = v$SEL7_2877_out0;
assign v$G65_12942_out0 = v$HALT_8544_out0 || v$G64_4407_out0;
assign v$G65_12943_out0 = v$HALT_8545_out0 || v$G64_4408_out0;
assign v$G13_186_out0 = v$EQ12_10420_out0 && v$WEN_2398_out0;
assign v$G13_187_out0 = v$EQ12_10421_out0 && v$WEN_2399_out0;
assign v$MUX6_542_out0 = v$FF1_11440_out0 ? v$S$REG_2143_out0 : v$_8810_out0;
assign v$MUX6_543_out0 = v$FF1_11441_out0 ? v$S$REG_2144_out0 : v$_8811_out0;
assign v$G37_744_out0 = !((v$B4_11980_out0 && !v$A4_10324_out0) || (!v$B4_11980_out0) && v$A4_10324_out0);
assign v$G37_746_out0 = !((v$B4_11982_out0 && !v$A4_10326_out0) || (!v$B4_11982_out0) && v$A4_10326_out0);
assign v$A2$COMP$B2_1115_out0 = v$G14_8284_out0;
assign v$A2$COMP$B2_1127_out0 = v$G14_8286_out0;
assign v$B$MANTISSA_1575_out0 = v$B$MANTISA_10857_out0;
assign v$B$MANTISSA_1576_out0 = v$B$MANTISA_10858_out0;
assign v$ADD_1721_out0 = v$RAMAddress_1183_out0;
assign v$ADD_1722_out0 = v$RAMAddress_1184_out0;
assign v$G21_2225_out0 = ! v$B1_9618_out0;
assign v$G21_2226_out0 = ! v$B1_9619_out0;
assign v$G21_2233_out0 = ! v$B1_9626_out0;
assign v$G21_2237_out0 = ! v$B1_9630_out0;
assign v$G21_2238_out0 = ! v$B1_9631_out0;
assign v$G21_2245_out0 = ! v$B1_9638_out0;
assign v$G8_2440_out0 = !((v$A3_7019_out0 && !v$B3_12639_out0) || (!v$A3_7019_out0) && v$B3_12639_out0);
assign v$G8_2441_out0 = !((v$A3_7020_out0 && !v$B3_12640_out0) || (!v$A3_7020_out0) && v$B3_12640_out0);
assign v$G8_2448_out0 = !((v$A3_7027_out0 && !v$B3_12647_out0) || (!v$A3_7027_out0) && v$B3_12647_out0);
assign v$G8_2452_out0 = !((v$A3_7031_out0 && !v$B3_12651_out0) || (!v$A3_7031_out0) && v$B3_12651_out0);
assign v$G8_2453_out0 = !((v$A3_7032_out0 && !v$B3_12652_out0) || (!v$A3_7032_out0) && v$B3_12652_out0);
assign v$G8_2460_out0 = !((v$A3_7039_out0 && !v$B3_12659_out0) || (!v$A3_7039_out0) && v$B3_12659_out0);
assign v$G30_3316_out0 = !(v$EXTHALT_4456_out0 || v$STPHALT_2988_out0);
assign v$G30_3317_out0 = !(v$EXTHALT_4457_out0 || v$STPHALT_2989_out0);
assign v$G36_3924_out0 = !((v$B3_12639_out0 && !v$A3_7019_out0) || (!v$B3_12639_out0) && v$A3_7019_out0);
assign v$G36_3925_out0 = !((v$B3_12640_out0 && !v$A3_7020_out0) || (!v$B3_12640_out0) && v$A3_7020_out0);
assign v$G36_3932_out0 = !((v$B3_12647_out0 && !v$A3_7027_out0) || (!v$B3_12647_out0) && v$A3_7027_out0);
assign v$G36_3936_out0 = !((v$B3_12651_out0 && !v$A3_7031_out0) || (!v$B3_12651_out0) && v$A3_7031_out0);
assign v$G36_3937_out0 = !((v$B3_12652_out0 && !v$A3_7032_out0) || (!v$B3_12652_out0) && v$A3_7032_out0);
assign v$G36_3944_out0 = !((v$B3_12659_out0 && !v$A3_7039_out0) || (!v$B3_12659_out0) && v$A3_7039_out0);
assign v$G6_4555_out0 = ! v$B3_12639_out0;
assign v$G6_4556_out0 = ! v$B3_12640_out0;
assign v$G6_4563_out0 = ! v$B3_12647_out0;
assign v$G6_4567_out0 = ! v$B3_12651_out0;
assign v$G6_4568_out0 = ! v$B3_12652_out0;
assign v$G6_4575_out0 = ! v$B3_12659_out0;
assign v$MUX6_4683_out0 = v$G70_9421_out0 ? v$REG12_2023_out0 : v$RAMADDR1_8300_out0;
assign v$SEL4_4936_out0 = v$A_7356_out0[1:1];
assign v$SEL4_4937_out0 = v$A_7357_out0[1:1];
assign v$SEL4_4939_out0 = v$A_7360_out0[1:1];
assign v$SEL4_4940_out0 = v$A_7361_out0[1:1];
assign v$SEL4_4948_out0 = v$A_7372_out0[1:1];
assign v$SEL4_4949_out0 = v$A_7373_out0[1:1];
assign v$SEL4_4951_out0 = v$A_7376_out0[1:1];
assign v$SEL4_4952_out0 = v$A_7377_out0[1:1];
assign v$G3_5063_out0 = !((v$A4_10324_out0 && !v$B4_11980_out0) || (!v$A4_10324_out0) && v$B4_11980_out0);
assign v$G3_5065_out0 = !((v$A4_10326_out0 && !v$B4_11982_out0) || (!v$A4_10326_out0) && v$B4_11982_out0);
assign v$G3_5080_out0 = v$EQ2_11951_out0 && v$WEN_2398_out0;
assign v$G3_5081_out0 = v$EQ2_11952_out0 && v$WEN_2399_out0;
assign v$S_5522_out0 = v$S_10768_out0;
assign v$S_5523_out0 = v$S_10769_out0;
assign v$G17_5671_out0 = !((v$A0_906_out0 && !v$B0_2349_out0) || (!v$A0_906_out0) && v$B0_2349_out0);
assign v$G17_5672_out0 = !((v$A0_907_out0 && !v$B0_2350_out0) || (!v$A0_907_out0) && v$B0_2350_out0);
assign v$G17_5679_out0 = !((v$A0_914_out0 && !v$B0_2357_out0) || (!v$A0_914_out0) && v$B0_2357_out0);
assign v$G17_5683_out0 = !((v$A0_918_out0 && !v$B0_2361_out0) || (!v$A0_918_out0) && v$B0_2361_out0);
assign v$G17_5684_out0 = !((v$A0_919_out0 && !v$B0_2362_out0) || (!v$A0_919_out0) && v$B0_2362_out0);
assign v$G17_5691_out0 = !((v$A0_926_out0 && !v$B0_2369_out0) || (!v$A0_926_out0) && v$B0_2369_out0);
assign v$SEL3_5884_out0 = v$A_7356_out0[2:2];
assign v$SEL3_5885_out0 = v$A_7357_out0[2:2];
assign v$SEL3_5887_out0 = v$A_7360_out0[2:2];
assign v$SEL3_5888_out0 = v$A_7361_out0[2:2];
assign v$SEL3_5896_out0 = v$A_7372_out0[2:2];
assign v$SEL3_5897_out0 = v$A_7373_out0[2:2];
assign v$SEL3_5899_out0 = v$A_7376_out0[2:2];
assign v$SEL3_5900_out0 = v$A_7377_out0[2:2];
assign v$G66_5924_out0 = ! v$G65_12942_out0;
assign v$G66_5925_out0 = ! v$G65_12943_out0;
assign v$SEL3_6298_out0 = v$B_9820_out0[7:4];
assign v$SEL3_6302_out0 = v$B_9836_out0[7:4];
assign v$MUX3_6357_out0 = v$G66_6177_out0 ? v$REG9_11269_out0 : v$RAMADDR0_12041_out0;
assign v$G19_6817_out0 = v$A4XNORB4_597_out0 && v$G18_3366_out0;
assign v$G19_6819_out0 = v$A4XNORB4_599_out0 && v$G18_3378_out0;
assign v$G23_7949_out0 = ! v$B0_2349_out0;
assign v$G23_7950_out0 = ! v$B0_2350_out0;
assign v$G23_7957_out0 = ! v$B0_2357_out0;
assign v$G23_7961_out0 = ! v$B0_2361_out0;
assign v$G23_7962_out0 = ! v$B0_2362_out0;
assign v$G23_7969_out0 = ! v$B0_2369_out0;
assign v$G5_8400_out0 = v$EQ5_2252_out0 && v$WEN_2398_out0;
assign v$G5_8401_out0 = v$EQ5_2253_out0 && v$WEN_2399_out0;
assign v$SEL5_8434_out0 = v$A_7356_out0[0:0];
assign v$SEL5_8435_out0 = v$A_7357_out0[0:0];
assign v$SEL5_8437_out0 = v$A_7360_out0[0:0];
assign v$SEL5_8438_out0 = v$A_7361_out0[0:0];
assign v$SEL5_8446_out0 = v$A_7372_out0[0:0];
assign v$SEL5_8447_out0 = v$A_7373_out0[0:0];
assign v$SEL5_8449_out0 = v$A_7376_out0[0:0];
assign v$SEL5_8450_out0 = v$A_7377_out0[0:0];
assign v$G33_8723_out0 = !((v$A0_906_out0 && !v$B0_2349_out0) || (!v$A0_906_out0) && v$B0_2349_out0);
assign v$G33_8724_out0 = !((v$A0_907_out0 && !v$B0_2350_out0) || (!v$A0_907_out0) && v$B0_2350_out0);
assign v$G33_8731_out0 = !((v$A0_914_out0 && !v$B0_2357_out0) || (!v$A0_914_out0) && v$B0_2357_out0);
assign v$G33_8735_out0 = !((v$A0_918_out0 && !v$B0_2361_out0) || (!v$A0_918_out0) && v$B0_2361_out0);
assign v$G33_8736_out0 = !((v$A0_919_out0 && !v$B0_2362_out0) || (!v$A0_919_out0) && v$B0_2362_out0);
assign v$G33_8743_out0 = !((v$A0_926_out0 && !v$B0_2369_out0) || (!v$A0_926_out0) && v$B0_2369_out0);
assign v$G1_8793_out0 = ! v$B4_11980_out0;
assign v$G1_8795_out0 = ! v$B4_11982_out0;
assign v$G15_9196_out0 = !((v$A2_5565_out0 && !v$B2_11697_out0) || (!v$A2_5565_out0) && v$B2_11697_out0);
assign v$G15_9197_out0 = !((v$A2_5566_out0 && !v$B2_11698_out0) || (!v$A2_5566_out0) && v$B2_11698_out0);
assign v$G15_9204_out0 = !((v$A2_5573_out0 && !v$B2_11705_out0) || (!v$A2_5573_out0) && v$B2_11705_out0);
assign v$G15_9208_out0 = !((v$A2_5577_out0 && !v$B2_11709_out0) || (!v$A2_5577_out0) && v$B2_11709_out0);
assign v$G15_9209_out0 = !((v$A2_5578_out0 && !v$B2_11710_out0) || (!v$A2_5578_out0) && v$B2_11710_out0);
assign v$G15_9216_out0 = !((v$A2_5585_out0 && !v$B2_11717_out0) || (!v$A2_5585_out0) && v$B2_11717_out0);
assign v$G2_9239_out0 = v$EQ3_7532_out0 && v$WEN_2398_out0;
assign v$G2_9240_out0 = v$EQ3_7533_out0 && v$WEN_2399_out0;
assign v$VALID_9883_out0 = v$V0_6376_out0;
assign v$VALID_9884_out0 = v$V1_12627_out0;
assign v$G35_9912_out0 = !((v$A2_5565_out0 && !v$B2_11697_out0) || (!v$A2_5565_out0) && v$B2_11697_out0);
assign v$G35_9913_out0 = !((v$A2_5566_out0 && !v$B2_11698_out0) || (!v$A2_5566_out0) && v$B2_11698_out0);
assign v$G35_9920_out0 = !((v$A2_5573_out0 && !v$B2_11705_out0) || (!v$A2_5573_out0) && v$B2_11705_out0);
assign v$G35_9924_out0 = !((v$A2_5577_out0 && !v$B2_11709_out0) || (!v$A2_5577_out0) && v$B2_11709_out0);
assign v$G35_9925_out0 = !((v$A2_5578_out0 && !v$B2_11710_out0) || (!v$A2_5578_out0) && v$B2_11710_out0);
assign v$G35_9932_out0 = !((v$A2_5585_out0 && !v$B2_11717_out0) || (!v$A2_5585_out0) && v$B2_11717_out0);
assign v$G4_10436_out0 = v$EQ1_1719_out0 && v$WEN_2398_out0;
assign v$G4_10437_out0 = v$EQ1_1720_out0 && v$WEN_2399_out0;
assign v$G24_10947_out0 = v$A3XNORB3_10072_out0 && v$G27_3185_out0;
assign v$G24_10959_out0 = v$A3XNORB3_10084_out0 && v$G27_3197_out0;
assign v$MUX4_11179_out0 = v$EN_12030_out0 ? v$_710_out0 : v$IN_6533_out0;
assign v$MUX4_11183_out0 = v$EN_12034_out0 ? v$_714_out0 : v$IN_6537_out0;
assign v$G12_11547_out0 = ! v$B2_11697_out0;
assign v$G12_11548_out0 = ! v$B2_11698_out0;
assign v$G12_11555_out0 = ! v$B2_11705_out0;
assign v$G12_11559_out0 = ! v$B2_11709_out0;
assign v$G12_11560_out0 = ! v$B2_11710_out0;
assign v$G12_11567_out0 = ! v$B2_11717_out0;
assign v$G1_11574_out0 = v$EQ4_11654_out0 && v$WEN_2398_out0;
assign v$G1_11575_out0 = v$EQ4_11655_out0 && v$WEN_2399_out0;
assign v$SEL2_11676_out0 = v$A_7356_out0[3:3];
assign v$SEL2_11677_out0 = v$A_7357_out0[3:3];
assign v$SEL2_11679_out0 = v$A_7360_out0[3:3];
assign v$SEL2_11680_out0 = v$A_7361_out0[3:3];
assign v$SEL2_11688_out0 = v$A_7372_out0[3:3];
assign v$SEL2_11689_out0 = v$A_7373_out0[3:3];
assign v$SEL2_11691_out0 = v$A_7376_out0[3:3];
assign v$SEL2_11692_out0 = v$A_7377_out0[3:3];
assign v$G16_11912_out0 = !((v$A1_9727_out0 && !v$B1_9618_out0) || (!v$A1_9727_out0) && v$B1_9618_out0);
assign v$G16_11913_out0 = !((v$A1_9728_out0 && !v$B1_9619_out0) || (!v$A1_9728_out0) && v$B1_9619_out0);
assign v$G16_11920_out0 = !((v$A1_9735_out0 && !v$B1_9626_out0) || (!v$A1_9735_out0) && v$B1_9626_out0);
assign v$G16_11924_out0 = !((v$A1_9739_out0 && !v$B1_9630_out0) || (!v$A1_9739_out0) && v$B1_9630_out0);
assign v$G16_11925_out0 = !((v$A1_9740_out0 && !v$B1_9631_out0) || (!v$A1_9740_out0) && v$B1_9631_out0);
assign v$G16_11932_out0 = !((v$A1_9747_out0 && !v$B1_9638_out0) || (!v$A1_9747_out0) && v$B1_9638_out0);
assign v$G34_12122_out0 = !((v$A1_9727_out0 && !v$B1_9618_out0) || (!v$A1_9727_out0) && v$B1_9618_out0);
assign v$G34_12123_out0 = !((v$A1_9728_out0 && !v$B1_9619_out0) || (!v$A1_9728_out0) && v$B1_9619_out0);
assign v$G34_12130_out0 = !((v$A1_9735_out0 && !v$B1_9626_out0) || (!v$A1_9735_out0) && v$B1_9626_out0);
assign v$G34_12134_out0 = !((v$A1_9739_out0 && !v$B1_9630_out0) || (!v$A1_9739_out0) && v$B1_9630_out0);
assign v$G34_12135_out0 = !((v$A1_9740_out0 && !v$B1_9631_out0) || (!v$A1_9740_out0) && v$B1_9631_out0);
assign v$G34_12142_out0 = !((v$A1_9747_out0 && !v$B1_9638_out0) || (!v$A1_9747_out0) && v$B1_9638_out0);
assign v$SEL2_12245_out0 = v$B_9820_out0[3:0];
assign v$SEL2_12249_out0 = v$B_9836_out0[3:0];
assign v$SAME_13351_out0 = v$G41_7156_out0;
assign v$SAME_13367_out0 = v$G41_7168_out0;
assign v$I3REGISTERWRITE_521_out0 = v$G1_11574_out0;
assign v$I3REGISTERWRITE_522_out0 = v$G1_11575_out0;
assign v$SEL4_589_out0 = v$B$MANTISSA_1575_out0[23:12];
assign v$SEL4_590_out0 = v$B$MANTISSA_1576_out0[23:12];
assign v$A4XNORB4_598_out0 = v$G3_5063_out0;
assign v$A4XNORB4_600_out0 = v$G3_5065_out0;
assign v$A0XNORB0_670_out0 = v$G17_5671_out0;
assign v$A0XNORB0_671_out0 = v$G17_5672_out0;
assign v$A0XNORB0_678_out0 = v$G17_5679_out0;
assign v$A0XNORB0_682_out0 = v$G17_5683_out0;
assign v$A0XNORB0_683_out0 = v$G17_5684_out0;
assign v$A0XNORB0_690_out0 = v$G17_5691_out0;
assign v$COUNTEREN_828_out0 = v$G13_186_out0;
assign v$COUNTEREN_829_out0 = v$G13_187_out0;
assign v$A0_909_out0 = v$SEL5_8434_out0;
assign v$A0_910_out0 = v$SEL5_8435_out0;
assign v$A0_912_out0 = v$SEL5_8437_out0;
assign v$A0_913_out0 = v$SEL5_8438_out0;
assign v$A0_921_out0 = v$SEL5_8446_out0;
assign v$A0_922_out0 = v$SEL5_8447_out0;
assign v$A0_924_out0 = v$SEL5_8449_out0;
assign v$A0_925_out0 = v$SEL5_8450_out0;
assign v$MUX1_1023_out0 = v$SELIN_12946_out0 ? v$MUX6_4683_out0 : v$MUX3_6357_out0;
assign v$I1REGISTERWRITE_1698_out0 = v$G3_5080_out0;
assign v$I1REGISTERWRITE_1699_out0 = v$G3_5081_out0;
assign v$I0REGISTERWRITE_2048_out0 = v$G4_10436_out0;
assign v$I0REGISTERWRITE_2049_out0 = v$G4_10437_out0;
assign v$ModeRegAdd_2724_out0 = v$ADD_1721_out0 == 12'hffc;
assign v$ModeRegAdd_2725_out0 = v$ADD_1722_out0 == 12'hffc;
assign v$A2XNORB2_3126_out0 = v$G15_9196_out0;
assign v$A2XNORB2_3127_out0 = v$G15_9197_out0;
assign v$A2XNORB2_3134_out0 = v$G15_9204_out0;
assign v$A2XNORB2_3138_out0 = v$G15_9208_out0;
assign v$A2XNORB2_3139_out0 = v$G15_9209_out0;
assign v$A2XNORB2_3146_out0 = v$G15_9216_out0;
assign v$MODEEN_3782_out0 = v$G5_8400_out0;
assign v$MODEEN_3783_out0 = v$G5_8401_out0;
assign v$G5_4705_out0 = v$A3_7019_out0 && v$G6_4555_out0;
assign v$G5_4706_out0 = v$A3_7020_out0 && v$G6_4556_out0;
assign v$G5_4713_out0 = v$A3_7027_out0 && v$G6_4563_out0;
assign v$G5_4717_out0 = v$A3_7031_out0 && v$G6_4567_out0;
assign v$G5_4718_out0 = v$A3_7032_out0 && v$G6_4568_out0;
assign v$G5_4725_out0 = v$A3_7039_out0 && v$G6_4575_out0;
assign v$G38_4890_out0 = v$G33_8723_out0 && v$G34_12122_out0;
assign v$G38_4891_out0 = v$G33_8724_out0 && v$G34_12123_out0;
assign v$G38_4898_out0 = v$G33_8731_out0 && v$G34_12130_out0;
assign v$G38_4902_out0 = v$G33_8735_out0 && v$G34_12134_out0;
assign v$G38_4903_out0 = v$G33_8736_out0 && v$G34_12135_out0;
assign v$G38_4910_out0 = v$G33_8743_out0 && v$G34_12142_out0;
assign v$StatRegAdd_5285_out0 = v$ADD_1721_out0 == 12'hffd;
assign v$StatRegAdd_5286_out0 = v$ADD_1722_out0 == 12'hffd;
assign v$A2_5568_out0 = v$SEL3_5884_out0;
assign v$A2_5569_out0 = v$SEL3_5885_out0;
assign v$A2_5571_out0 = v$SEL3_5887_out0;
assign v$A2_5572_out0 = v$SEL3_5888_out0;
assign v$A2_5580_out0 = v$SEL3_5896_out0;
assign v$A2_5581_out0 = v$SEL3_5897_out0;
assign v$A2_5583_out0 = v$SEL3_5899_out0;
assign v$A2_5584_out0 = v$SEL3_5900_out0;
assign v$EN_6318_out0 = v$G30_3316_out0;
assign v$EN_6319_out0 = v$G30_3317_out0;
assign v$G20_6620_out0 = v$A1_9727_out0 && v$G21_2225_out0;
assign v$G20_6621_out0 = v$A1_9728_out0 && v$G21_2226_out0;
assign v$G20_6628_out0 = v$A1_9735_out0 && v$G21_2233_out0;
assign v$G20_6632_out0 = v$A1_9739_out0 && v$G21_2237_out0;
assign v$G20_6633_out0 = v$A1_9740_out0 && v$G21_2238_out0;
assign v$G20_6640_out0 = v$A1_9747_out0 && v$G21_2245_out0;
assign v$G2_6950_out0 = v$A4_10324_out0 && v$G1_8793_out0;
assign v$G2_6952_out0 = v$A4_10326_out0 && v$G1_8795_out0;
assign v$A3_7022_out0 = v$SEL2_11676_out0;
assign v$A3_7023_out0 = v$SEL2_11677_out0;
assign v$A3_7025_out0 = v$SEL2_11679_out0;
assign v$A3_7026_out0 = v$SEL2_11680_out0;
assign v$A3_7034_out0 = v$SEL2_11688_out0;
assign v$A3_7035_out0 = v$SEL2_11689_out0;
assign v$A3_7037_out0 = v$SEL2_11691_out0;
assign v$A3_7038_out0 = v$SEL2_11692_out0;
assign v$G25_7204_out0 = v$A0_906_out0 && v$G23_7949_out0;
assign v$G25_7205_out0 = v$A0_907_out0 && v$G23_7950_out0;
assign v$G25_7212_out0 = v$A0_914_out0 && v$G23_7957_out0;
assign v$G25_7216_out0 = v$A0_918_out0 && v$G23_7961_out0;
assign v$G25_7217_out0 = v$A0_919_out0 && v$G23_7962_out0;
assign v$G25_7224_out0 = v$A0_926_out0 && v$G23_7969_out0;
assign v$G26_7414_out0 = v$A4XNORB4_597_out0 && v$G24_10947_out0;
assign v$G26_7416_out0 = v$A4XNORB4_599_out0 && v$G24_10959_out0;
assign v$_7609_out0 = { v$_10003_out0,v$MUX6_542_out0 };
assign v$_7613_out0 = { v$_10007_out0,v$MUX6_543_out0 };
assign v$I2REGISTERWRITE_7720_out0 = v$G2_9239_out0;
assign v$I2REGISTERWRITE_7721_out0 = v$G2_9240_out0;
assign v$MUX2_7823_out0 = v$G3_1508_out0 ? v$_6442_out0 : v$MUX4_11179_out0;
assign v$MUX2_7827_out0 = v$G3_1512_out0 ? v$_6446_out0 : v$MUX4_11183_out0;
assign v$A1$COMP$B1_8127_out0 = v$G19_6817_out0;
assign v$A1$COMP$B1_8139_out0 = v$G19_6819_out0;
assign v$RXRegAdd_8613_out0 = v$ADD_1721_out0 == 12'hffe;
assign v$RXRegAdd_8614_out0 = v$ADD_1722_out0 == 12'hffe;
assign v$G40_8935_out0 = v$G35_9912_out0 && v$G36_3924_out0;
assign v$G40_8936_out0 = v$G35_9913_out0 && v$G36_3925_out0;
assign v$G40_8947_out0 = v$G35_9924_out0 && v$G36_3936_out0;
assign v$G40_8948_out0 = v$G35_9925_out0 && v$G36_3937_out0;
assign v$SEL2_9281_out0 = v$B$MANTISSA_1575_out0[11:0];
assign v$SEL2_9282_out0 = v$B$MANTISSA_1576_out0[11:0];
assign v$A1_9730_out0 = v$SEL4_4936_out0;
assign v$A1_9731_out0 = v$SEL4_4937_out0;
assign v$A1_9733_out0 = v$SEL4_4939_out0;
assign v$A1_9734_out0 = v$SEL4_4940_out0;
assign v$A1_9742_out0 = v$SEL4_4948_out0;
assign v$A1_9743_out0 = v$SEL4_4949_out0;
assign v$A1_9745_out0 = v$SEL4_4951_out0;
assign v$A1_9746_out0 = v$SEL4_4952_out0;
assign v$B_9821_out0 = v$SEL3_6298_out0;
assign v$B_9822_out0 = v$SEL2_12245_out0;
assign v$B_9837_out0 = v$SEL3_6302_out0;
assign v$B_9838_out0 = v$SEL2_12249_out0;
assign v$StatRegAdd1_9943_out0 = v$ADD_1721_out0 == 12'hffd;
assign v$StatRegAdd1_9944_out0 = v$ADD_1722_out0 == 12'hffd;
assign v$A3XNORB3_10073_out0 = v$G8_2440_out0;
assign v$A3XNORB3_10074_out0 = v$G8_2441_out0;
assign v$A3XNORB3_10081_out0 = v$G8_2448_out0;
assign v$A3XNORB3_10085_out0 = v$G8_2452_out0;
assign v$A3XNORB3_10086_out0 = v$G8_2453_out0;
assign v$A3XNORB3_10093_out0 = v$G8_2460_out0;
assign v$TXRegAdd_10869_out0 = v$ADD_1721_out0 == 12'hfff;
assign v$TXRegAdd_10870_out0 = v$ADD_1722_out0 == 12'hfff;
assign v$G11_10907_out0 = v$A2_5565_out0 && v$G12_11547_out0;
assign v$G11_10908_out0 = v$A2_5566_out0 && v$G12_11548_out0;
assign v$G11_10915_out0 = v$A2_5573_out0 && v$G12_11555_out0;
assign v$G11_10919_out0 = v$A2_5577_out0 && v$G12_11559_out0;
assign v$G11_10920_out0 = v$A2_5578_out0 && v$G12_11560_out0;
assign v$G11_10927_out0 = v$A2_5585_out0 && v$G12_11567_out0;
assign v$A1XNORB1_11226_out0 = v$G16_11912_out0;
assign v$A1XNORB1_11227_out0 = v$G16_11913_out0;
assign v$A1XNORB1_11234_out0 = v$G16_11920_out0;
assign v$A1XNORB1_11238_out0 = v$G16_11924_out0;
assign v$A1XNORB1_11239_out0 = v$G16_11925_out0;
assign v$A1XNORB1_11246_out0 = v$G16_11932_out0;
assign v$G39_12168_out0 = v$G36_3932_out0 && v$G37_744_out0;
assign v$G39_12170_out0 = v$G36_3944_out0 && v$G37_746_out0;
assign v$SAME_13064_out0 = v$SAME_13351_out0;
assign v$SAME_13068_out0 = v$SAME_13367_out0;
assign v$VALID_13300_out0 = v$VALID_9883_out0;
assign v$VALID_13301_out0 = v$VALID_9884_out0;
assign v$G7_1165_out0 = v$A4XNORB4_598_out0 && v$G5_4713_out0;
assign v$G7_1167_out0 = v$A4XNORB4_600_out0 && v$G5_4725_out0;
assign v$SEL7_2866_out0 = v$B_9821_out0[3:3];
assign v$SEL7_2867_out0 = v$B_9822_out0[3:3];
assign v$SEL7_2878_out0 = v$B_9837_out0[3:3];
assign v$SEL7_2879_out0 = v$B_9838_out0[3:3];
assign v$G13_3055_out0 = v$A3XNORB3_10073_out0 && v$G11_10907_out0;
assign v$G13_3056_out0 = v$A3XNORB3_10074_out0 && v$G11_10908_out0;
assign v$G13_3063_out0 = v$A3XNORB3_10081_out0 && v$G11_10915_out0;
assign v$G13_3067_out0 = v$A3XNORB3_10085_out0 && v$G11_10919_out0;
assign v$G13_3068_out0 = v$A3XNORB3_10086_out0 && v$G11_10920_out0;
assign v$G13_3075_out0 = v$A3XNORB3_10093_out0 && v$G11_10927_out0;
assign v$A3$COMP$B3_3339_out0 = v$G5_4705_out0;
assign v$A3$COMP$B3_3340_out0 = v$G5_4706_out0;
assign v$A3$COMP$B3_3351_out0 = v$G5_4717_out0;
assign v$A3$COMP$B3_3352_out0 = v$G5_4718_out0;
assign v$MUX1_4668_out0 = v$G4_2747_out0 ? v$_7609_out0 : v$MUX2_7823_out0;
assign v$MUX1_4672_out0 = v$G4_2751_out0 ? v$_7613_out0 : v$MUX2_7827_out0;
assign v$A4$COMP$B4_4998_out0 = v$G2_6950_out0;
assign v$A4$COMP$B4_5000_out0 = v$G2_6952_out0;
assign v$G3_5136_out0 = v$TXRegAdd_10869_out0 && v$WEN_13084_out0;
assign v$G3_5137_out0 = v$TXRegAdd_10870_out0 && v$WEN_13085_out0;
assign v$G7_5269_out0 = v$StatRegAdd1_9943_out0 && v$G8_8973_out0;
assign v$G7_5270_out0 = v$StatRegAdd1_9944_out0 && v$G8_8974_out0;
assign v$A0$COMP$B0_5492_out0 = v$G26_7414_out0;
assign v$A0$COMP$B0_5504_out0 = v$G26_7416_out0;
assign v$I0EN_5551_out0 = v$I0REGISTERWRITE_2048_out0;
assign v$I0EN_5552_out0 = v$I0REGISTERWRITE_2049_out0;
assign v$G5_5904_out0 = v$RXRegAdd_8613_out0 && v$G6_382_out0;
assign v$G5_5905_out0 = v$RXRegAdd_8614_out0 && v$G6_383_out0;
assign v$SEL9_7138_out0 = v$B_9821_out0[1:1];
assign v$SEL9_7139_out0 = v$B_9822_out0[1:1];
assign v$SEL9_7150_out0 = v$B_9837_out0[1:1];
assign v$SEL9_7151_out0 = v$B_9838_out0[1:1];
assign v$G41_7157_out0 = v$G38_4890_out0 && v$G40_8935_out0;
assign v$G41_7158_out0 = v$G38_4891_out0 && v$G40_8936_out0;
assign v$G41_7169_out0 = v$G38_4902_out0 && v$G40_8947_out0;
assign v$G41_7170_out0 = v$G38_4903_out0 && v$G40_8948_out0;
assign v$B_7905_out0 = v$SEL4_589_out0;
assign v$B_7906_out0 = v$SEL2_9281_out0;
assign v$B_7907_out0 = v$SEL4_590_out0;
assign v$B_7908_out0 = v$SEL2_9282_out0;
assign v$SEL10_8258_out0 = v$B_9821_out0[0:0];
assign v$SEL10_8259_out0 = v$B_9822_out0[0:0];
assign v$SEL10_8270_out0 = v$B_9837_out0[0:0];
assign v$SEL10_8271_out0 = v$B_9838_out0[0:0];
assign v$SEL8_8569_out0 = v$B_9821_out0[2:2];
assign v$SEL8_8570_out0 = v$B_9822_out0[2:2];
assign v$SEL8_8581_out0 = v$B_9837_out0[2:2];
assign v$SEL8_8582_out0 = v$B_9838_out0[2:2];
assign v$G28_8639_out0 = v$A1XNORB1_11226_out0 && v$G25_7204_out0;
assign v$G28_8640_out0 = v$A1XNORB1_11227_out0 && v$G25_7205_out0;
assign v$G28_8647_out0 = v$A1XNORB1_11234_out0 && v$G25_7212_out0;
assign v$G28_8651_out0 = v$A1XNORB1_11238_out0 && v$G25_7216_out0;
assign v$G28_8652_out0 = v$A1XNORB1_11239_out0 && v$G25_7217_out0;
assign v$G28_8659_out0 = v$A1XNORB1_11246_out0 && v$G25_7224_out0;
assign v$G22_8902_out0 = v$A2XNORB2_3126_out0 && v$G20_6620_out0;
assign v$G22_8903_out0 = v$A2XNORB2_3127_out0 && v$G20_6621_out0;
assign v$G22_8910_out0 = v$A2XNORB2_3134_out0 && v$G20_6628_out0;
assign v$G22_8914_out0 = v$A2XNORB2_3138_out0 && v$G20_6632_out0;
assign v$G22_8915_out0 = v$A2XNORB2_3139_out0 && v$G20_6633_out0;
assign v$G22_8922_out0 = v$A2XNORB2_3146_out0 && v$G20_6640_out0;
assign v$G40_8943_out0 = v$G35_9920_out0 && v$G39_12168_out0;
assign v$G40_8955_out0 = v$G35_9932_out0 && v$G39_12170_out0;
assign v$COUNTEREN_9016_out0 = v$COUNTEREN_828_out0;
assign v$COUNTEREN_9017_out0 = v$COUNTEREN_829_out0;
assign v$RAMADDR_9169_out0 = v$MUX1_1023_out0;
assign v$ENMODE_9952_out0 = v$MODEEN_3782_out0;
assign v$ENMODE_9953_out0 = v$MODEEN_3783_out0;
assign v$G9_10859_out0 = v$ModeRegAdd_2724_out0 && v$WEN_13084_out0;
assign v$G9_10860_out0 = v$ModeRegAdd_2725_out0 && v$WEN_13085_out0;
assign v$I2EN_10989_out0 = v$I2REGISTERWRITE_7720_out0;
assign v$I2EN_10990_out0 = v$I2REGISTERWRITE_7721_out0;
assign v$G1_11506_out0 = v$StatRegAdd_5285_out0 && v$WEN_13084_out0;
assign v$G1_11507_out0 = v$StatRegAdd_5286_out0 && v$WEN_13085_out0;
assign v$I3EN_12565_out0 = v$I3REGISTERWRITE_521_out0;
assign v$I3EN_12566_out0 = v$I3REGISTERWRITE_522_out0;
assign v$VALID_12693_out0 = v$VALID_13300_out0;
assign v$VALID_12694_out0 = v$VALID_13301_out0;
assign v$I1EN_13089_out0 = v$I1REGISTERWRITE_1698_out0;
assign v$I1EN_13090_out0 = v$I1REGISTERWRITE_1699_out0;
assign v$G32_321_out0 = v$A1$COMP$B1_8127_out0 || v$A0$COMP$B0_5492_out0;
assign v$G32_333_out0 = v$A1$COMP$B1_8139_out0 || v$A0$COMP$B0_5504_out0;
assign v$MUX3_1099_out0 = v$G8_1037_out0 ? v$_8878_out0 : v$MUX1_4668_out0;
assign v$MUX3_1103_out0 = v$G8_1041_out0 ? v$_8882_out0 : v$MUX1_4672_out0;
assign v$A2$COMP$B2_1116_out0 = v$G13_3055_out0;
assign v$A2$COMP$B2_1117_out0 = v$G13_3056_out0;
assign v$A2$COMP$B2_1128_out0 = v$G13_3067_out0;
assign v$A2$COMP$B2_1129_out0 = v$G13_3068_out0;
assign v$B0_2358_out0 = v$SEL10_8258_out0;
assign v$B0_2359_out0 = v$SEL10_8259_out0;
assign v$B0_2370_out0 = v$SEL10_8270_out0;
assign v$B0_2371_out0 = v$SEL10_8271_out0;
assign v$VALID_2425_out0 = v$VALID_12693_out0;
assign v$VALID_2426_out0 = v$VALID_12694_out0;
assign v$ModeWrite_3091_out0 = v$G9_10859_out0;
assign v$ModeWrite_3092_out0 = v$G9_10860_out0;
assign v$G27_3186_out0 = v$A2XNORB2_3126_out0 && v$G28_8639_out0;
assign v$G27_3187_out0 = v$A2XNORB2_3127_out0 && v$G28_8640_out0;
assign v$G27_3194_out0 = v$A2XNORB2_3134_out0 && v$G28_8647_out0;
assign v$G27_3198_out0 = v$A2XNORB2_3138_out0 && v$G28_8651_out0;
assign v$G27_3199_out0 = v$A2XNORB2_3139_out0 && v$G28_8652_out0;
assign v$G27_3206_out0 = v$A2XNORB2_3146_out0 && v$G28_8659_out0;
assign v$A3$COMP$B3_3347_out0 = v$G7_1165_out0;
assign v$A3$COMP$B3_3359_out0 = v$G7_1167_out0;
assign v$G18_3367_out0 = v$A3XNORB3_10073_out0 && v$G22_8902_out0;
assign v$G18_3368_out0 = v$A3XNORB3_10074_out0 && v$G22_8903_out0;
assign v$G18_3375_out0 = v$A3XNORB3_10081_out0 && v$G22_8910_out0;
assign v$G18_3379_out0 = v$A3XNORB3_10085_out0 && v$G22_8914_out0;
assign v$G18_3380_out0 = v$A3XNORB3_10086_out0 && v$G22_8915_out0;
assign v$G18_3387_out0 = v$A3XNORB3_10093_out0 && v$G22_8922_out0;
assign v$THRESHOLD$WRITE_4845_out0 = v$COUNTEREN_9016_out0;
assign v$THRESHOLD$WRITE_4846_out0 = v$COUNTEREN_9017_out0;
assign v$ENMODE_5281_out0 = v$ENMODE_9952_out0;
assign v$ENMODE_5282_out0 = v$ENMODE_9953_out0;
assign v$RAMADDR_6006_out0 = v$RAMADDR_9169_out0;
assign v$SEL4_6540_out0 = v$B_7905_out0[11:8];
assign v$SEL4_6541_out0 = v$B_7906_out0[11:8];
assign v$SEL4_6542_out0 = v$B_7907_out0[11:8];
assign v$SEL4_6543_out0 = v$B_7908_out0[11:8];
assign v$STRead_6652_out0 = v$G7_5269_out0;
assign v$STRead_6653_out0 = v$G7_5270_out0;
assign v$STClr_6793_out0 = v$G1_11506_out0;
assign v$STClr_6794_out0 = v$G1_11507_out0;
assign v$G41_7165_out0 = v$G38_4898_out0 && v$G40_8943_out0;
assign v$G41_7177_out0 = v$G38_4910_out0 && v$G40_8955_out0;
assign v$G14_8285_out0 = v$A4XNORB4_598_out0 && v$G13_3063_out0;
assign v$G14_8287_out0 = v$A4XNORB4_600_out0 && v$G13_3075_out0;
assign v$B1_9627_out0 = v$SEL9_7138_out0;
assign v$B1_9628_out0 = v$SEL9_7139_out0;
assign v$B1_9639_out0 = v$SEL9_7150_out0;
assign v$B1_9640_out0 = v$SEL9_7151_out0;
assign v$RXRead_11475_out0 = v$G5_5904_out0;
assign v$RXRead_11476_out0 = v$G5_5905_out0;
assign v$B2_11706_out0 = v$SEL8_8569_out0;
assign v$B2_11707_out0 = v$SEL8_8570_out0;
assign v$B2_11718_out0 = v$SEL8_8581_out0;
assign v$B2_11719_out0 = v$SEL8_8582_out0;
assign v$TXWrite_12290_out0 = v$G3_5136_out0;
assign v$TXWrite_12291_out0 = v$G3_5137_out0;
assign v$SEL2_12312_out0 = v$B_7905_out0[7:0];
assign v$SEL2_12313_out0 = v$B_7906_out0[7:0];
assign v$SEL2_12314_out0 = v$B_7907_out0[7:0];
assign v$SEL2_12315_out0 = v$B_7908_out0[7:0];
assign v$B3_12648_out0 = v$SEL7_2866_out0;
assign v$B3_12649_out0 = v$SEL7_2867_out0;
assign v$B3_12660_out0 = v$SEL7_2878_out0;
assign v$B3_12661_out0 = v$SEL7_2879_out0;
assign v$SAME_13353_out0 = v$G41_7157_out0;
assign v$SAME_13354_out0 = v$G41_7158_out0;
assign v$SAME_13369_out0 = v$G41_7169_out0;
assign v$SAME_13370_out0 = v$G41_7170_out0;
assign v$R_719_out0 = v$VALID_2425_out0;
assign v$R_720_out0 = v$VALID_2426_out0;
assign v$STATUSREAD_835_out0 = v$STRead_6652_out0;
assign v$STATUSREAD_836_out0 = v$STRead_6653_out0;
assign v$A2$COMP$B2_1124_out0 = v$G14_8285_out0;
assign v$A2$COMP$B2_1136_out0 = v$G14_8287_out0;
assign v$OUT_1900_out0 = v$MUX3_1099_out0;
assign v$OUT_1904_out0 = v$MUX3_1103_out0;
assign v$G21_2234_out0 = ! v$B1_9627_out0;
assign v$G21_2235_out0 = ! v$B1_9628_out0;
assign v$G21_2246_out0 = ! v$B1_9639_out0;
assign v$G21_2247_out0 = ! v$B1_9640_out0;
assign v$G8_2449_out0 = !((v$A3_7028_out0 && !v$B3_12648_out0) || (!v$A3_7028_out0) && v$B3_12648_out0);
assign v$G8_2450_out0 = !((v$A3_7029_out0 && !v$B3_12649_out0) || (!v$A3_7029_out0) && v$B3_12649_out0);
assign v$G8_2461_out0 = !((v$A3_7040_out0 && !v$B3_12660_out0) || (!v$A3_7040_out0) && v$B3_12660_out0);
assign v$G8_2462_out0 = !((v$A3_7041_out0 && !v$B3_12661_out0) || (!v$A3_7041_out0) && v$B3_12661_out0);
assign v$G36_3933_out0 = !((v$B3_12648_out0 && !v$A3_7028_out0) || (!v$B3_12648_out0) && v$A3_7028_out0);
assign v$G36_3934_out0 = !((v$B3_12649_out0 && !v$A3_7029_out0) || (!v$B3_12649_out0) && v$A3_7029_out0);
assign v$G36_3945_out0 = !((v$B3_12660_out0 && !v$A3_7040_out0) || (!v$B3_12660_out0) && v$A3_7040_out0);
assign v$G36_3946_out0 = !((v$B3_12661_out0 && !v$A3_7041_out0) || (!v$B3_12661_out0) && v$A3_7041_out0);
assign v$STATUSCLR_3955_out0 = v$STClr_6793_out0;
assign v$STATUSCLR_3956_out0 = v$STClr_6794_out0;
assign v$G6_4564_out0 = ! v$B3_12648_out0;
assign v$G6_4565_out0 = ! v$B3_12649_out0;
assign v$G6_4576_out0 = ! v$B3_12660_out0;
assign v$G6_4577_out0 = ! v$B3_12661_out0;
assign v$G17_5680_out0 = !((v$A0_915_out0 && !v$B0_2358_out0) || (!v$A0_915_out0) && v$B0_2358_out0);
assign v$G17_5681_out0 = !((v$A0_916_out0 && !v$B0_2359_out0) || (!v$A0_916_out0) && v$B0_2359_out0);
assign v$G17_5692_out0 = !((v$A0_927_out0 && !v$B0_2370_out0) || (!v$A0_927_out0) && v$B0_2370_out0);
assign v$G17_5693_out0 = !((v$A0_928_out0 && !v$B0_2371_out0) || (!v$A0_928_out0) && v$B0_2371_out0);
assign v$LOWER$SAME_6757_out0 = v$SAME_13354_out0;
assign v$LOWER$SAME_6761_out0 = v$SAME_13370_out0;
assign v$G19_6818_out0 = v$A4XNORB4_598_out0 && v$G18_3375_out0;
assign v$G19_6820_out0 = v$A4XNORB4_600_out0 && v$G18_3387_out0;
assign v$TXWRITE_7348_out0 = v$TXWrite_12290_out0;
assign v$TXWRITE_7349_out0 = v$TXWrite_12291_out0;
assign v$G23_7958_out0 = ! v$B0_2358_out0;
assign v$G23_7959_out0 = ! v$B0_2359_out0;
assign v$G23_7970_out0 = ! v$B0_2370_out0;
assign v$G23_7971_out0 = ! v$B0_2371_out0;
assign v$A1$COMP$B1_8128_out0 = v$G18_3367_out0;
assign v$A1$COMP$B1_8129_out0 = v$G18_3368_out0;
assign v$A1$COMP$B1_8140_out0 = v$G18_3379_out0;
assign v$A1$COMP$B1_8141_out0 = v$G18_3380_out0;
assign v$G33_8732_out0 = !((v$A0_915_out0 && !v$B0_2358_out0) || (!v$A0_915_out0) && v$B0_2358_out0);
assign v$G33_8733_out0 = !((v$A0_916_out0 && !v$B0_2359_out0) || (!v$A0_916_out0) && v$B0_2359_out0);
assign v$G33_8744_out0 = !((v$A0_927_out0 && !v$B0_2370_out0) || (!v$A0_927_out0) && v$B0_2370_out0);
assign v$G33_8745_out0 = !((v$A0_928_out0 && !v$B0_2371_out0) || (!v$A0_928_out0) && v$B0_2371_out0);
assign v$G5_9119_out0 = v$EQUAL_11046_out0 || v$THRESHOLD$WRITE_4845_out0;
assign v$G5_9120_out0 = v$EQUAL_11047_out0 || v$THRESHOLD$WRITE_4846_out0;
assign v$G15_9205_out0 = !((v$A2_5574_out0 && !v$B2_11706_out0) || (!v$A2_5574_out0) && v$B2_11706_out0);
assign v$G15_9206_out0 = !((v$A2_5575_out0 && !v$B2_11707_out0) || (!v$A2_5575_out0) && v$B2_11707_out0);
assign v$G15_9217_out0 = !((v$A2_5586_out0 && !v$B2_11718_out0) || (!v$A2_5586_out0) && v$B2_11718_out0);
assign v$G15_9218_out0 = !((v$A2_5587_out0 && !v$B2_11719_out0) || (!v$A2_5587_out0) && v$B2_11719_out0);
assign v$B_9811_out0 = v$SEL4_6540_out0;
assign v$B_9812_out0 = v$SEL2_12312_out0;
assign v$B_9815_out0 = v$SEL4_6541_out0;
assign v$B_9816_out0 = v$SEL2_12313_out0;
assign v$B_9827_out0 = v$SEL4_6542_out0;
assign v$B_9828_out0 = v$SEL2_12314_out0;
assign v$B_9831_out0 = v$SEL4_6543_out0;
assign v$B_9832_out0 = v$SEL2_12315_out0;
assign v$G35_9921_out0 = !((v$A2_5574_out0 && !v$B2_11706_out0) || (!v$A2_5574_out0) && v$B2_11706_out0);
assign v$G35_9922_out0 = !((v$A2_5575_out0 && !v$B2_11707_out0) || (!v$A2_5575_out0) && v$B2_11707_out0);
assign v$G35_9933_out0 = !((v$A2_5586_out0 && !v$B2_11718_out0) || (!v$A2_5586_out0) && v$B2_11718_out0);
assign v$G35_9934_out0 = !((v$A2_5587_out0 && !v$B2_11719_out0) || (!v$A2_5587_out0) && v$B2_11719_out0);
assign v$MODEWRITE_10070_out0 = v$ModeWrite_3091_out0;
assign v$MODEWRITE_10071_out0 = v$ModeWrite_3092_out0;
assign v$HIGHER$SAME_10331_out0 = v$SAME_13353_out0;
assign v$HIGHER$SAME_10335_out0 = v$SAME_13369_out0;
assign v$G31_10787_out0 = v$A2$COMP$B2_1115_out0 || v$G32_321_out0;
assign v$G31_10799_out0 = v$A2$COMP$B2_1127_out0 || v$G32_333_out0;
assign v$G24_10948_out0 = v$A3XNORB3_10073_out0 && v$G27_3186_out0;
assign v$G24_10949_out0 = v$A3XNORB3_10074_out0 && v$G27_3187_out0;
assign v$G24_10956_out0 = v$A3XNORB3_10081_out0 && v$G27_3194_out0;
assign v$G24_10960_out0 = v$A3XNORB3_10085_out0 && v$G27_3198_out0;
assign v$G24_10961_out0 = v$A3XNORB3_10086_out0 && v$G27_3199_out0;
assign v$G24_10968_out0 = v$A3XNORB3_10093_out0 && v$G27_3206_out0;
assign v$RXREAD_11072_out0 = v$RXRead_11475_out0;
assign v$RXREAD_11073_out0 = v$RXRead_11476_out0;
assign v$EN_11112_out0 = v$ENMODE_5281_out0;
assign v$EN_11113_out0 = v$ENMODE_5282_out0;
assign v$G12_11556_out0 = ! v$B2_11706_out0;
assign v$G12_11557_out0 = ! v$B2_11707_out0;
assign v$G12_11568_out0 = ! v$B2_11718_out0;
assign v$G12_11569_out0 = ! v$B2_11719_out0;
assign v$G16_11921_out0 = !((v$A1_9736_out0 && !v$B1_9627_out0) || (!v$A1_9736_out0) && v$B1_9627_out0);
assign v$G16_11922_out0 = !((v$A1_9737_out0 && !v$B1_9628_out0) || (!v$A1_9737_out0) && v$B1_9628_out0);
assign v$G16_11933_out0 = !((v$A1_9748_out0 && !v$B1_9639_out0) || (!v$A1_9748_out0) && v$B1_9639_out0);
assign v$G16_11934_out0 = !((v$A1_9749_out0 && !v$B1_9640_out0) || (!v$A1_9749_out0) && v$B1_9640_out0);
assign v$G34_12131_out0 = !((v$A1_9736_out0 && !v$B1_9627_out0) || (!v$A1_9736_out0) && v$B1_9627_out0);
assign v$G34_12132_out0 = !((v$A1_9737_out0 && !v$B1_9628_out0) || (!v$A1_9737_out0) && v$B1_9628_out0);
assign v$G34_12143_out0 = !((v$A1_9748_out0 && !v$B1_9639_out0) || (!v$A1_9748_out0) && v$B1_9639_out0);
assign v$G34_12144_out0 = !((v$A1_9749_out0 && !v$B1_9640_out0) || (!v$A1_9749_out0) && v$B1_9640_out0);
assign v$RAMADDR_13293_out0 = v$RAMADDR_6006_out0;
assign v$SAME_13363_out0 = v$G41_7165_out0;
assign v$SAME_13379_out0 = v$G41_7177_out0;
assign v$A0XNORB0_679_out0 = v$G17_5680_out0;
assign v$A0XNORB0_680_out0 = v$G17_5681_out0;
assign v$A0XNORB0_691_out0 = v$G17_5692_out0;
assign v$A0XNORB0_692_out0 = v$G17_5693_out0;
assign v$R_789_out0 = v$R_719_out0;
assign v$R_790_out0 = v$R_720_out0;
assign v$G30_948_out0 = v$A3$COMP$B3_3338_out0 || v$G31_10787_out0;
assign v$G30_960_out0 = v$A3$COMP$B3_3350_out0 || v$G31_10799_out0;
assign v$WREN_1443_out0 = v$TXWRITE_7348_out0;
assign v$WREN_1444_out0 = v$TXWRITE_7349_out0;
assign v$SEL7_2859_out0 = v$B_9811_out0[3:3];
assign v$SEL7_2862_out0 = v$B_9815_out0[3:3];
assign v$SEL7_2871_out0 = v$B_9827_out0[3:3];
assign v$SEL7_2874_out0 = v$B_9831_out0[3:3];
assign v$G1_2894_out0 = v$STATUSREAD_835_out0 || v$RXREAD_11072_out0;
assign v$G1_2895_out0 = v$STATUSREAD_836_out0 || v$RXREAD_11073_out0;
assign v$IN_3018_out0 = v$OUT_1900_out0;
assign v$IN_3022_out0 = v$OUT_1904_out0;
assign v$A2XNORB2_3135_out0 = v$G15_9205_out0;
assign v$A2XNORB2_3136_out0 = v$G15_9206_out0;
assign v$A2XNORB2_3147_out0 = v$G15_9217_out0;
assign v$A2XNORB2_3148_out0 = v$G15_9218_out0;
assign v$RXreset_3961_out0 = v$RXREAD_11072_out0;
assign v$RXreset_3962_out0 = v$RXREAD_11073_out0;
assign v$G5_4714_out0 = v$A3_7028_out0 && v$G6_4564_out0;
assign v$G5_4715_out0 = v$A3_7029_out0 && v$G6_4565_out0;
assign v$G5_4726_out0 = v$A3_7040_out0 && v$G6_4576_out0;
assign v$G5_4727_out0 = v$A3_7041_out0 && v$G6_4577_out0;
assign v$_4875_out0 = v$RAMADDR_13293_out0[3:0];
assign v$_4875_out1 = v$RAMADDR_13293_out0[11:8];
assign v$G38_4899_out0 = v$G33_8732_out0 && v$G34_12131_out0;
assign v$G38_4900_out0 = v$G33_8733_out0 && v$G34_12132_out0;
assign v$G38_4911_out0 = v$G33_8744_out0 && v$G34_12143_out0;
assign v$G38_4912_out0 = v$G33_8745_out0 && v$G34_12144_out0;
assign v$A0$COMP$B0_5493_out0 = v$G24_10948_out0;
assign v$A0$COMP$B0_5494_out0 = v$G24_10949_out0;
assign v$A0$COMP$B0_5505_out0 = v$G24_10960_out0;
assign v$A0$COMP$B0_5506_out0 = v$G24_10961_out0;
assign v$SEL3_6296_out0 = v$B_9812_out0[7:4];
assign v$SEL3_6297_out0 = v$B_9816_out0[7:4];
assign v$SEL3_6300_out0 = v$B_9828_out0[7:4];
assign v$SEL3_6301_out0 = v$B_9832_out0[7:4];
assign v$G1_6387_out0 = v$LOWER$SAME_6757_out0 && v$HIGHER$SAME_10331_out0;
assign v$G1_6391_out0 = v$LOWER$SAME_6761_out0 && v$HIGHER$SAME_10335_out0;
assign v$G20_6629_out0 = v$A1_9736_out0 && v$G21_2234_out0;
assign v$G20_6630_out0 = v$A1_9737_out0 && v$G21_2235_out0;
assign v$G20_6641_out0 = v$A1_9748_out0 && v$G21_2246_out0;
assign v$G20_6642_out0 = v$A1_9749_out0 && v$G21_2247_out0;
assign v$SEL9_7131_out0 = v$B_9811_out0[1:1];
assign v$SEL9_7134_out0 = v$B_9815_out0[1:1];
assign v$SEL9_7143_out0 = v$B_9827_out0[1:1];
assign v$SEL9_7146_out0 = v$B_9831_out0[1:1];
assign v$G25_7213_out0 = v$A0_915_out0 && v$G23_7958_out0;
assign v$G25_7214_out0 = v$A0_916_out0 && v$G23_7959_out0;
assign v$G25_7225_out0 = v$A0_927_out0 && v$G23_7970_out0;
assign v$G25_7226_out0 = v$A0_928_out0 && v$G23_7971_out0;
assign v$G26_7415_out0 = v$A4XNORB4_598_out0 && v$G24_10956_out0;
assign v$G26_7417_out0 = v$A4XNORB4_600_out0 && v$G24_10968_out0;
assign v$A1$COMP$B1_8136_out0 = v$G19_6818_out0;
assign v$A1$COMP$B1_8148_out0 = v$G19_6820_out0;
assign v$SEL10_8251_out0 = v$B_9811_out0[0:0];
assign v$SEL10_8254_out0 = v$B_9815_out0[0:0];
assign v$SEL10_8263_out0 = v$B_9827_out0[0:0];
assign v$SEL10_8266_out0 = v$B_9831_out0[0:0];
assign v$Clear_8404_out0 = v$STATUSCLR_3955_out0;
assign v$Clear_8405_out0 = v$STATUSCLR_3956_out0;
assign v$SEL8_8562_out0 = v$B_9811_out0[2:2];
assign v$SEL8_8565_out0 = v$B_9815_out0[2:2];
assign v$SEL8_8574_out0 = v$B_9827_out0[2:2];
assign v$SEL8_8577_out0 = v$B_9831_out0[2:2];
assign v$G40_8944_out0 = v$G35_9921_out0 && v$G36_3933_out0;
assign v$G40_8945_out0 = v$G35_9922_out0 && v$G36_3934_out0;
assign v$G40_8956_out0 = v$G35_9933_out0 && v$G36_3945_out0;
assign v$G40_8957_out0 = v$G35_9934_out0 && v$G36_3946_out0;
assign v$TXSet_9724_out0 = v$TXWRITE_7348_out0;
assign v$TXSet_9725_out0 = v$TXWRITE_7349_out0;
assign v$A3XNORB3_10082_out0 = v$G8_2449_out0;
assign v$A3XNORB3_10083_out0 = v$G8_2450_out0;
assign v$A3XNORB3_10094_out0 = v$G8_2461_out0;
assign v$A3XNORB3_10095_out0 = v$G8_2462_out0;
assign v$G11_10916_out0 = v$A2_5574_out0 && v$G12_11556_out0;
assign v$G11_10917_out0 = v$A2_5575_out0 && v$G12_11557_out0;
assign v$G11_10928_out0 = v$A2_5586_out0 && v$G12_11568_out0;
assign v$G11_10929_out0 = v$A2_5587_out0 && v$G12_11569_out0;
assign v$A1XNORB1_11235_out0 = v$G16_11921_out0;
assign v$A1XNORB1_11236_out0 = v$G16_11922_out0;
assign v$A1XNORB1_11247_out0 = v$G16_11933_out0;
assign v$A1XNORB1_11248_out0 = v$G16_11934_out0;
assign v$SEL2_12243_out0 = v$B_9812_out0[3:0];
assign v$SEL2_12244_out0 = v$B_9816_out0[3:0];
assign v$SEL2_12247_out0 = v$B_9828_out0[3:0];
assign v$SEL2_12248_out0 = v$B_9832_out0[3:0];
assign v$MUX1_13028_out0 = v$G5_9119_out0 ? v$C3_7978_out0 : v$A1_9247_out0;
assign v$MUX1_13029_out0 = v$G5_9120_out0 ? v$C3_7979_out0 : v$A1_9248_out0;
assign v$SAME_13066_out0 = v$SAME_13363_out0;
assign v$SAME_13070_out0 = v$SAME_13379_out0;
assign v$G32_322_out0 = v$A1$COMP$B1_8128_out0 || v$A0$COMP$B0_5493_out0;
assign v$G32_323_out0 = v$A1$COMP$B1_8129_out0 || v$A0$COMP$B0_5494_out0;
assign v$G32_334_out0 = v$A1$COMP$B1_8140_out0 || v$A0$COMP$B0_5505_out0;
assign v$G32_335_out0 = v$A1$COMP$B1_8141_out0 || v$A0$COMP$B0_5506_out0;
assign v$SEL8_1110_out0 = v$_4875_out1[7:7];
assign v$SEL3_1872_out0 = v$_4875_out1[2:2];
assign v$B0_2351_out0 = v$SEL10_8251_out0;
assign v$B0_2354_out0 = v$SEL10_8254_out0;
assign v$B0_2363_out0 = v$SEL10_8263_out0;
assign v$B0_2366_out0 = v$SEL10_8266_out0;
assign v$G13_3064_out0 = v$A3XNORB3_10082_out0 && v$G11_10916_out0;
assign v$G13_3065_out0 = v$A3XNORB3_10083_out0 && v$G11_10917_out0;
assign v$G13_3076_out0 = v$A3XNORB3_10094_out0 && v$G11_10928_out0;
assign v$G13_3077_out0 = v$A3XNORB3_10095_out0 && v$G11_10929_out0;
assign v$A3$COMP$B3_3348_out0 = v$G5_4714_out0;
assign v$A3$COMP$B3_3349_out0 = v$G5_4715_out0;
assign v$A3$COMP$B3_3360_out0 = v$G5_4726_out0;
assign v$A3$COMP$B3_3361_out0 = v$G5_4727_out0;
assign v$SEL1_4765_out0 = v$_4875_out1[0:0];
assign v$A0$COMP$B0_5501_out0 = v$G26_7415_out0;
assign v$A0$COMP$B0_5513_out0 = v$G26_7417_out0;
assign v$IN_6534_out0 = v$IN_3018_out0;
assign v$IN_6538_out0 = v$IN_3022_out0;
assign v$G29_6859_out0 = v$A4$COMP$B4_4997_out0 || v$G30_948_out0;
assign v$G29_6861_out0 = v$A4$COMP$B4_4999_out0 || v$G30_960_out0;
assign v$G41_7166_out0 = v$G38_4899_out0 && v$G40_8944_out0;
assign v$G41_7167_out0 = v$G38_4900_out0 && v$G40_8945_out0;
assign v$G41_7178_out0 = v$G38_4911_out0 && v$G40_8956_out0;
assign v$G41_7179_out0 = v$G38_4912_out0 && v$G40_8957_out0;
assign v$WREN_7251_out0 = v$WREN_1443_out0;
assign v$WREN_7252_out0 = v$WREN_1444_out0;
assign v$SEL5_7466_out0 = v$_4875_out1[4:4];
assign v$TXSet_8294_out0 = v$TXSet_9724_out0;
assign v$TXSet_8295_out0 = v$TXSet_9725_out0;
assign v$G28_8648_out0 = v$A1XNORB1_11235_out0 && v$G25_7213_out0;
assign v$G28_8649_out0 = v$A1XNORB1_11236_out0 && v$G25_7214_out0;
assign v$G28_8660_out0 = v$A1XNORB1_11247_out0 && v$G25_7225_out0;
assign v$G28_8661_out0 = v$A1XNORB1_11248_out0 && v$G25_7226_out0;
assign v$G22_8911_out0 = v$A2XNORB2_3135_out0 && v$G20_6629_out0;
assign v$G22_8912_out0 = v$A2XNORB2_3136_out0 && v$G20_6630_out0;
assign v$G22_8923_out0 = v$A2XNORB2_3147_out0 && v$G20_6641_out0;
assign v$G22_8924_out0 = v$A2XNORB2_3148_out0 && v$G20_6642_out0;
assign v$B1_9620_out0 = v$SEL9_7131_out0;
assign v$B1_9623_out0 = v$SEL9_7134_out0;
assign v$B1_9632_out0 = v$SEL9_7143_out0;
assign v$B1_9635_out0 = v$SEL9_7146_out0;
assign v$SEL6_9641_out0 = v$_4875_out1[5:5];
assign v$B_9813_out0 = v$SEL3_6296_out0;
assign v$B_9814_out0 = v$SEL2_12243_out0;
assign v$B_9817_out0 = v$SEL3_6297_out0;
assign v$B_9818_out0 = v$SEL2_12244_out0;
assign v$B_9829_out0 = v$SEL3_6300_out0;
assign v$B_9830_out0 = v$SEL2_12247_out0;
assign v$B_9833_out0 = v$SEL3_6301_out0;
assign v$B_9834_out0 = v$SEL2_12248_out0;
assign v$Clear_10010_out0 = v$Clear_8404_out0;
assign v$Clear_10011_out0 = v$Clear_8405_out0;
assign v$USELESS_10774_out0 = v$_4875_out0;
assign v$SEL2_11054_out0 = v$_4875_out1[1:1];
assign v$SEL4_11518_out0 = v$_4875_out1[3:3];
assign v$B2_11699_out0 = v$SEL8_8562_out0;
assign v$B2_11702_out0 = v$SEL8_8565_out0;
assign v$B2_11711_out0 = v$SEL8_8574_out0;
assign v$B2_11714_out0 = v$SEL8_8577_out0;
assign v$SEL7_12068_out0 = v$_4875_out1[6:6];
assign v$G3_12513_out0 = ! v$R_789_out0;
assign v$G3_12514_out0 = ! v$R_790_out0;
assign v$B3_12641_out0 = v$SEL7_2859_out0;
assign v$B3_12644_out0 = v$SEL7_2862_out0;
assign v$B3_12653_out0 = v$SEL7_2871_out0;
assign v$B3_12656_out0 = v$SEL7_2874_out0;
assign v$G18_12843_out0 = v$WREN_1443_out0 || v$G19_5745_out0;
assign v$G18_12844_out0 = v$WREN_1444_out0 || v$G19_5746_out0;
assign v$R_13039_out0 = v$RXreset_3961_out0;
assign v$R_13050_out0 = v$RXreset_3962_out0;
assign v$SAME_13352_out0 = v$G1_6387_out0;
assign v$SAME_13368_out0 = v$G1_6391_out0;
assign v$G32_330_out0 = v$A1$COMP$B1_8136_out0 || v$A0$COMP$B0_5501_out0;
assign v$G32_342_out0 = v$A1$COMP$B1_8148_out0 || v$A0$COMP$B0_5513_out0;
assign v$_765_out0 = v$IN_6534_out0[15:15];
assign v$_766_out0 = v$IN_6538_out0[15:15];
assign v$A2$COMP$B2_1125_out0 = v$G13_3064_out0;
assign v$A2$COMP$B2_1126_out0 = v$G13_3065_out0;
assign v$A2$COMP$B2_1137_out0 = v$G13_3076_out0;
assign v$A2$COMP$B2_1138_out0 = v$G13_3077_out0;
assign v$G21_2227_out0 = ! v$B1_9620_out0;
assign v$G21_2230_out0 = ! v$B1_9623_out0;
assign v$G21_2239_out0 = ! v$B1_9632_out0;
assign v$G21_2242_out0 = ! v$B1_9635_out0;
assign v$G8_2442_out0 = !((v$A3_7021_out0 && !v$B3_12641_out0) || (!v$A3_7021_out0) && v$B3_12641_out0);
assign v$G8_2445_out0 = !((v$A3_7024_out0 && !v$B3_12644_out0) || (!v$A3_7024_out0) && v$B3_12644_out0);
assign v$G8_2454_out0 = !((v$A3_7033_out0 && !v$B3_12653_out0) || (!v$A3_7033_out0) && v$B3_12653_out0);
assign v$G8_2457_out0 = !((v$A3_7036_out0 && !v$B3_12656_out0) || (!v$A3_7036_out0) && v$B3_12656_out0);
assign v$OUT_2622_out0 = v$G29_6859_out0;
assign v$OUT_2638_out0 = v$G29_6861_out0;
assign v$SEL7_2860_out0 = v$B_9813_out0[3:3];
assign v$SEL7_2861_out0 = v$B_9814_out0[3:3];
assign v$SEL7_2863_out0 = v$B_9817_out0[3:3];
assign v$SEL7_2864_out0 = v$B_9818_out0[3:3];
assign v$SEL7_2872_out0 = v$B_9829_out0[3:3];
assign v$SEL7_2873_out0 = v$B_9830_out0[3:3];
assign v$SEL7_2875_out0 = v$B_9833_out0[3:3];
assign v$SEL7_2876_out0 = v$B_9834_out0[3:3];
assign v$G27_3195_out0 = v$A2XNORB2_3135_out0 && v$G28_8648_out0;
assign v$G27_3196_out0 = v$A2XNORB2_3136_out0 && v$G28_8649_out0;
assign v$G27_3207_out0 = v$A2XNORB2_3147_out0 && v$G28_8660_out0;
assign v$G27_3208_out0 = v$A2XNORB2_3148_out0 && v$G28_8661_out0;
assign v$_3211_out0 = v$IN_6534_out0[11:0];
assign v$_3215_out0 = v$IN_6538_out0[11:0];
assign v$G18_3376_out0 = v$A3XNORB3_10082_out0 && v$G22_8911_out0;
assign v$G18_3377_out0 = v$A3XNORB3_10083_out0 && v$G22_8912_out0;
assign v$G18_3388_out0 = v$A3XNORB3_10094_out0 && v$G22_8923_out0;
assign v$G18_3389_out0 = v$A3XNORB3_10095_out0 && v$G22_8924_out0;
assign v$G3_3394_out0 = v$SEL5_7466_out0 && v$SEL6_9641_out0;
assign v$G36_3926_out0 = !((v$B3_12641_out0 && !v$A3_7021_out0) || (!v$B3_12641_out0) && v$A3_7021_out0);
assign v$G36_3929_out0 = !((v$B3_12644_out0 && !v$A3_7024_out0) || (!v$B3_12644_out0) && v$A3_7024_out0);
assign v$G36_3938_out0 = !((v$B3_12653_out0 && !v$A3_7033_out0) || (!v$B3_12653_out0) && v$A3_7033_out0);
assign v$G36_3941_out0 = !((v$B3_12656_out0 && !v$A3_7036_out0) || (!v$B3_12656_out0) && v$A3_7036_out0);
assign v$G4_4429_out0 = v$SEL7_12068_out0 && v$SEL8_1110_out0;
assign v$G6_4557_out0 = ! v$B3_12641_out0;
assign v$G6_4560_out0 = ! v$B3_12644_out0;
assign v$G6_4569_out0 = ! v$B3_12653_out0;
assign v$G6_4572_out0 = ! v$B3_12656_out0;
assign v$_4977_out0 = v$IN_6534_out0[3:0];
assign v$_4978_out0 = v$IN_6538_out0[3:0];
assign v$ShiftEN_5265_out0 = v$G18_12843_out0;
assign v$ShiftEN_5266_out0 = v$G18_12844_out0;
assign v$G17_5673_out0 = !((v$A0_908_out0 && !v$B0_2351_out0) || (!v$A0_908_out0) && v$B0_2351_out0);
assign v$G17_5676_out0 = !((v$A0_911_out0 && !v$B0_2354_out0) || (!v$A0_911_out0) && v$B0_2354_out0);
assign v$G17_5685_out0 = !((v$A0_920_out0 && !v$B0_2363_out0) || (!v$A0_920_out0) && v$B0_2363_out0);
assign v$G17_5688_out0 = !((v$A0_923_out0 && !v$B0_2366_out0) || (!v$A0_923_out0) && v$B0_2366_out0);
assign v$G9_5922_out0 = v$TXSet_8294_out0 && v$TXLast_7426_out0;
assign v$G9_5923_out0 = v$TXSet_8295_out0 && v$TXLast_7427_out0;
assign v$G17_6145_out0 = ! v$WREN_7251_out0;
assign v$G17_6146_out0 = ! v$WREN_7252_out0;
assign v$SEL9_7132_out0 = v$B_9813_out0[1:1];
assign v$SEL9_7133_out0 = v$B_9814_out0[1:1];
assign v$SEL9_7135_out0 = v$B_9817_out0[1:1];
assign v$SEL9_7136_out0 = v$B_9818_out0[1:1];
assign v$SEL9_7144_out0 = v$B_9829_out0[1:1];
assign v$SEL9_7145_out0 = v$B_9830_out0[1:1];
assign v$SEL9_7147_out0 = v$B_9833_out0[1:1];
assign v$SEL9_7148_out0 = v$B_9834_out0[1:1];
assign v$G2_7517_out0 = v$SEL3_1872_out0 && v$SEL4_11518_out0;
assign v$G23_7951_out0 = ! v$B0_2351_out0;
assign v$G23_7954_out0 = ! v$B0_2354_out0;
assign v$G23_7963_out0 = ! v$B0_2363_out0;
assign v$G23_7966_out0 = ! v$B0_2366_out0;
assign v$SEL10_8252_out0 = v$B_9813_out0[0:0];
assign v$SEL10_8253_out0 = v$B_9814_out0[0:0];
assign v$SEL10_8255_out0 = v$B_9817_out0[0:0];
assign v$SEL10_8256_out0 = v$B_9818_out0[0:0];
assign v$SEL10_8264_out0 = v$B_9829_out0[0:0];
assign v$SEL10_8265_out0 = v$B_9830_out0[0:0];
assign v$SEL10_8267_out0 = v$B_9833_out0[0:0];
assign v$SEL10_8268_out0 = v$B_9834_out0[0:0];
assign v$SEL8_8563_out0 = v$B_9813_out0[2:2];
assign v$SEL8_8564_out0 = v$B_9814_out0[2:2];
assign v$SEL8_8566_out0 = v$B_9817_out0[2:2];
assign v$SEL8_8567_out0 = v$B_9818_out0[2:2];
assign v$SEL8_8575_out0 = v$B_9829_out0[2:2];
assign v$SEL8_8576_out0 = v$B_9830_out0[2:2];
assign v$SEL8_8578_out0 = v$B_9833_out0[2:2];
assign v$SEL8_8579_out0 = v$B_9834_out0[2:2];
assign v$G1_8621_out0 = v$STATE_11196_out0 && v$G3_12513_out0;
assign v$G1_8622_out0 = v$STATE_11197_out0 && v$G3_12514_out0;
assign v$G33_8725_out0 = !((v$A0_908_out0 && !v$B0_2351_out0) || (!v$A0_908_out0) && v$B0_2351_out0);
assign v$G33_8728_out0 = !((v$A0_911_out0 && !v$B0_2354_out0) || (!v$A0_911_out0) && v$B0_2354_out0);
assign v$G33_8737_out0 = !((v$A0_920_out0 && !v$B0_2363_out0) || (!v$A0_920_out0) && v$B0_2363_out0);
assign v$G33_8740_out0 = !((v$A0_923_out0 && !v$B0_2366_out0) || (!v$A0_923_out0) && v$B0_2366_out0);
assign v$_8853_out0 = v$IN_6534_out0[3:0];
assign v$_8856_out0 = v$IN_6538_out0[3:0];
assign v$G15_9198_out0 = !((v$A2_5567_out0 && !v$B2_11699_out0) || (!v$A2_5567_out0) && v$B2_11699_out0);
assign v$G15_9201_out0 = !((v$A2_5570_out0 && !v$B2_11702_out0) || (!v$A2_5570_out0) && v$B2_11702_out0);
assign v$G15_9210_out0 = !((v$A2_5579_out0 && !v$B2_11711_out0) || (!v$A2_5579_out0) && v$B2_11711_out0);
assign v$G15_9213_out0 = !((v$A2_5582_out0 && !v$B2_11714_out0) || (!v$A2_5582_out0) && v$B2_11714_out0);
assign v$G1_9792_out0 = v$SEL1_4765_out0 && v$SEL2_11054_out0;
assign v$G35_9914_out0 = !((v$A2_5567_out0 && !v$B2_11699_out0) || (!v$A2_5567_out0) && v$B2_11699_out0);
assign v$G35_9917_out0 = !((v$A2_5570_out0 && !v$B2_11702_out0) || (!v$A2_5570_out0) && v$B2_11702_out0);
assign v$G35_9926_out0 = !((v$A2_5579_out0 && !v$B2_11711_out0) || (!v$A2_5579_out0) && v$B2_11711_out0);
assign v$G35_9929_out0 = !((v$A2_5582_out0 && !v$B2_11714_out0) || (!v$A2_5582_out0) && v$B2_11714_out0);
assign v$_9978_out0 = v$IN_6534_out0[15:4];
assign v$_9982_out0 = v$IN_6538_out0[15:4];
assign v$_10004_out0 = v$IN_6534_out0[15:4];
assign v$_10008_out0 = v$IN_6538_out0[15:4];
assign v$G31_10788_out0 = v$A2$COMP$B2_1116_out0 || v$G32_322_out0;
assign v$G31_10789_out0 = v$A2$COMP$B2_1117_out0 || v$G32_323_out0;
assign v$G31_10800_out0 = v$A2$COMP$B2_1128_out0 || v$G32_334_out0;
assign v$G31_10801_out0 = v$A2$COMP$B2_1129_out0 || v$G32_335_out0;
assign v$G6_10840_out0 = ! v$R_13039_out0;
assign v$G6_10851_out0 = ! v$R_13050_out0;
assign v$G12_11549_out0 = ! v$B2_11699_out0;
assign v$G12_11552_out0 = ! v$B2_11702_out0;
assign v$G12_11561_out0 = ! v$B2_11711_out0;
assign v$G12_11564_out0 = ! v$B2_11714_out0;
assign v$_11796_out0 = v$IN_6534_out0[15:4];
assign v$_11800_out0 = v$IN_6538_out0[15:4];
assign v$G16_11914_out0 = !((v$A1_9729_out0 && !v$B1_9620_out0) || (!v$A1_9729_out0) && v$B1_9620_out0);
assign v$G16_11917_out0 = !((v$A1_9732_out0 && !v$B1_9623_out0) || (!v$A1_9732_out0) && v$B1_9623_out0);
assign v$G16_11926_out0 = !((v$A1_9741_out0 && !v$B1_9632_out0) || (!v$A1_9741_out0) && v$B1_9632_out0);
assign v$G16_11929_out0 = !((v$A1_9744_out0 && !v$B1_9635_out0) || (!v$A1_9744_out0) && v$B1_9635_out0);
assign v$S_11989_out0 = v$TXSet_8294_out0;
assign v$S_12000_out0 = v$TXSet_8295_out0;
assign v$G34_12124_out0 = !((v$A1_9729_out0 && !v$B1_9620_out0) || (!v$A1_9729_out0) && v$B1_9620_out0);
assign v$G34_12127_out0 = !((v$A1_9732_out0 && !v$B1_9623_out0) || (!v$A1_9732_out0) && v$B1_9623_out0);
assign v$G34_12136_out0 = !((v$A1_9741_out0 && !v$B1_9632_out0) || (!v$A1_9741_out0) && v$B1_9632_out0);
assign v$G34_12139_out0 = !((v$A1_9744_out0 && !v$B1_9635_out0) || (!v$A1_9744_out0) && v$B1_9635_out0);
assign v$R_13040_out0 = v$Clear_10010_out0;
assign v$R_13041_out0 = v$Clear_10010_out0;
assign v$R_13042_out0 = v$Clear_10010_out0;
assign v$R_13051_out0 = v$Clear_10011_out0;
assign v$R_13052_out0 = v$Clear_10011_out0;
assign v$R_13053_out0 = v$Clear_10011_out0;
assign v$SAME_13065_out0 = v$SAME_13352_out0;
assign v$SAME_13069_out0 = v$SAME_13368_out0;
assign v$SAME_13365_out0 = v$G41_7166_out0;
assign v$SAME_13366_out0 = v$G41_7167_out0;
assign v$SAME_13381_out0 = v$G41_7178_out0;
assign v$SAME_13382_out0 = v$G41_7179_out0;
assign v$MUX1_345_out0 = v$G17_6145_out0 ? v$FF2_1717_out0 : v$_2193_out0;
assign v$MUX1_346_out0 = v$G17_6146_out0 ? v$FF2_1718_out0 : v$_2194_out0;
assign v$G5_424_out0 = v$FF2_8669_out0 && v$G6_10840_out0;
assign v$G5_429_out0 = v$FF2_8680_out0 && v$G6_10851_out0;
assign v$A0XNORB0_672_out0 = v$G17_5673_out0;
assign v$A0XNORB0_675_out0 = v$G17_5676_out0;
assign v$A0XNORB0_684_out0 = v$G17_5685_out0;
assign v$A0XNORB0_687_out0 = v$G17_5688_out0;
assign v$_711_out0 = { v$C1_5480_out0,v$_3211_out0 };
assign v$_715_out0 = { v$C1_5484_out0,v$_3215_out0 };
assign v$MUX8_725_out0 = v$G17_6145_out0 ? v$C1_8496_out0 : v$_6383_out1;
assign v$MUX8_726_out0 = v$G17_6146_out0 ? v$C1_8497_out0 : v$_6384_out1;
assign v$G30_949_out0 = v$A3$COMP$B3_3339_out0 || v$G31_10788_out0;
assign v$G30_950_out0 = v$A3$COMP$B3_3340_out0 || v$G31_10789_out0;
assign v$G30_961_out0 = v$A3$COMP$B3_3351_out0 || v$G31_10800_out0;
assign v$G30_962_out0 = v$A3$COMP$B3_3352_out0 || v$G31_10801_out0;
assign v$MUX3_2097_out0 = v$OUT_2622_out0 ? v$A$EXP_236_out0 : v$B$EXP_11734_out0;
assign v$MUX3_2101_out0 = v$OUT_2638_out0 ? v$A$EXP_240_out0 : v$B$EXP_11738_out0;
assign v$B0_2352_out0 = v$SEL10_8252_out0;
assign v$B0_2353_out0 = v$SEL10_8253_out0;
assign v$B0_2355_out0 = v$SEL10_8255_out0;
assign v$B0_2356_out0 = v$SEL10_8256_out0;
assign v$B0_2364_out0 = v$SEL10_8264_out0;
assign v$B0_2365_out0 = v$SEL10_8265_out0;
assign v$B0_2367_out0 = v$SEL10_8267_out0;
assign v$B0_2368_out0 = v$SEL10_8268_out0;
assign v$A2XNORB2_3128_out0 = v$G15_9198_out0;
assign v$A2XNORB2_3131_out0 = v$G15_9201_out0;
assign v$A2XNORB2_3140_out0 = v$G15_9210_out0;
assign v$A2XNORB2_3143_out0 = v$G15_9213_out0;
assign v$G5_3817_out0 = v$G1_9792_out0 && v$G2_7517_out0;
assign v$G5_4707_out0 = v$A3_7021_out0 && v$G6_4557_out0;
assign v$G5_4710_out0 = v$A3_7024_out0 && v$G6_4560_out0;
assign v$G5_4719_out0 = v$A3_7033_out0 && v$G6_4569_out0;
assign v$G5_4722_out0 = v$A3_7036_out0 && v$G6_4572_out0;
assign v$G38_4892_out0 = v$G33_8725_out0 && v$G34_12124_out0;
assign v$G38_4895_out0 = v$G33_8728_out0 && v$G34_12127_out0;
assign v$G38_4904_out0 = v$G33_8737_out0 && v$G34_12136_out0;
assign v$G38_4907_out0 = v$G33_8740_out0 && v$G34_12139_out0;
assign v$G2_5115_out0 = v$G1_8621_out0 || v$S_5522_out0;
assign v$G2_5116_out0 = v$G1_8622_out0 || v$S_5523_out0;
assign v$MUX6_6364_out0 = v$G17_6145_out0 ? v$FF7_12855_out0 : v$_5597_out1;
assign v$MUX6_6365_out0 = v$G17_6146_out0 ? v$FF7_12856_out0 : v$_5598_out1;
assign v$_6443_out0 = { v$_11796_out0,v$LSBS_10623_out0 };
assign v$_6447_out0 = { v$_11800_out0,v$LSBS_10624_out0 };
assign v$MUX7_6471_out0 = v$G17_6145_out0 ? v$FF8_5529_out0 : v$_6383_out0;
assign v$MUX7_6472_out0 = v$G17_6146_out0 ? v$FF8_5530_out0 : v$_6384_out0;
assign v$G20_6622_out0 = v$A1_9729_out0 && v$G21_2227_out0;
assign v$G20_6625_out0 = v$A1_9732_out0 && v$G21_2230_out0;
assign v$G20_6634_out0 = v$A1_9741_out0 && v$G21_2239_out0;
assign v$G20_6637_out0 = v$A1_9744_out0 && v$G21_2242_out0;
assign v$_6643_out0 = { v$_765_out0,v$_765_out0 };
assign v$_6644_out0 = { v$_766_out0,v$_766_out0 };
assign v$LOWER$SAME_6760_out0 = v$SAME_13366_out0;
assign v$LOWER$SAME_6764_out0 = v$SAME_13382_out0;
assign v$G25_7206_out0 = v$A0_908_out0 && v$G23_7951_out0;
assign v$G25_7209_out0 = v$A0_911_out0 && v$G23_7954_out0;
assign v$G25_7218_out0 = v$A0_920_out0 && v$G23_7963_out0;
assign v$G25_7221_out0 = v$A0_923_out0 && v$G23_7966_out0;
assign v$MUX4_7488_out0 = v$IS$32$BITS_527_out0 ? v$SAME_13065_out0 : v$SAME_13064_out0;
assign v$MUX4_7489_out0 = v$IS$32$BITS_528_out0 ? v$SAME_13069_out0 : v$SAME_13068_out0;
assign v$G4_7633_out0 = v$G5_423_out0 || v$S_11989_out0;
assign v$G4_7638_out0 = v$G5_428_out0 || v$S_12000_out0;
assign v$A1$COMP$B1_8137_out0 = v$G18_3376_out0;
assign v$A1$COMP$B1_8138_out0 = v$G18_3377_out0;
assign v$A1$COMP$B1_8149_out0 = v$G18_3388_out0;
assign v$A1$COMP$B1_8150_out0 = v$G18_3389_out0;
assign v$MUX2_8870_out0 = v$G17_6145_out0 ? v$FF3_227_out0 : v$_2193_out1;
assign v$MUX2_8871_out0 = v$G17_6146_out0 ? v$FF3_228_out0 : v$_2194_out1;
assign v$_8879_out0 = { v$_9978_out0,v$_8853_out0 };
assign v$_8883_out0 = { v$_9982_out0,v$_8856_out0 };
assign v$G40_8937_out0 = v$G35_9914_out0 && v$G36_3926_out0;
assign v$G40_8940_out0 = v$G35_9917_out0 && v$G36_3929_out0;
assign v$G40_8949_out0 = v$G35_9926_out0 && v$G36_3938_out0;
assign v$G40_8952_out0 = v$G35_9929_out0 && v$G36_3941_out0;
assign v$OUT_9286_out0 = v$OUT_2622_out0;
assign v$OUT_9290_out0 = v$OUT_2638_out0;
assign v$B1_9621_out0 = v$SEL9_7132_out0;
assign v$B1_9622_out0 = v$SEL9_7133_out0;
assign v$B1_9624_out0 = v$SEL9_7135_out0;
assign v$B1_9625_out0 = v$SEL9_7136_out0;
assign v$B1_9633_out0 = v$SEL9_7144_out0;
assign v$B1_9634_out0 = v$SEL9_7145_out0;
assign v$B1_9636_out0 = v$SEL9_7147_out0;
assign v$B1_9637_out0 = v$SEL9_7148_out0;
assign v$MUX5_9877_out0 = v$S_6897_out0 ? v$_4977_out0 : v$C1_8474_out0;
assign v$MUX5_9878_out0 = v$S_6898_out0 ? v$_4978_out0 : v$C1_8475_out0;
assign v$A3XNORB3_10075_out0 = v$G8_2442_out0;
assign v$A3XNORB3_10078_out0 = v$G8_2445_out0;
assign v$A3XNORB3_10087_out0 = v$G8_2454_out0;
assign v$A3XNORB3_10090_out0 = v$G8_2457_out0;
assign v$HIGHER$SAME_10334_out0 = v$SAME_13365_out0;
assign v$HIGHER$SAME_10338_out0 = v$SAME_13381_out0;
assign v$G31_10796_out0 = v$A2$COMP$B2_1124_out0 || v$G32_330_out0;
assign v$G31_10808_out0 = v$A2$COMP$B2_1136_out0 || v$G32_342_out0;
assign v$G6_10841_out0 = ! v$R_13040_out0;
assign v$G6_10842_out0 = ! v$R_13041_out0;
assign v$G6_10843_out0 = ! v$R_13042_out0;
assign v$G6_10852_out0 = ! v$R_13051_out0;
assign v$G6_10853_out0 = ! v$R_13052_out0;
assign v$G6_10854_out0 = ! v$R_13053_out0;
assign v$MUX4_10904_out0 = v$G17_6145_out0 ? v$FF5_11452_out0 : v$_9470_out1;
assign v$MUX4_10905_out0 = v$G17_6146_out0 ? v$FF5_11453_out0 : v$_9471_out1;
assign v$G11_10909_out0 = v$A2_5567_out0 && v$G12_11549_out0;
assign v$G11_10912_out0 = v$A2_5570_out0 && v$G12_11552_out0;
assign v$G11_10921_out0 = v$A2_5579_out0 && v$G12_11561_out0;
assign v$G11_10924_out0 = v$A2_5582_out0 && v$G12_11564_out0;
assign v$G24_10957_out0 = v$A3XNORB3_10082_out0 && v$G27_3195_out0;
assign v$G24_10958_out0 = v$A3XNORB3_10083_out0 && v$G27_3196_out0;
assign v$G24_10969_out0 = v$A3XNORB3_10094_out0 && v$G27_3207_out0;
assign v$G24_10970_out0 = v$A3XNORB3_10095_out0 && v$G27_3208_out0;
assign v$A1XNORB1_11228_out0 = v$G16_11914_out0;
assign v$A1XNORB1_11231_out0 = v$G16_11917_out0;
assign v$A1XNORB1_11240_out0 = v$G16_11926_out0;
assign v$A1XNORB1_11243_out0 = v$G16_11929_out0;
assign v$B2_11700_out0 = v$SEL8_8563_out0;
assign v$B2_11701_out0 = v$SEL8_8564_out0;
assign v$B2_11703_out0 = v$SEL8_8566_out0;
assign v$B2_11704_out0 = v$SEL8_8567_out0;
assign v$B2_11712_out0 = v$SEL8_8575_out0;
assign v$B2_11713_out0 = v$SEL8_8576_out0;
assign v$B2_11715_out0 = v$SEL8_8578_out0;
assign v$B2_11716_out0 = v$SEL8_8579_out0;
assign v$S_11991_out0 = v$G9_5922_out0;
assign v$S_12002_out0 = v$G9_5923_out0;
assign v$G6_12207_out0 = v$G3_3394_out0 && v$G4_4429_out0;
assign v$MUX3_12536_out0 = v$G17_6145_out0 ? v$FF4_1281_out0 : v$_9470_out0;
assign v$MUX3_12537_out0 = v$G17_6146_out0 ? v$FF4_1282_out0 : v$_9471_out0;
assign v$B3_12642_out0 = v$SEL7_2860_out0;
assign v$B3_12643_out0 = v$SEL7_2861_out0;
assign v$B3_12645_out0 = v$SEL7_2863_out0;
assign v$B3_12646_out0 = v$SEL7_2864_out0;
assign v$B3_12654_out0 = v$SEL7_2872_out0;
assign v$B3_12655_out0 = v$SEL7_2873_out0;
assign v$B3_12657_out0 = v$SEL7_2875_out0;
assign v$B3_12658_out0 = v$SEL7_2876_out0;
assign v$MUX1_12699_out0 = v$OUT_2622_out0 ? v$B$EXP_11734_out0 : v$A$EXP_236_out0;
assign v$MUX1_12703_out0 = v$OUT_2638_out0 ? v$B$EXP_11738_out0 : v$A$EXP_240_out0;
assign v$MUX5_13207_out0 = v$G17_6145_out0 ? v$FF6_10631_out0 : v$_5597_out0;
assign v$MUX5_13208_out0 = v$G17_6146_out0 ? v$FF6_10632_out0 : v$_5598_out0;
assign v$G5_425_out0 = v$FF2_8670_out0 && v$G6_10841_out0;
assign v$G5_426_out0 = v$FF2_8671_out0 && v$G6_10842_out0;
assign v$G5_427_out0 = v$FF2_8672_out0 && v$G6_10843_out0;
assign v$G5_430_out0 = v$FF2_8681_out0 && v$G6_10852_out0;
assign v$G5_431_out0 = v$FF2_8682_out0 && v$G6_10853_out0;
assign v$G5_432_out0 = v$FF2_8683_out0 && v$G6_10854_out0;
assign v$G30_957_out0 = v$A3$COMP$B3_3347_out0 || v$G31_10796_out0;
assign v$G30_969_out0 = v$A3$COMP$B3_3359_out0 || v$G31_10808_out0;
assign v$G21_2228_out0 = ! v$B1_9621_out0;
assign v$G21_2229_out0 = ! v$B1_9622_out0;
assign v$G21_2231_out0 = ! v$B1_9624_out0;
assign v$G21_2232_out0 = ! v$B1_9625_out0;
assign v$G21_2240_out0 = ! v$B1_9633_out0;
assign v$G21_2241_out0 = ! v$B1_9634_out0;
assign v$G21_2243_out0 = ! v$B1_9636_out0;
assign v$G21_2244_out0 = ! v$B1_9637_out0;
assign v$G8_2443_out0 = !((v$A3_7022_out0 && !v$B3_12642_out0) || (!v$A3_7022_out0) && v$B3_12642_out0);
assign v$G8_2444_out0 = !((v$A3_7023_out0 && !v$B3_12643_out0) || (!v$A3_7023_out0) && v$B3_12643_out0);
assign v$G8_2446_out0 = !((v$A3_7025_out0 && !v$B3_12645_out0) || (!v$A3_7025_out0) && v$B3_12645_out0);
assign v$G8_2447_out0 = !((v$A3_7026_out0 && !v$B3_12646_out0) || (!v$A3_7026_out0) && v$B3_12646_out0);
assign v$G8_2455_out0 = !((v$A3_7034_out0 && !v$B3_12654_out0) || (!v$A3_7034_out0) && v$B3_12654_out0);
assign v$G8_2456_out0 = !((v$A3_7035_out0 && !v$B3_12655_out0) || (!v$A3_7035_out0) && v$B3_12655_out0);
assign v$G8_2458_out0 = !((v$A3_7037_out0 && !v$B3_12657_out0) || (!v$A3_7037_out0) && v$B3_12657_out0);
assign v$G8_2459_out0 = !((v$A3_7038_out0 && !v$B3_12658_out0) || (!v$A3_7038_out0) && v$B3_12658_out0);
assign v$OUT_2624_out0 = v$G30_949_out0;
assign v$OUT_2625_out0 = v$G30_950_out0;
assign v$OUT_2640_out0 = v$G30_961_out0;
assign v$OUT_2641_out0 = v$G30_962_out0;
assign v$G13_3057_out0 = v$A3XNORB3_10075_out0 && v$G11_10909_out0;
assign v$G13_3060_out0 = v$A3XNORB3_10078_out0 && v$G11_10912_out0;
assign v$G13_3069_out0 = v$A3XNORB3_10087_out0 && v$G11_10921_out0;
assign v$G13_3072_out0 = v$A3XNORB3_10090_out0 && v$G11_10924_out0;
assign v$A3$COMP$B3_3341_out0 = v$G5_4707_out0;
assign v$A3$COMP$B3_3344_out0 = v$G5_4710_out0;
assign v$A3$COMP$B3_3353_out0 = v$G5_4719_out0;
assign v$A3$COMP$B3_3356_out0 = v$G5_4722_out0;
assign v$G36_3927_out0 = !((v$B3_12642_out0 && !v$A3_7022_out0) || (!v$B3_12642_out0) && v$A3_7022_out0);
assign v$G36_3928_out0 = !((v$B3_12643_out0 && !v$A3_7023_out0) || (!v$B3_12643_out0) && v$A3_7023_out0);
assign v$G36_3930_out0 = !((v$B3_12645_out0 && !v$A3_7025_out0) || (!v$B3_12645_out0) && v$A3_7025_out0);
assign v$G36_3931_out0 = !((v$B3_12646_out0 && !v$A3_7026_out0) || (!v$B3_12646_out0) && v$A3_7026_out0);
assign v$G36_3939_out0 = !((v$B3_12654_out0 && !v$A3_7034_out0) || (!v$B3_12654_out0) && v$A3_7034_out0);
assign v$G36_3940_out0 = !((v$B3_12655_out0 && !v$A3_7035_out0) || (!v$B3_12655_out0) && v$A3_7035_out0);
assign v$G36_3942_out0 = !((v$B3_12657_out0 && !v$A3_7037_out0) || (!v$B3_12657_out0) && v$A3_7037_out0);
assign v$G36_3943_out0 = !((v$B3_12658_out0 && !v$A3_7038_out0) || (!v$B3_12658_out0) && v$A3_7038_out0);
assign v$G6_4558_out0 = ! v$B3_12642_out0;
assign v$G6_4559_out0 = ! v$B3_12643_out0;
assign v$G6_4561_out0 = ! v$B3_12645_out0;
assign v$G6_4562_out0 = ! v$B3_12646_out0;
assign v$G6_4570_out0 = ! v$B3_12654_out0;
assign v$G6_4571_out0 = ! v$B3_12655_out0;
assign v$G6_4573_out0 = ! v$B3_12657_out0;
assign v$G6_4574_out0 = ! v$B3_12658_out0;
assign v$_5102_out0 = { v$_6643_out0,v$_6643_out0 };
assign v$_5103_out0 = { v$_6644_out0,v$_6644_out0 };
assign v$XOR1_5128_out0 = v$C1_9147_out0 ^ v$MUX1_12699_out0;
assign v$XOR1_5132_out0 = v$C1_9151_out0 ^ v$MUX1_12703_out0;
assign v$A0$COMP$B0_5502_out0 = v$G24_10957_out0;
assign v$A0$COMP$B0_5503_out0 = v$G24_10958_out0;
assign v$A0$COMP$B0_5514_out0 = v$G24_10969_out0;
assign v$A0$COMP$B0_5515_out0 = v$G24_10970_out0;
assign v$G17_5674_out0 = !((v$A0_909_out0 && !v$B0_2352_out0) || (!v$A0_909_out0) && v$B0_2352_out0);
assign v$G17_5675_out0 = !((v$A0_910_out0 && !v$B0_2353_out0) || (!v$A0_910_out0) && v$B0_2353_out0);
assign v$G17_5677_out0 = !((v$A0_912_out0 && !v$B0_2355_out0) || (!v$A0_912_out0) && v$B0_2355_out0);
assign v$G17_5678_out0 = !((v$A0_913_out0 && !v$B0_2356_out0) || (!v$A0_913_out0) && v$B0_2356_out0);
assign v$G17_5686_out0 = !((v$A0_921_out0 && !v$B0_2364_out0) || (!v$A0_921_out0) && v$B0_2364_out0);
assign v$G17_5687_out0 = !((v$A0_922_out0 && !v$B0_2365_out0) || (!v$A0_922_out0) && v$B0_2365_out0);
assign v$G17_5689_out0 = !((v$A0_924_out0 && !v$B0_2367_out0) || (!v$A0_924_out0) && v$B0_2367_out0);
assign v$G17_5690_out0 = !((v$A0_925_out0 && !v$B0_2368_out0) || (!v$A0_925_out0) && v$B0_2368_out0);
assign v$G1_6390_out0 = v$LOWER$SAME_6760_out0 && v$HIGHER$SAME_10334_out0;
assign v$G1_6394_out0 = v$LOWER$SAME_6764_out0 && v$HIGHER$SAME_10338_out0;
assign v$G41_7159_out0 = v$G38_4892_out0 && v$G40_8937_out0;
assign v$G41_7162_out0 = v$G38_4895_out0 && v$G40_8940_out0;
assign v$G41_7171_out0 = v$G38_4904_out0 && v$G40_8949_out0;
assign v$G41_7174_out0 = v$G38_4907_out0 && v$G40_8952_out0;
assign v$G4_7634_out0 = v$G5_424_out0 || v$S_11990_out0;
assign v$G4_7639_out0 = v$G5_429_out0 || v$S_12001_out0;
assign v$G23_7952_out0 = ! v$B0_2352_out0;
assign v$G23_7953_out0 = ! v$B0_2353_out0;
assign v$G23_7955_out0 = ! v$B0_2355_out0;
assign v$G23_7956_out0 = ! v$B0_2356_out0;
assign v$G23_7964_out0 = ! v$B0_2364_out0;
assign v$G23_7965_out0 = ! v$B0_2365_out0;
assign v$G23_7967_out0 = ! v$B0_2367_out0;
assign v$G23_7968_out0 = ! v$B0_2368_out0;
assign v$G28_8641_out0 = v$A1XNORB1_11228_out0 && v$G25_7206_out0;
assign v$G28_8644_out0 = v$A1XNORB1_11231_out0 && v$G25_7209_out0;
assign v$G28_8653_out0 = v$A1XNORB1_11240_out0 && v$G25_7218_out0;
assign v$G28_8656_out0 = v$A1XNORB1_11243_out0 && v$G25_7221_out0;
assign v$G33_8726_out0 = !((v$A0_909_out0 && !v$B0_2352_out0) || (!v$A0_909_out0) && v$B0_2352_out0);
assign v$G33_8727_out0 = !((v$A0_910_out0 && !v$B0_2353_out0) || (!v$A0_910_out0) && v$B0_2353_out0);
assign v$G33_8729_out0 = !((v$A0_912_out0 && !v$B0_2355_out0) || (!v$A0_912_out0) && v$B0_2355_out0);
assign v$G33_8730_out0 = !((v$A0_913_out0 && !v$B0_2356_out0) || (!v$A0_913_out0) && v$B0_2356_out0);
assign v$G33_8738_out0 = !((v$A0_921_out0 && !v$B0_2364_out0) || (!v$A0_921_out0) && v$B0_2364_out0);
assign v$G33_8739_out0 = !((v$A0_922_out0 && !v$B0_2365_out0) || (!v$A0_922_out0) && v$B0_2365_out0);
assign v$G33_8741_out0 = !((v$A0_924_out0 && !v$B0_2367_out0) || (!v$A0_924_out0) && v$B0_2367_out0);
assign v$G33_8742_out0 = !((v$A0_925_out0 && !v$B0_2368_out0) || (!v$A0_925_out0) && v$B0_2368_out0);
assign v$G22_8904_out0 = v$A2XNORB2_3128_out0 && v$G20_6622_out0;
assign v$G22_8907_out0 = v$A2XNORB2_3131_out0 && v$G20_6625_out0;
assign v$G22_8916_out0 = v$A2XNORB2_3140_out0 && v$G20_6634_out0;
assign v$G22_8919_out0 = v$A2XNORB2_3143_out0 && v$G20_6637_out0;
assign v$NEXTSTATE_9107_out0 = v$G2_5115_out0;
assign v$NEXTSTATE_9108_out0 = v$G2_5116_out0;
assign v$G15_9199_out0 = !((v$A2_5568_out0 && !v$B2_11700_out0) || (!v$A2_5568_out0) && v$B2_11700_out0);
assign v$G15_9200_out0 = !((v$A2_5569_out0 && !v$B2_11701_out0) || (!v$A2_5569_out0) && v$B2_11701_out0);
assign v$G15_9202_out0 = !((v$A2_5571_out0 && !v$B2_11703_out0) || (!v$A2_5571_out0) && v$B2_11703_out0);
assign v$G15_9203_out0 = !((v$A2_5572_out0 && !v$B2_11704_out0) || (!v$A2_5572_out0) && v$B2_11704_out0);
assign v$G15_9211_out0 = !((v$A2_5580_out0 && !v$B2_11712_out0) || (!v$A2_5580_out0) && v$B2_11712_out0);
assign v$G15_9212_out0 = !((v$A2_5581_out0 && !v$B2_11713_out0) || (!v$A2_5581_out0) && v$B2_11713_out0);
assign v$G15_9214_out0 = !((v$A2_5583_out0 && !v$B2_11715_out0) || (!v$A2_5583_out0) && v$B2_11715_out0);
assign v$G15_9215_out0 = !((v$A2_5584_out0 && !v$B2_11716_out0) || (!v$A2_5584_out0) && v$B2_11716_out0);
assign v$Q_9534_out0 = v$G4_7633_out0;
assign v$Q_9545_out0 = v$G4_7638_out0;
assign v$G35_9915_out0 = !((v$A2_5568_out0 && !v$B2_11700_out0) || (!v$A2_5568_out0) && v$B2_11700_out0);
assign v$G35_9916_out0 = !((v$A2_5569_out0 && !v$B2_11701_out0) || (!v$A2_5569_out0) && v$B2_11701_out0);
assign v$G35_9918_out0 = !((v$A2_5571_out0 && !v$B2_11703_out0) || (!v$A2_5571_out0) && v$B2_11703_out0);
assign v$G35_9919_out0 = !((v$A2_5572_out0 && !v$B2_11704_out0) || (!v$A2_5572_out0) && v$B2_11704_out0);
assign v$G35_9927_out0 = !((v$A2_5580_out0 && !v$B2_11712_out0) || (!v$A2_5580_out0) && v$B2_11712_out0);
assign v$G35_9928_out0 = !((v$A2_5581_out0 && !v$B2_11713_out0) || (!v$A2_5581_out0) && v$B2_11713_out0);
assign v$G35_9930_out0 = !((v$A2_5583_out0 && !v$B2_11715_out0) || (!v$A2_5583_out0) && v$B2_11715_out0);
assign v$G35_9931_out0 = !((v$A2_5584_out0 && !v$B2_11716_out0) || (!v$A2_5584_out0) && v$B2_11716_out0);
assign v$G7_10153_out0 = v$G5_3817_out0 && v$G6_12207_out0;
assign v$MUX4_11180_out0 = v$EN_12031_out0 ? v$_711_out0 : v$IN_6534_out0;
assign v$MUX4_11184_out0 = v$EN_12035_out0 ? v$_715_out0 : v$IN_6538_out0;
assign v$G12_11550_out0 = ! v$B2_11700_out0;
assign v$G12_11551_out0 = ! v$B2_11701_out0;
assign v$G12_11553_out0 = ! v$B2_11703_out0;
assign v$G12_11554_out0 = ! v$B2_11704_out0;
assign v$G12_11562_out0 = ! v$B2_11712_out0;
assign v$G12_11563_out0 = ! v$B2_11713_out0;
assign v$G12_11565_out0 = ! v$B2_11715_out0;
assign v$G12_11566_out0 = ! v$B2_11716_out0;
assign v$EXP$SAME_11626_out0 = v$MUX4_7488_out0;
assign v$EXP$SAME_11627_out0 = v$MUX4_7489_out0;
assign v$G16_11915_out0 = !((v$A1_9730_out0 && !v$B1_9621_out0) || (!v$A1_9730_out0) && v$B1_9621_out0);
assign v$G16_11916_out0 = !((v$A1_9731_out0 && !v$B1_9622_out0) || (!v$A1_9731_out0) && v$B1_9622_out0);
assign v$G16_11918_out0 = !((v$A1_9733_out0 && !v$B1_9624_out0) || (!v$A1_9733_out0) && v$B1_9624_out0);
assign v$G16_11919_out0 = !((v$A1_9734_out0 && !v$B1_9625_out0) || (!v$A1_9734_out0) && v$B1_9625_out0);
assign v$G16_11927_out0 = !((v$A1_9742_out0 && !v$B1_9633_out0) || (!v$A1_9742_out0) && v$B1_9633_out0);
assign v$G16_11928_out0 = !((v$A1_9743_out0 && !v$B1_9634_out0) || (!v$A1_9743_out0) && v$B1_9634_out0);
assign v$G16_11930_out0 = !((v$A1_9745_out0 && !v$B1_9636_out0) || (!v$A1_9745_out0) && v$B1_9636_out0);
assign v$G16_11931_out0 = !((v$A1_9746_out0 && !v$B1_9637_out0) || (!v$A1_9746_out0) && v$B1_9637_out0);
assign v$G34_12125_out0 = !((v$A1_9730_out0 && !v$B1_9621_out0) || (!v$A1_9730_out0) && v$B1_9621_out0);
assign v$G34_12126_out0 = !((v$A1_9731_out0 && !v$B1_9622_out0) || (!v$A1_9731_out0) && v$B1_9622_out0);
assign v$G34_12128_out0 = !((v$A1_9733_out0 && !v$B1_9624_out0) || (!v$A1_9733_out0) && v$B1_9624_out0);
assign v$G34_12129_out0 = !((v$A1_9734_out0 && !v$B1_9625_out0) || (!v$A1_9734_out0) && v$B1_9625_out0);
assign v$G34_12137_out0 = !((v$A1_9742_out0 && !v$B1_9633_out0) || (!v$A1_9742_out0) && v$B1_9633_out0);
assign v$G34_12138_out0 = !((v$A1_9743_out0 && !v$B1_9634_out0) || (!v$A1_9743_out0) && v$B1_9634_out0);
assign v$G34_12140_out0 = !((v$A1_9745_out0 && !v$B1_9636_out0) || (!v$A1_9745_out0) && v$B1_9636_out0);
assign v$G34_12141_out0 = !((v$A1_9746_out0 && !v$B1_9637_out0) || (!v$A1_9746_out0) && v$B1_9637_out0);
assign v$G32_331_out0 = v$A1$COMP$B1_8137_out0 || v$A0$COMP$B0_5502_out0;
assign v$G32_332_out0 = v$A1$COMP$B1_8138_out0 || v$A0$COMP$B0_5503_out0;
assign v$G32_343_out0 = v$A1$COMP$B1_8149_out0 || v$A0$COMP$B0_5514_out0;
assign v$G32_344_out0 = v$A1$COMP$B1_8150_out0 || v$A0$COMP$B0_5515_out0;
assign v$A0XNORB0_673_out0 = v$G17_5674_out0;
assign v$A0XNORB0_674_out0 = v$G17_5675_out0;
assign v$A0XNORB0_676_out0 = v$G17_5677_out0;
assign v$A0XNORB0_677_out0 = v$G17_5678_out0;
assign v$A0XNORB0_685_out0 = v$G17_5686_out0;
assign v$A0XNORB0_686_out0 = v$G17_5687_out0;
assign v$A0XNORB0_688_out0 = v$G17_5689_out0;
assign v$A0XNORB0_689_out0 = v$G17_5690_out0;
assign v$A2$COMP$B2_1118_out0 = v$G13_3057_out0;
assign v$A2$COMP$B2_1121_out0 = v$G13_3060_out0;
assign v$A2$COMP$B2_1130_out0 = v$G13_3069_out0;
assign v$A2$COMP$B2_1133_out0 = v$G13_3072_out0;
assign v$MUX6_1605_out0 = v$FF1_9226_out0 ? v$LSBS_10623_out0 : v$_5102_out0;
assign v$MUX6_1606_out0 = v$FF1_9227_out0 ? v$LSBS_10624_out0 : v$_5103_out0;
assign v$HIGHER$OUT_2537_out0 = v$OUT_2624_out0;
assign v$HIGHER$OUT_2541_out0 = v$OUT_2640_out0;
assign v$LOWER$OUT_2902_out0 = v$OUT_2625_out0;
assign v$LOWER$OUT_2906_out0 = v$OUT_2641_out0;
assign v$A2XNORB2_3129_out0 = v$G15_9199_out0;
assign v$A2XNORB2_3130_out0 = v$G15_9200_out0;
assign v$A2XNORB2_3132_out0 = v$G15_9202_out0;
assign v$A2XNORB2_3133_out0 = v$G15_9203_out0;
assign v$A2XNORB2_3141_out0 = v$G15_9211_out0;
assign v$A2XNORB2_3142_out0 = v$G15_9212_out0;
assign v$A2XNORB2_3144_out0 = v$G15_9214_out0;
assign v$A2XNORB2_3145_out0 = v$G15_9215_out0;
assign v$G27_3188_out0 = v$A2XNORB2_3128_out0 && v$G28_8641_out0;
assign v$G27_3191_out0 = v$A2XNORB2_3131_out0 && v$G28_8644_out0;
assign v$G27_3200_out0 = v$A2XNORB2_3140_out0 && v$G28_8653_out0;
assign v$G27_3203_out0 = v$A2XNORB2_3143_out0 && v$G28_8656_out0;
assign v$G18_3369_out0 = v$A3XNORB3_10075_out0 && v$G22_8904_out0;
assign v$G18_3372_out0 = v$A3XNORB3_10078_out0 && v$G22_8907_out0;
assign v$G18_3381_out0 = v$A3XNORB3_10087_out0 && v$G22_8916_out0;
assign v$G18_3384_out0 = v$A3XNORB3_10090_out0 && v$G22_8919_out0;
assign {v$A1_3809_out1,v$A1_3809_out0 } = v$MUX3_2097_out0 + v$XOR1_5128_out0 + v$CIN_12952_out0;
assign {v$A1_3813_out1,v$A1_3813_out0 } = v$MUX3_2101_out0 + v$XOR1_5132_out0 + v$CIN_12956_out0;
assign v$G5_4708_out0 = v$A3_7022_out0 && v$G6_4558_out0;
assign v$G5_4709_out0 = v$A3_7023_out0 && v$G6_4559_out0;
assign v$G5_4711_out0 = v$A3_7025_out0 && v$G6_4561_out0;
assign v$G5_4712_out0 = v$A3_7026_out0 && v$G6_4562_out0;
assign v$G5_4720_out0 = v$A3_7034_out0 && v$G6_4570_out0;
assign v$G5_4721_out0 = v$A3_7035_out0 && v$G6_4571_out0;
assign v$G5_4723_out0 = v$A3_7037_out0 && v$G6_4573_out0;
assign v$G5_4724_out0 = v$A3_7038_out0 && v$G6_4574_out0;
assign v$G38_4893_out0 = v$G33_8726_out0 && v$G34_12125_out0;
assign v$G38_4894_out0 = v$G33_8727_out0 && v$G34_12126_out0;
assign v$G38_4896_out0 = v$G33_8729_out0 && v$G34_12128_out0;
assign v$G38_4897_out0 = v$G33_8730_out0 && v$G34_12129_out0;
assign v$G38_4905_out0 = v$G33_8738_out0 && v$G34_12137_out0;
assign v$G38_4906_out0 = v$G33_8739_out0 && v$G34_12138_out0;
assign v$G38_4908_out0 = v$G33_8741_out0 && v$G34_12140_out0;
assign v$G38_4909_out0 = v$G33_8742_out0 && v$G34_12141_out0;
assign v$TXFlag_5261_out0 = v$Q_9534_out0;
assign v$TXFlag_5262_out0 = v$Q_9545_out0;
assign v$IGNORE_5757_out0 = v$G7_10153_out0;
assign v$G20_6623_out0 = v$A1_9730_out0 && v$G21_2228_out0;
assign v$G20_6624_out0 = v$A1_9731_out0 && v$G21_2229_out0;
assign v$G20_6626_out0 = v$A1_9733_out0 && v$G21_2231_out0;
assign v$G20_6627_out0 = v$A1_9734_out0 && v$G21_2232_out0;
assign v$G20_6635_out0 = v$A1_9742_out0 && v$G21_2240_out0;
assign v$G20_6636_out0 = v$A1_9743_out0 && v$G21_2241_out0;
assign v$G20_6638_out0 = v$A1_9745_out0 && v$G21_2243_out0;
assign v$G20_6639_out0 = v$A1_9746_out0 && v$G21_2244_out0;
assign v$G29_6860_out0 = v$A4$COMP$B4_4998_out0 || v$G30_957_out0;
assign v$G29_6862_out0 = v$A4$COMP$B4_5000_out0 || v$G30_969_out0;
assign v$G25_7207_out0 = v$A0_909_out0 && v$G23_7952_out0;
assign v$G25_7208_out0 = v$A0_910_out0 && v$G23_7953_out0;
assign v$G25_7210_out0 = v$A0_912_out0 && v$G23_7955_out0;
assign v$G25_7211_out0 = v$A0_913_out0 && v$G23_7956_out0;
assign v$G25_7219_out0 = v$A0_921_out0 && v$G23_7964_out0;
assign v$G25_7220_out0 = v$A0_922_out0 && v$G23_7965_out0;
assign v$G25_7222_out0 = v$A0_924_out0 && v$G23_7967_out0;
assign v$G25_7223_out0 = v$A0_925_out0 && v$G23_7968_out0;
assign v$G4_7635_out0 = v$G5_425_out0 || v$S_11991_out0;
assign v$G4_7636_out0 = v$G5_426_out0 || v$S_11992_out0;
assign v$G4_7637_out0 = v$G5_427_out0 || v$S_11993_out0;
assign v$G4_7640_out0 = v$G5_430_out0 || v$S_12002_out0;
assign v$G4_7641_out0 = v$G5_431_out0 || v$S_12003_out0;
assign v$G4_7642_out0 = v$G5_432_out0 || v$S_12004_out0;
assign v$MUX2_7824_out0 = v$G3_1509_out0 ? v$_6443_out0 : v$MUX4_11180_out0;
assign v$MUX2_7828_out0 = v$G3_1513_out0 ? v$_6447_out0 : v$MUX4_11184_out0;
assign v$G40_8938_out0 = v$G35_9915_out0 && v$G36_3927_out0;
assign v$G40_8939_out0 = v$G35_9916_out0 && v$G36_3928_out0;
assign v$G40_8941_out0 = v$G35_9918_out0 && v$G36_3930_out0;
assign v$G40_8942_out0 = v$G35_9919_out0 && v$G36_3931_out0;
assign v$G40_8950_out0 = v$G35_9927_out0 && v$G36_3939_out0;
assign v$G40_8951_out0 = v$G35_9928_out0 && v$G36_3940_out0;
assign v$G40_8953_out0 = v$G35_9930_out0 && v$G36_3942_out0;
assign v$G40_8954_out0 = v$G35_9931_out0 && v$G36_3943_out0;
assign v$Q_9535_out0 = v$G4_7634_out0;
assign v$Q_9546_out0 = v$G4_7639_out0;
assign v$A3XNORB3_10076_out0 = v$G8_2443_out0;
assign v$A3XNORB3_10077_out0 = v$G8_2444_out0;
assign v$A3XNORB3_10079_out0 = v$G8_2446_out0;
assign v$A3XNORB3_10080_out0 = v$G8_2447_out0;
assign v$A3XNORB3_10088_out0 = v$G8_2455_out0;
assign v$A3XNORB3_10089_out0 = v$G8_2456_out0;
assign v$A3XNORB3_10091_out0 = v$G8_2458_out0;
assign v$A3XNORB3_10092_out0 = v$G8_2459_out0;
assign v$G11_10910_out0 = v$A2_5568_out0 && v$G12_11550_out0;
assign v$G11_10911_out0 = v$A2_5569_out0 && v$G12_11551_out0;
assign v$G11_10913_out0 = v$A2_5571_out0 && v$G12_11553_out0;
assign v$G11_10914_out0 = v$A2_5572_out0 && v$G12_11554_out0;
assign v$G11_10922_out0 = v$A2_5580_out0 && v$G12_11562_out0;
assign v$G11_10923_out0 = v$A2_5581_out0 && v$G12_11563_out0;
assign v$G11_10925_out0 = v$A2_5583_out0 && v$G12_11565_out0;
assign v$G11_10926_out0 = v$A2_5584_out0 && v$G12_11566_out0;
assign v$A1XNORB1_11229_out0 = v$G16_11915_out0;
assign v$A1XNORB1_11230_out0 = v$G16_11916_out0;
assign v$A1XNORB1_11232_out0 = v$G16_11918_out0;
assign v$A1XNORB1_11233_out0 = v$G16_11919_out0;
assign v$A1XNORB1_11241_out0 = v$G16_11927_out0;
assign v$A1XNORB1_11242_out0 = v$G16_11928_out0;
assign v$A1XNORB1_11244_out0 = v$G16_11930_out0;
assign v$A1XNORB1_11245_out0 = v$G16_11931_out0;
assign v$SAME_13355_out0 = v$G41_7159_out0;
assign v$SAME_13359_out0 = v$G41_7162_out0;
assign v$SAME_13364_out0 = v$G1_6390_out0;
assign v$SAME_13371_out0 = v$G41_7171_out0;
assign v$SAME_13375_out0 = v$G41_7174_out0;
assign v$SAME_13380_out0 = v$G1_6394_out0;
assign v$OUT_2634_out0 = v$G29_6860_out0;
assign v$OUT_2650_out0 = v$G29_6862_out0;
assign v$G13_3058_out0 = v$A3XNORB3_10076_out0 && v$G11_10910_out0;
assign v$G13_3059_out0 = v$A3XNORB3_10077_out0 && v$G11_10911_out0;
assign v$G13_3061_out0 = v$A3XNORB3_10079_out0 && v$G11_10913_out0;
assign v$G13_3062_out0 = v$A3XNORB3_10080_out0 && v$G11_10914_out0;
assign v$G13_3070_out0 = v$A3XNORB3_10088_out0 && v$G11_10922_out0;
assign v$G13_3071_out0 = v$A3XNORB3_10089_out0 && v$G11_10923_out0;
assign v$G13_3073_out0 = v$A3XNORB3_10091_out0 && v$G11_10925_out0;
assign v$G13_3074_out0 = v$A3XNORB3_10092_out0 && v$G11_10926_out0;
assign v$A3$COMP$B3_3342_out0 = v$G5_4708_out0;
assign v$A3$COMP$B3_3343_out0 = v$G5_4709_out0;
assign v$A3$COMP$B3_3345_out0 = v$G5_4711_out0;
assign v$A3$COMP$B3_3346_out0 = v$G5_4712_out0;
assign v$A3$COMP$B3_3354_out0 = v$G5_4720_out0;
assign v$A3$COMP$B3_3355_out0 = v$G5_4721_out0;
assign v$A3$COMP$B3_3357_out0 = v$G5_4723_out0;
assign v$A3$COMP$B3_3358_out0 = v$G5_4724_out0;
assign v$G3_6059_out0 = v$HIGHER$SAME_10331_out0 && v$LOWER$OUT_2902_out0;
assign v$G3_6063_out0 = v$HIGHER$SAME_10335_out0 && v$LOWER$OUT_2906_out0;
assign v$DIFF_6326_out0 = v$A1_3809_out0;
assign v$DIFF_6330_out0 = v$A1_3813_out0;
assign v$HIGHER$SAME_6366_out0 = v$SAME_13355_out0;
assign v$HIGHER$SAME_6367_out0 = v$SAME_13359_out0;
assign v$HIGHER$SAME_6368_out0 = v$SAME_13371_out0;
assign v$HIGHER$SAME_6369_out0 = v$SAME_13375_out0;
assign v$G41_7160_out0 = v$G38_4893_out0 && v$G40_8938_out0;
assign v$G41_7161_out0 = v$G38_4894_out0 && v$G40_8939_out0;
assign v$G41_7163_out0 = v$G38_4896_out0 && v$G40_8941_out0;
assign v$G41_7164_out0 = v$G38_4897_out0 && v$G40_8942_out0;
assign v$G41_7172_out0 = v$G38_4905_out0 && v$G40_8950_out0;
assign v$G41_7173_out0 = v$G38_4906_out0 && v$G40_8951_out0;
assign v$G41_7175_out0 = v$G38_4908_out0 && v$G40_8953_out0;
assign v$G41_7176_out0 = v$G38_4909_out0 && v$G40_8954_out0;
assign v$_7610_out0 = { v$_10004_out0,v$MUX6_1605_out0 };
assign v$_7614_out0 = { v$_10008_out0,v$MUX6_1606_out0 };
assign v$A1$COMP$B1_8130_out0 = v$G18_3369_out0;
assign v$A1$COMP$B1_8133_out0 = v$G18_3372_out0;
assign v$A1$COMP$B1_8142_out0 = v$G18_3381_out0;
assign v$A1$COMP$B1_8145_out0 = v$G18_3384_out0;
assign v$G28_8642_out0 = v$A1XNORB1_11229_out0 && v$G25_7207_out0;
assign v$G28_8643_out0 = v$A1XNORB1_11230_out0 && v$G25_7208_out0;
assign v$G28_8645_out0 = v$A1XNORB1_11232_out0 && v$G25_7210_out0;
assign v$G28_8646_out0 = v$A1XNORB1_11233_out0 && v$G25_7211_out0;
assign v$G28_8654_out0 = v$A1XNORB1_11241_out0 && v$G25_7219_out0;
assign v$G28_8655_out0 = v$A1XNORB1_11242_out0 && v$G25_7220_out0;
assign v$G28_8657_out0 = v$A1XNORB1_11244_out0 && v$G25_7222_out0;
assign v$G28_8658_out0 = v$A1XNORB1_11245_out0 && v$G25_7223_out0;
assign v$G22_8905_out0 = v$A2XNORB2_3129_out0 && v$G20_6623_out0;
assign v$G22_8906_out0 = v$A2XNORB2_3130_out0 && v$G20_6624_out0;
assign v$G22_8908_out0 = v$A2XNORB2_3132_out0 && v$G20_6626_out0;
assign v$G22_8909_out0 = v$A2XNORB2_3133_out0 && v$G20_6627_out0;
assign v$G22_8917_out0 = v$A2XNORB2_3141_out0 && v$G20_6635_out0;
assign v$G22_8918_out0 = v$A2XNORB2_3142_out0 && v$G20_6636_out0;
assign v$G22_8920_out0 = v$A2XNORB2_3144_out0 && v$G20_6638_out0;
assign v$G22_8921_out0 = v$A2XNORB2_3145_out0 && v$G20_6639_out0;
assign v$Q_9536_out0 = v$G4_7635_out0;
assign v$Q_9537_out0 = v$G4_7636_out0;
assign v$Q_9538_out0 = v$G4_7637_out0;
assign v$Q_9547_out0 = v$G4_7640_out0;
assign v$Q_9548_out0 = v$G4_7641_out0;
assign v$Q_9549_out0 = v$G4_7642_out0;
assign v$NOT$USED1_9760_out0 = v$A1_3809_out1;
assign v$NOT$USED1_9764_out0 = v$A1_3813_out1;
assign v$TXFlag_10569_out0 = v$TXFlag_5261_out0;
assign v$TXFlag_10570_out0 = v$TXFlag_5262_out0;
assign v$G31_10797_out0 = v$A2$COMP$B2_1125_out0 || v$G32_331_out0;
assign v$G31_10798_out0 = v$A2$COMP$B2_1126_out0 || v$G32_332_out0;
assign v$G31_10809_out0 = v$A2$COMP$B2_1137_out0 || v$G32_343_out0;
assign v$G31_10810_out0 = v$A2$COMP$B2_1138_out0 || v$G32_344_out0;
assign v$G24_10950_out0 = v$A3XNORB3_10075_out0 && v$G27_3188_out0;
assign v$G24_10953_out0 = v$A3XNORB3_10078_out0 && v$G27_3191_out0;
assign v$G24_10962_out0 = v$A3XNORB3_10087_out0 && v$G27_3200_out0;
assign v$G24_10965_out0 = v$A3XNORB3_10090_out0 && v$G27_3203_out0;
assign v$RXflag_11059_out0 = v$Q_9535_out0;
assign v$RXflag_11060_out0 = v$Q_9546_out0;
assign v$G6_11846_out0 = ! v$IGNORE_5757_out0;
assign v$SAME_13067_out0 = v$SAME_13364_out0;
assign v$SAME_13071_out0 = v$SAME_13380_out0;
assign v$G30_958_out0 = v$A3$COMP$B3_3348_out0 || v$G31_10797_out0;
assign v$G30_959_out0 = v$A3$COMP$B3_3349_out0 || v$G31_10798_out0;
assign v$G30_970_out0 = v$A3$COMP$B3_3360_out0 || v$G31_10809_out0;
assign v$G30_971_out0 = v$A3$COMP$B3_3361_out0 || v$G31_10810_out0;
assign v$A2$COMP$B2_1119_out0 = v$G13_3058_out0;
assign v$A2$COMP$B2_1120_out0 = v$G13_3059_out0;
assign v$A2$COMP$B2_1122_out0 = v$G13_3061_out0;
assign v$A2$COMP$B2_1123_out0 = v$G13_3062_out0;
assign v$A2$COMP$B2_1131_out0 = v$G13_3070_out0;
assign v$A2$COMP$B2_1132_out0 = v$G13_3071_out0;
assign v$A2$COMP$B2_1134_out0 = v$G13_3073_out0;
assign v$A2$COMP$B2_1135_out0 = v$G13_3074_out0;
assign v$MUX14_1723_out0 = v$IS$32$BIT_7152_out0 ? v$SAME_13067_out0 : v$SAME_13066_out0;
assign v$MUX14_1724_out0 = v$IS$32$BIT_7153_out0 ? v$SAME_13071_out0 : v$SAME_13070_out0;
assign v$MUX3_2099_out0 = v$OUT_2634_out0 ? v$A$EXP_238_out0 : v$B$EXP_11736_out0;
assign v$MUX3_2103_out0 = v$OUT_2650_out0 ? v$A$EXP_242_out0 : v$B$EXP_11740_out0;
assign v$Error_2475_out0 = v$Q_9538_out0;
assign v$Error_2476_out0 = v$Q_9549_out0;
assign v$TXoverflow_2807_out0 = v$Q_9536_out0;
assign v$TXoverflow_2808_out0 = v$Q_9547_out0;
assign v$G27_3189_out0 = v$A2XNORB2_3129_out0 && v$G28_8642_out0;
assign v$G27_3190_out0 = v$A2XNORB2_3130_out0 && v$G28_8643_out0;
assign v$G27_3192_out0 = v$A2XNORB2_3132_out0 && v$G28_8645_out0;
assign v$G27_3193_out0 = v$A2XNORB2_3133_out0 && v$G28_8646_out0;
assign v$G27_3201_out0 = v$A2XNORB2_3141_out0 && v$G28_8654_out0;
assign v$G27_3202_out0 = v$A2XNORB2_3142_out0 && v$G28_8655_out0;
assign v$G27_3204_out0 = v$A2XNORB2_3144_out0 && v$G28_8657_out0;
assign v$G27_3205_out0 = v$A2XNORB2_3145_out0 && v$G28_8658_out0;
assign v$G18_3370_out0 = v$A3XNORB3_10076_out0 && v$G22_8905_out0;
assign v$G18_3371_out0 = v$A3XNORB3_10077_out0 && v$G22_8906_out0;
assign v$G18_3373_out0 = v$A3XNORB3_10079_out0 && v$G22_8908_out0;
assign v$G18_3374_out0 = v$A3XNORB3_10080_out0 && v$G22_8909_out0;
assign v$G18_3382_out0 = v$A3XNORB3_10088_out0 && v$G22_8917_out0;
assign v$G18_3383_out0 = v$A3XNORB3_10089_out0 && v$G22_8918_out0;
assign v$G18_3385_out0 = v$A3XNORB3_10091_out0 && v$G22_8920_out0;
assign v$G18_3386_out0 = v$A3XNORB3_10092_out0 && v$G22_8921_out0;
assign v$MUX1_4669_out0 = v$G4_2748_out0 ? v$_7610_out0 : v$MUX2_7824_out0;
assign v$MUX1_4673_out0 = v$G4_2752_out0 ? v$_7614_out0 : v$MUX2_7828_out0;
assign v$A0$COMP$B0_5495_out0 = v$G24_10950_out0;
assign v$A0$COMP$B0_5498_out0 = v$G24_10953_out0;
assign v$A0$COMP$B0_5507_out0 = v$G24_10962_out0;
assign v$A0$COMP$B0_5510_out0 = v$G24_10965_out0;
assign v$RXoverflow_6516_out0 = v$Q_9537_out0;
assign v$RXoverflow_6517_out0 = v$Q_9548_out0;
assign v$RXFLAG_7909_out0 = v$RXflag_11059_out0;
assign v$RXFLAG_7910_out0 = v$RXflag_11060_out0;
assign v$G2_8548_out0 = v$HIGHER$OUT_2537_out0 || v$G3_6059_out0;
assign v$G2_8552_out0 = v$HIGHER$OUT_2541_out0 || v$G3_6063_out0;
assign v$OUT_9288_out0 = v$OUT_2634_out0;
assign v$OUT_9292_out0 = v$OUT_2650_out0;
assign v$TXFLAG_10050_out0 = v$TXFlag_10569_out0;
assign v$TXFLAG_10051_out0 = v$TXFlag_10570_out0;
assign v$_12214_out0 = { v$DIFF_6326_out0,v$C2_8899_out0 };
assign v$_12215_out0 = { v$DIFF_6330_out0,v$C2_8900_out0 };
assign v$G7_12491_out0 = v$G5_1570_out0 && v$G6_11846_out0;
assign v$MUX1_12701_out0 = v$OUT_2634_out0 ? v$B$EXP_11736_out0 : v$A$EXP_238_out0;
assign v$MUX1_12705_out0 = v$OUT_2650_out0 ? v$B$EXP_11740_out0 : v$A$EXP_242_out0;
assign v$SAME_13357_out0 = v$G41_7160_out0;
assign v$SAME_13358_out0 = v$G41_7161_out0;
assign v$SAME_13361_out0 = v$G41_7163_out0;
assign v$SAME_13362_out0 = v$G41_7164_out0;
assign v$SAME_13373_out0 = v$G41_7172_out0;
assign v$SAME_13374_out0 = v$G41_7173_out0;
assign v$SAME_13377_out0 = v$G41_7175_out0;
assign v$SAME_13378_out0 = v$G41_7176_out0;
assign v$G32_324_out0 = v$A1$COMP$B1_8130_out0 || v$A0$COMP$B0_5495_out0;
assign v$G32_327_out0 = v$A1$COMP$B1_8133_out0 || v$A0$COMP$B0_5498_out0;
assign v$G32_336_out0 = v$A1$COMP$B1_8142_out0 || v$A0$COMP$B0_5507_out0;
assign v$G32_339_out0 = v$A1$COMP$B1_8145_out0 || v$A0$COMP$B0_5510_out0;
assign v$EXP$SAME_408_out0 = v$MUX14_1723_out0;
assign v$EXP$SAME_409_out0 = v$MUX14_1724_out0;
assign v$MUX3_1100_out0 = v$G8_1038_out0 ? v$_8879_out0 : v$MUX1_4669_out0;
assign v$MUX3_1104_out0 = v$G8_1042_out0 ? v$_8883_out0 : v$MUX1_4673_out0;
assign v$TXFLAG_2586_out0 = v$TXFLAG_10050_out0;
assign v$TXFLAG_2587_out0 = v$TXFLAG_10051_out0;
assign v$OUT_2623_out0 = v$G2_8548_out0;
assign v$OUT_2636_out0 = v$G30_958_out0;
assign v$OUT_2637_out0 = v$G30_959_out0;
assign v$OUT_2639_out0 = v$G2_8552_out0;
assign v$OUT_2652_out0 = v$G30_970_out0;
assign v$OUT_2653_out0 = v$G30_971_out0;
assign v$XOR1_5130_out0 = v$C1_9149_out0 ^ v$MUX1_12701_out0;
assign v$XOR1_5134_out0 = v$C1_9153_out0 ^ v$MUX1_12705_out0;
assign v$_6649_out0 = { v$RXoverflow_6516_out0,v$Error_2475_out0 };
assign v$_6650_out0 = { v$RXoverflow_6517_out0,v$Error_2476_out0 };
assign v$LOWER$SAME_6758_out0 = v$SAME_13358_out0;
assign v$LOWER$SAME_6759_out0 = v$SAME_13362_out0;
assign v$LOWER$SAME_6762_out0 = v$SAME_13374_out0;
assign v$LOWER$SAME_6763_out0 = v$SAME_13378_out0;
assign v$A1$COMP$B1_8131_out0 = v$G18_3370_out0;
assign v$A1$COMP$B1_8132_out0 = v$G18_3371_out0;
assign v$A1$COMP$B1_8134_out0 = v$G18_3373_out0;
assign v$A1$COMP$B1_8135_out0 = v$G18_3374_out0;
assign v$A1$COMP$B1_8143_out0 = v$G18_3382_out0;
assign v$A1$COMP$B1_8144_out0 = v$G18_3383_out0;
assign v$A1$COMP$B1_8146_out0 = v$G18_3385_out0;
assign v$A1$COMP$B1_8147_out0 = v$G18_3386_out0;
assign v$RXFLAG_10319_out0 = v$RXFLAG_7909_out0;
assign v$RXFLAG_10320_out0 = v$RXFLAG_7910_out0;
assign v$HIGHER$SAME_10332_out0 = v$SAME_13357_out0;
assign v$HIGHER$SAME_10333_out0 = v$SAME_13361_out0;
assign v$HIGHER$SAME_10336_out0 = v$SAME_13373_out0;
assign v$HIGHER$SAME_10337_out0 = v$SAME_13377_out0;
assign v$_10615_out0 = { v$TXFlag_5261_out0,v$TXoverflow_2807_out0 };
assign v$_10616_out0 = { v$TXFlag_5262_out0,v$TXoverflow_2808_out0 };
assign v$G24_10951_out0 = v$A3XNORB3_10076_out0 && v$G27_3189_out0;
assign v$G24_10952_out0 = v$A3XNORB3_10077_out0 && v$G27_3190_out0;
assign v$G24_10954_out0 = v$A3XNORB3_10079_out0 && v$G27_3192_out0;
assign v$G24_10955_out0 = v$A3XNORB3_10080_out0 && v$G27_3193_out0;
assign v$G24_10963_out0 = v$A3XNORB3_10088_out0 && v$G27_3201_out0;
assign v$G24_10964_out0 = v$A3XNORB3_10089_out0 && v$G27_3202_out0;
assign v$G24_10966_out0 = v$A3XNORB3_10091_out0 && v$G27_3204_out0;
assign v$G24_10967_out0 = v$A3XNORB3_10092_out0 && v$G27_3205_out0;
assign v$RAMWEN_12732_out0 = v$G7_12491_out0;
assign v$F_1111_out0 = v$TXFLAG_2586_out0;
assign v$F_1112_out0 = v$TXFLAG_2587_out0;
assign v$OUT_1901_out0 = v$MUX3_1100_out0;
assign v$OUT_1905_out0 = v$MUX3_1104_out0;
assign v$MUX3_2098_out0 = v$OUT_2623_out0 ? v$A$EXP_237_out0 : v$B$EXP_11735_out0;
assign v$MUX3_2102_out0 = v$OUT_2639_out0 ? v$A$EXP_241_out0 : v$B$EXP_11739_out0;
assign v$HIGHER$OUT_2540_out0 = v$OUT_2636_out0;
assign v$HIGHER$OUT_2544_out0 = v$OUT_2652_out0;
assign v$LOWER$OUT_2905_out0 = v$OUT_2637_out0;
assign v$LOWER$OUT_2909_out0 = v$OUT_2653_out0;
assign {v$A1_3811_out1,v$A1_3811_out0 } = v$MUX3_2099_out0 + v$XOR1_5130_out0 + v$CIN_12954_out0;
assign {v$A1_3815_out1,v$A1_3815_out0 } = v$MUX3_2103_out0 + v$XOR1_5134_out0 + v$CIN_12958_out0;
assign v$A0$COMP$B0_5496_out0 = v$G24_10951_out0;
assign v$A0$COMP$B0_5497_out0 = v$G24_10952_out0;
assign v$A0$COMP$B0_5499_out0 = v$G24_10954_out0;
assign v$A0$COMP$B0_5500_out0 = v$G24_10955_out0;
assign v$A0$COMP$B0_5508_out0 = v$G24_10963_out0;
assign v$A0$COMP$B0_5509_out0 = v$G24_10964_out0;
assign v$A0$COMP$B0_5511_out0 = v$G24_10966_out0;
assign v$A0$COMP$B0_5512_out0 = v$G24_10967_out0;
assign v$G1_6388_out0 = v$LOWER$SAME_6758_out0 && v$HIGHER$SAME_10332_out0;
assign v$G1_6389_out0 = v$LOWER$SAME_6759_out0 && v$HIGHER$SAME_10333_out0;
assign v$G1_6392_out0 = v$LOWER$SAME_6762_out0 && v$HIGHER$SAME_10336_out0;
assign v$G1_6393_out0 = v$LOWER$SAME_6763_out0 && v$HIGHER$SAME_10337_out0;
assign v$OUT_9287_out0 = v$OUT_2623_out0;
assign v$OUT_9291_out0 = v$OUT_2639_out0;
assign v$G31_10790_out0 = v$A2$COMP$B2_1118_out0 || v$G32_324_out0;
assign v$G31_10793_out0 = v$A2$COMP$B2_1121_out0 || v$G32_327_out0;
assign v$G31_10802_out0 = v$A2$COMP$B2_1130_out0 || v$G32_336_out0;
assign v$G31_10805_out0 = v$A2$COMP$B2_1133_out0 || v$G32_339_out0;
assign v$MUX1_12700_out0 = v$OUT_2623_out0 ? v$B$EXP_11735_out0 : v$A$EXP_237_out0;
assign v$MUX1_12704_out0 = v$OUT_2639_out0 ? v$B$EXP_11739_out0 : v$A$EXP_241_out0;
assign v$_13197_out0 = { v$RXflag_11059_out0,v$_6649_out0 };
assign v$_13198_out0 = { v$RXflag_11060_out0,v$_6650_out0 };
assign v$G32_325_out0 = v$A1$COMP$B1_8131_out0 || v$A0$COMP$B0_5496_out0;
assign v$G32_326_out0 = v$A1$COMP$B1_8132_out0 || v$A0$COMP$B0_5497_out0;
assign v$G32_328_out0 = v$A1$COMP$B1_8134_out0 || v$A0$COMP$B0_5499_out0;
assign v$G32_329_out0 = v$A1$COMP$B1_8135_out0 || v$A0$COMP$B0_5500_out0;
assign v$G32_337_out0 = v$A1$COMP$B1_8143_out0 || v$A0$COMP$B0_5508_out0;
assign v$G32_338_out0 = v$A1$COMP$B1_8144_out0 || v$A0$COMP$B0_5509_out0;
assign v$G32_340_out0 = v$A1$COMP$B1_8146_out0 || v$A0$COMP$B0_5511_out0;
assign v$G32_341_out0 = v$A1$COMP$B1_8147_out0 || v$A0$COMP$B0_5512_out0;
assign v$G30_951_out0 = v$A3$COMP$B3_3341_out0 || v$G31_10790_out0;
assign v$G30_954_out0 = v$A3$COMP$B3_3344_out0 || v$G31_10793_out0;
assign v$G30_963_out0 = v$A3$COMP$B3_3353_out0 || v$G31_10802_out0;
assign v$G30_966_out0 = v$A3$COMP$B3_3356_out0 || v$G31_10805_out0;
assign v$G51_2159_out0 = v$NQ1_7276_out0 && v$F_1111_out0;
assign v$G51_2160_out0 = v$NQ1_7277_out0 && v$F_1112_out0;
assign v$G28_2473_out0 = ! v$F_1111_out0;
assign v$G28_2474_out0 = ! v$F_1112_out0;
assign v$IN_3019_out0 = v$OUT_1901_out0;
assign v$IN_3023_out0 = v$OUT_1905_out0;
assign v$_4353_out0 = { v$_10615_out0,v$_13197_out0 };
assign v$_4354_out0 = { v$_10616_out0,v$_13198_out0 };
assign v$XOR1_5129_out0 = v$C1_9148_out0 ^ v$MUX1_12700_out0;
assign v$XOR1_5133_out0 = v$C1_9152_out0 ^ v$MUX1_12704_out0;
assign v$G3_6062_out0 = v$HIGHER$SAME_10334_out0 && v$LOWER$OUT_2905_out0;
assign v$G3_6066_out0 = v$HIGHER$SAME_10338_out0 && v$LOWER$OUT_2909_out0;
assign v$DIFF_6328_out0 = v$A1_3811_out0;
assign v$DIFF_6332_out0 = v$A1_3815_out0;
assign v$NOT$USED1_9762_out0 = v$A1_3811_out1;
assign v$NOT$USED1_9766_out0 = v$A1_3815_out1;
assign v$MUX5_10781_out0 = v$IS$32$BITS_527_out0 ? v$OUT_9287_out0 : v$OUT_9286_out0;
assign v$MUX5_10782_out0 = v$IS$32$BITS_528_out0 ? v$OUT_9291_out0 : v$OUT_9290_out0;
assign v$SAME_13356_out0 = v$G1_6388_out0;
assign v$SAME_13360_out0 = v$G1_6389_out0;
assign v$SAME_13372_out0 = v$G1_6392_out0;
assign v$SAME_13376_out0 = v$G1_6393_out0;
assign v$LOWER$SAME_2501_out0 = v$SAME_13356_out0;
assign v$LOWER$SAME_2502_out0 = v$SAME_13360_out0;
assign v$LOWER$SAME_2503_out0 = v$SAME_13372_out0;
assign v$LOWER$SAME_2504_out0 = v$SAME_13376_out0;
assign v$OUT_2626_out0 = v$G30_951_out0;
assign v$OUT_2630_out0 = v$G30_954_out0;
assign v$OUT_2642_out0 = v$G30_963_out0;
assign v$OUT_2646_out0 = v$G30_966_out0;
assign {v$A1_3810_out1,v$A1_3810_out0 } = v$MUX3_2098_out0 + v$XOR1_5129_out0 + v$CIN_12953_out0;
assign {v$A1_3814_out1,v$A1_3814_out0 } = v$MUX3_2102_out0 + v$XOR1_5133_out0 + v$CIN_12957_out0;
assign v$_5148_out0 = { v$DIFF_6328_out0,v$C4_4630_out0 };
assign v$_5149_out0 = { v$DIFF_6332_out0,v$C4_4631_out0 };
assign v$A$EXP$LARGER_6437_out0 = v$MUX5_10781_out0;
assign v$A$EXP$LARGER_6438_out0 = v$MUX5_10782_out0;
assign v$IN_6535_out0 = v$IN_3019_out0;
assign v$IN_6539_out0 = v$IN_3023_out0;
assign v$G49_7290_out0 = v$G50_12147_out0 || v$G51_2159_out0;
assign v$G49_7291_out0 = v$G50_12148_out0 || v$G51_2160_out0;
assign v$G2_8551_out0 = v$HIGHER$OUT_2540_out0 || v$G3_6062_out0;
assign v$G2_8555_out0 = v$HIGHER$OUT_2544_out0 || v$G3_6066_out0;
assign v$NF_9947_out0 = v$G28_2473_out0;
assign v$NF_9948_out0 = v$G28_2474_out0;
assign v$G31_10791_out0 = v$A2$COMP$B2_1119_out0 || v$G32_325_out0;
assign v$G31_10792_out0 = v$A2$COMP$B2_1120_out0 || v$G32_326_out0;
assign v$G31_10794_out0 = v$A2$COMP$B2_1122_out0 || v$G32_328_out0;
assign v$G31_10795_out0 = v$A2$COMP$B2_1123_out0 || v$G32_329_out0;
assign v$G31_10803_out0 = v$A2$COMP$B2_1131_out0 || v$G32_337_out0;
assign v$G31_10804_out0 = v$A2$COMP$B2_1132_out0 || v$G32_338_out0;
assign v$G31_10806_out0 = v$A2$COMP$B2_1134_out0 || v$G32_340_out0;
assign v$G31_10807_out0 = v$A2$COMP$B2_1135_out0 || v$G32_341_out0;
assign v$_11334_out0 = { v$_4353_out0,v$C1_11890_out0 };
assign v$_11335_out0 = { v$_4354_out0,v$C1_11891_out0 };
assign v$G30_952_out0 = v$A3$COMP$B3_3342_out0 || v$G31_10791_out0;
assign v$G30_953_out0 = v$A3$COMP$B3_3343_out0 || v$G31_10792_out0;
assign v$G30_955_out0 = v$A3$COMP$B3_3345_out0 || v$G31_10794_out0;
assign v$G30_956_out0 = v$A3$COMP$B3_3346_out0 || v$G31_10795_out0;
assign v$G30_964_out0 = v$A3$COMP$B3_3354_out0 || v$G31_10803_out0;
assign v$G30_965_out0 = v$A3$COMP$B3_3355_out0 || v$G31_10804_out0;
assign v$G30_967_out0 = v$A3$COMP$B3_3357_out0 || v$G31_10806_out0;
assign v$G30_968_out0 = v$A3$COMP$B3_3358_out0 || v$G31_10807_out0;
assign v$G2_1044_out0 = v$EXP$SAME_11626_out0 || v$A$EXP$LARGER_6437_out0;
assign v$G2_1045_out0 = v$EXP$SAME_11627_out0 || v$A$EXP$LARGER_6438_out0;
assign v$Status_2499_out0 = v$_11334_out0;
assign v$Status_2500_out0 = v$_11335_out0;
assign v$OUT_2635_out0 = v$G2_8551_out0;
assign v$OUT_2651_out0 = v$G2_8555_out0;
assign v$_3212_out0 = v$IN_6535_out0[7:0];
assign v$_3216_out0 = v$IN_6539_out0[7:0];
assign v$_5052_out0 = v$IN_6535_out0[15:15];
assign v$_5053_out0 = v$IN_6539_out0[15:15];
assign v$HIGHER$OUT_5318_out0 = v$OUT_2626_out0;
assign v$HIGHER$OUT_5319_out0 = v$OUT_2630_out0;
assign v$HIGHER$OUT_5320_out0 = v$OUT_2642_out0;
assign v$HIGHER$OUT_5321_out0 = v$OUT_2646_out0;
assign v$DIFF_6327_out0 = v$A1_3810_out0;
assign v$DIFF_6331_out0 = v$A1_3814_out0;
assign v$_8854_out0 = v$IN_6535_out0[7:0];
assign v$_8857_out0 = v$IN_6539_out0[7:0];
assign v$_9482_out0 = v$IN_6535_out0[7:0];
assign v$_9483_out0 = v$IN_6539_out0[7:0];
assign v$NOT$USED1_9761_out0 = v$A1_3810_out1;
assign v$NOT$USED1_9765_out0 = v$A1_3814_out1;
assign v$_9979_out0 = v$IN_6535_out0[15:8];
assign v$_9983_out0 = v$IN_6539_out0[15:8];
assign v$_10005_out0 = v$IN_6535_out0[15:8];
assign v$_10009_out0 = v$IN_6539_out0[15:8];
assign v$IS$A$LARGER_10027_out0 = v$A$EXP$LARGER_6437_out0;
assign v$IS$A$LARGER_10028_out0 = v$A$EXP$LARGER_6438_out0;
assign v$G4_10637_out0 = v$EXP$SAME_11626_out0 || v$A$EXP$LARGER_6437_out0;
assign v$G4_10638_out0 = v$EXP$SAME_11627_out0 || v$A$EXP$LARGER_6438_out0;
assign v$_11797_out0 = v$IN_6535_out0[15:8];
assign v$_11801_out0 = v$IN_6539_out0[15:8];
assign v$G1_12250_out0 = v$LOWER$SAME_2501_out0 && v$HIGHER$SAME_6366_out0;
assign v$G1_12251_out0 = v$LOWER$SAME_2502_out0 && v$HIGHER$SAME_6367_out0;
assign v$G1_12252_out0 = v$LOWER$SAME_2503_out0 && v$HIGHER$SAME_6368_out0;
assign v$G1_12253_out0 = v$LOWER$SAME_2504_out0 && v$HIGHER$SAME_6369_out0;
assign v$G48_13173_out0 = v$NQ0_10890_out0 && v$G49_7290_out0;
assign v$G48_13174_out0 = v$NQ0_10891_out0 && v$G49_7291_out0;
assign v$_712_out0 = { v$C1_5481_out0,v$_3212_out0 };
assign v$_716_out0 = { v$C1_5485_out0,v$_3216_out0 };
assign v$MUX2_813_out0 = v$IS$A$LARGER_10027_out0 ? v$SEL4_1201_out0 : v$SEL3_7684_out0;
assign v$MUX2_814_out0 = v$IS$A$LARGER_10028_out0 ? v$SEL4_1202_out0 : v$SEL3_7685_out0;
assign v$MUX1_1084_out0 = v$IS$A$LARGER_10027_out0 ? v$SEL1_10991_out0 : v$SEL2_7265_out0;
assign v$MUX1_1085_out0 = v$IS$A$LARGER_10028_out0 ? v$SEL1_10992_out0 : v$SEL2_7266_out0;
assign v$MUX3_2100_out0 = v$OUT_2635_out0 ? v$A$EXP_239_out0 : v$B$EXP_11737_out0;
assign v$MUX3_2104_out0 = v$OUT_2651_out0 ? v$A$EXP_243_out0 : v$B$EXP_11741_out0;
assign v$OUT_2628_out0 = v$G30_952_out0;
assign v$OUT_2629_out0 = v$G30_953_out0;
assign v$OUT_2632_out0 = v$G30_955_out0;
assign v$OUT_2633_out0 = v$G30_956_out0;
assign v$OUT_2644_out0 = v$G30_964_out0;
assign v$OUT_2645_out0 = v$G30_965_out0;
assign v$OUT_2648_out0 = v$G30_967_out0;
assign v$OUT_2649_out0 = v$G30_968_out0;
assign v$MUX1_2758_out0 = v$G2_1044_out0 ? v$B_7913_out0 : v$A_11271_out0;
assign v$MUX1_2759_out0 = v$G2_1045_out0 ? v$B_7914_out0 : v$A_11272_out0;
assign v$MUX6_5444_out0 = v$IS$32$BITS_527_out0 ? v$DIFF_6327_out0 : v$_12214_out0;
assign v$MUX6_5445_out0 = v$IS$32$BITS_528_out0 ? v$DIFF_6331_out0 : v$_12215_out0;
assign v$STATUS_6055_out0 = v$Status_2499_out0;
assign v$STATUS_6056_out0 = v$Status_2500_out0;
assign v$SAME_6171_out0 = v$G1_12250_out0;
assign v$SAME_6172_out0 = v$G1_12251_out0;
assign v$SAME_6173_out0 = v$G1_12252_out0;
assign v$SAME_6174_out0 = v$G1_12253_out0;
assign v$_6444_out0 = { v$_11797_out0,v$LSBS_5438_out0 };
assign v$_6448_out0 = { v$_11801_out0,v$LSBS_5439_out0 };
assign v$_8880_out0 = { v$_9979_out0,v$_8854_out0 };
assign v$_8884_out0 = { v$_9983_out0,v$_8857_out0 };
assign v$MUX6_9251_out0 = v$S_12723_out0 ? v$_9482_out0 : v$C1_9014_out0;
assign v$MUX6_9252_out0 = v$S_12724_out0 ? v$_9483_out0 : v$C1_9015_out0;
assign v$OUT_9289_out0 = v$OUT_2635_out0;
assign v$OUT_9293_out0 = v$OUT_2651_out0;
assign v$MUX2_10495_out0 = v$G2_1044_out0 ? v$A_11271_out0 : v$B_7913_out0;
assign v$MUX2_10496_out0 = v$G2_1045_out0 ? v$A_11272_out0 : v$B_7914_out0;
assign v$MUX10_11878_out0 = v$G4_10637_out0 ? v$A_11271_out0 : v$B_7913_out0;
assign v$MUX10_11879_out0 = v$G4_10638_out0 ? v$A_11272_out0 : v$B_7914_out0;
assign v$G5_12662_out0 = v$G6_1891_out0 || v$G48_13173_out0;
assign v$G5_12663_out0 = v$G6_1892_out0 || v$G48_13174_out0;
assign v$MUX1_12702_out0 = v$OUT_2635_out0 ? v$B$EXP_11737_out0 : v$A$EXP_239_out0;
assign v$MUX1_12706_out0 = v$OUT_2651_out0 ? v$B$EXP_11741_out0 : v$A$EXP_243_out0;
assign v$MUX9_12717_out0 = v$G4_10637_out0 ? v$B_7913_out0 : v$A_11271_out0;
assign v$MUX9_12718_out0 = v$G4_10638_out0 ? v$B_7914_out0 : v$A_11272_out0;
assign v$_12735_out0 = { v$_5052_out0,v$_5052_out0 };
assign v$_12736_out0 = { v$_5053_out0,v$_5053_out0 };
assign v$SEL10_1771_out0 = v$MUX9_12717_out0[14:10];
assign v$SEL10_1772_out0 = v$MUX9_12718_out0[14:10];
assign v$SEL9_2481_out0 = v$MUX10_11878_out0[14:10];
assign v$SEL9_2482_out0 = v$MUX10_11879_out0[14:10];
assign v$HIGHER$OUT_2538_out0 = v$OUT_2628_out0;
assign v$HIGHER$OUT_2539_out0 = v$OUT_2632_out0;
assign v$HIGHER$OUT_2542_out0 = v$OUT_2644_out0;
assign v$HIGHER$OUT_2543_out0 = v$OUT_2648_out0;
assign v$LOWER$OUT_2903_out0 = v$OUT_2629_out0;
assign v$LOWER$OUT_2904_out0 = v$OUT_2633_out0;
assign v$LOWER$OUT_2907_out0 = v$OUT_2645_out0;
assign v$LOWER$OUT_2908_out0 = v$OUT_2649_out0;
assign v$MUX2_3252_out0 = v$IS$32$BIT_7152_out0 ? v$OUT_9289_out0 : v$OUT_9288_out0;
assign v$MUX2_3253_out0 = v$IS$32$BIT_7153_out0 ? v$OUT_9293_out0 : v$OUT_9292_out0;
assign v$XOR1_5131_out0 = v$C1_9150_out0 ^ v$MUX1_12702_out0;
assign v$XOR1_5135_out0 = v$C1_9154_out0 ^ v$MUX1_12706_out0;
assign v$MUX1_5175_out0 = v$G47_753_out0 ? v$C1_703_out0 : v$G5_12662_out0;
assign v$MUX1_5176_out0 = v$G47_754_out0 ? v$C1_704_out0 : v$G5_12663_out0;
assign v$SAME$H_6167_out0 = v$SAME_6171_out0;
assign v$SAME$H_6168_out0 = v$SAME_6173_out0;
assign v$_7269_out0 = { v$MUX2_813_out0,v$C2_2336_out0 };
assign v$_7270_out0 = { v$MUX2_814_out0,v$C2_2337_out0 };
assign v$SEL4_7972_out0 = v$MUX2_10495_out0[14:7];
assign v$SEL4_7973_out0 = v$MUX2_10496_out0[14:7];
assign v$EXP$DIFF_8111_out0 = v$MUX6_5444_out0;
assign v$EXP$DIFF_8112_out0 = v$MUX6_5445_out0;
assign v$_9480_out0 = { v$MUX1_1084_out0,v$C1_3012_out0 };
assign v$_9481_out0 = { v$MUX1_1085_out0,v$C1_3013_out0 };
assign v$MUX4_11181_out0 = v$EN_12032_out0 ? v$_712_out0 : v$IN_6535_out0;
assign v$MUX4_11185_out0 = v$EN_12036_out0 ? v$_716_out0 : v$IN_6539_out0;
assign v$SAME$L_11525_out0 = v$SAME_6172_out0;
assign v$SAME$L_11526_out0 = v$SAME_6174_out0;
assign v$_12218_out0 = { v$_12735_out0,v$_12735_out0 };
assign v$_12219_out0 = { v$_12736_out0,v$_12736_out0 };
assign v$MUX2_12550_out0 = v$FF2_6413_out0 ? v$STATUS_6055_out0 : v$RXBYTE_6584_out0;
assign v$MUX2_12551_out0 = v$FF2_6414_out0 ? v$STATUS_6056_out0 : v$RXBYTE_6585_out0;
assign v$SEL3_12613_out0 = v$MUX1_2758_out0[14:7];
assign v$SEL3_12614_out0 = v$MUX1_2759_out0[14:7];
assign v$SMALLER$EXP_1707_out0 = v$SEL10_1771_out0;
assign v$SMALLER$EXP_1708_out0 = v$SEL3_12613_out0;
assign v$SMALLER$EXP_1709_out0 = v$SEL10_1772_out0;
assign v$SMALLER$EXP_1710_out0 = v$SEL3_12614_out0;
assign {v$A1_3812_out1,v$A1_3812_out0 } = v$MUX3_2100_out0 + v$XOR1_5131_out0 + v$CIN_12955_out0;
assign {v$A1_3816_out1,v$A1_3816_out0 } = v$MUX3_2104_out0 + v$XOR1_5135_out0 + v$CIN_12959_out0;
assign v$_4688_out0 = { v$MUX2_12550_out0,v$C1_10160_out0 };
assign v$_4689_out0 = { v$MUX2_12551_out0,v$C1_10161_out0 };
assign v$G3_6060_out0 = v$HIGHER$SAME_10332_out0 && v$LOWER$OUT_2903_out0;
assign v$G3_6061_out0 = v$HIGHER$SAME_10333_out0 && v$LOWER$OUT_2904_out0;
assign v$G3_6064_out0 = v$HIGHER$SAME_10336_out0 && v$LOWER$OUT_2907_out0;
assign v$G3_6065_out0 = v$HIGHER$SAME_10337_out0 && v$LOWER$OUT_2908_out0;
assign v$LARGER$EXP_6839_out0 = v$SEL9_2481_out0;
assign v$LARGER$EXP_6840_out0 = v$SEL4_7972_out0;
assign v$LARGER$EXP_6841_out0 = v$SEL9_2482_out0;
assign v$LARGER$EXP_6842_out0 = v$SEL4_7973_out0;
assign v$MUX2_7825_out0 = v$G3_1510_out0 ? v$_6444_out0 : v$MUX4_11181_out0;
assign v$MUX2_7829_out0 = v$G3_1514_out0 ? v$_6448_out0 : v$MUX4_11185_out0;
assign v$IN_8774_out0 = v$_7269_out0;
assign v$IN_8778_out0 = v$_7270_out0;
assign v$_9705_out0 = { v$_12218_out0,v$_12218_out0 };
assign v$_9706_out0 = { v$_12219_out0,v$_12219_out0 };
assign v$EXP$DIFF_9717_out0 = v$EXP$DIFF_8111_out0;
assign v$EXP$DIFF_9718_out0 = v$EXP$DIFF_8112_out0;
assign v$SEL5_11341_out0 = v$_9480_out0[23:13];
assign v$SEL5_11342_out0 = v$_9481_out0[23:13];
assign v$Q0P_11821_out0 = v$MUX1_5175_out0;
assign v$Q0P_11822_out0 = v$MUX1_5176_out0;
assign v$DIFF_12292_out0 = v$EXP$DIFF_8111_out0;
assign v$DIFF_12293_out0 = v$EXP$DIFF_8111_out0;
assign v$DIFF_12294_out0 = v$EXP$DIFF_8112_out0;
assign v$DIFF_12295_out0 = v$EXP$DIFF_8112_out0;
assign v$A$EXP$LARGER_12968_out0 = v$MUX2_3252_out0;
assign v$A$EXP$LARGER_12969_out0 = v$MUX2_3253_out0;
assign v$G4_12987_out0 = v$SAME$L_11525_out0 && v$SAME$H_6167_out0;
assign v$G4_12988_out0 = v$SAME$L_11526_out0 && v$SAME$H_6168_out0;
assign v$MUX1_1139_out0 = v$FF1_7292_out0 ? v$_4688_out0 : v$RAMDOUT_11827_out0;
assign v$MUX1_1140_out0 = v$FF1_7293_out0 ? v$_4689_out0 : v$RAMDOUT_11828_out0;
assign v$IN_3523_out0 = v$IN_8774_out0;
assign v$IN_3555_out0 = v$IN_8778_out0;
assign v$SAME_4265_out0 = v$G4_12987_out0;
assign v$SAME_4266_out0 = v$G4_12988_out0;
assign v$DIFF_6329_out0 = v$A1_3812_out0;
assign v$DIFF_6333_out0 = v$A1_3816_out0;
assign v$_6744_out0 = { v$C4_1379_out0,v$SEL5_11341_out0 };
assign v$_6745_out0 = { v$C4_1380_out0,v$SEL5_11342_out0 };
assign v$G2_8549_out0 = v$HIGHER$OUT_2538_out0 || v$G3_6060_out0;
assign v$G2_8550_out0 = v$HIGHER$OUT_2539_out0 || v$G3_6061_out0;
assign v$G2_8553_out0 = v$HIGHER$OUT_2542_out0 || v$G3_6064_out0;
assign v$G2_8554_out0 = v$HIGHER$OUT_2543_out0 || v$G3_6065_out0;
assign v$MUX5_8784_out0 = v$FF1_5716_out0 ? v$LSBS_5438_out0 : v$_9705_out0;
assign v$MUX5_8785_out0 = v$FF1_5717_out0 ? v$LSBS_5439_out0 : v$_9706_out0;
assign v$N_9462_out0 = v$DIFF_12292_out0;
assign v$N_9463_out0 = v$DIFF_12293_out0;
assign v$N_9464_out0 = v$DIFF_12294_out0;
assign v$N_9465_out0 = v$DIFF_12295_out0;
assign v$NOT$USED1_9763_out0 = v$A1_3812_out1;
assign v$NOT$USED1_9767_out0 = v$A1_3816_out1;
assign v$_11300_out0 = { v$Q0P_11821_out0,v$Q1P_3774_out0 };
assign v$_11301_out0 = { v$Q0P_11822_out0,v$Q1P_3775_out0 };
assign v$EXP$DIFF_12503_out0 = v$EXP$DIFF_9717_out0;
assign v$EXP$DIFF_12504_out0 = v$EXP$DIFF_9718_out0;
assign v$MANTISA$SAME_1363_out0 = v$SAME_4265_out0;
assign v$MANTISA$SAME_1364_out0 = v$SAME_4266_out0;
assign v$MUX3_1862_out0 = v$IS$32$BITS_2837_out0 ? v$_9480_out0 : v$_6744_out0;
assign v$MUX3_1863_out0 = v$IS$32$BITS_2838_out0 ? v$_9481_out0 : v$_6745_out0;
assign v$RAMDOutOut_1911_out0 = v$MUX1_1139_out0;
assign v$RAMDOutOut_1912_out0 = v$MUX1_1140_out0;
assign v$IN_2566_out0 = v$IN_3523_out0;
assign v$IN_2576_out0 = v$IN_3555_out0;
assign v$OUT_2627_out0 = v$G2_8549_out0;
assign v$OUT_2631_out0 = v$G2_8550_out0;
assign v$OUT_2643_out0 = v$G2_8553_out0;
assign v$OUT_2647_out0 = v$G2_8554_out0;
assign v$SEL26_3242_out0 = v$N_9462_out0[7:5];
assign v$SEL26_3243_out0 = v$N_9463_out0[7:5];
assign v$SEL26_3244_out0 = v$N_9464_out0[7:5];
assign v$SEL26_3245_out0 = v$N_9465_out0[7:5];
assign v$SHIFT$AMOUNT_4980_out0 = v$EXP$DIFF_12503_out0;
assign v$SHIFT$AMOUNT_4984_out0 = v$EXP$DIFF_12504_out0;
assign v$_6427_out0 = { v$_11300_out0,v$_1571_out0 };
assign v$_6428_out0 = { v$_11301_out0,v$_1572_out0 };
assign v$MUX13_6905_out0 = v$IS$32$BIT_7152_out0 ? v$DIFF_6329_out0 : v$_5148_out0;
assign v$MUX13_6906_out0 = v$IS$32$BIT_7153_out0 ? v$DIFF_6333_out0 : v$_5149_out0;
assign v$_7611_out0 = { v$_10005_out0,v$MUX5_8784_out0 };
assign v$_7615_out0 = { v$_10009_out0,v$MUX5_8785_out0 };
assign v$SEL25_9020_out0 = v$N_9462_out0[4:0];
assign v$SEL25_9021_out0 = v$N_9463_out0[4:0];
assign v$SEL25_9022_out0 = v$N_9464_out0[4:0];
assign v$SEL25_9023_out0 = v$N_9465_out0[4:0];
assign v$SEL3_437_out0 = v$SHIFT$AMOUNT_4980_out0[2:2];
assign v$SEL3_441_out0 = v$SHIFT$AMOUNT_4984_out0[2:2];
assign v$SEL1_1191_out0 = v$SHIFT$AMOUNT_4980_out0[0:0];
assign v$SEL1_1195_out0 = v$SHIFT$AMOUNT_4984_out0[0:0];
assign v$OP1_2798_out0 = v$MUX3_1862_out0;
assign v$OP1_2799_out0 = v$MUX3_1863_out0;
assign v$SEL4_3330_out0 = v$SHIFT$AMOUNT_4980_out0[3:3];
assign v$SEL4_3334_out0 = v$SHIFT$AMOUNT_4984_out0[3:3];
assign v$SEL7_4357_out0 = v$SHIFT$AMOUNT_4980_out0[5:5];
assign v$SEL7_4361_out0 = v$SHIFT$AMOUNT_4984_out0[5:5];
assign v$LOWER$OUT_4434_out0 = v$OUT_2627_out0;
assign v$LOWER$OUT_4435_out0 = v$OUT_2631_out0;
assign v$LOWER$OUT_4436_out0 = v$OUT_2643_out0;
assign v$LOWER$OUT_4437_out0 = v$OUT_2647_out0;
assign v$MUX1_4670_out0 = v$G4_2749_out0 ? v$_7611_out0 : v$MUX2_7825_out0;
assign v$MUX1_4674_out0 = v$G4_2753_out0 ? v$_7615_out0 : v$MUX2_7829_out0;
assign v$SEL1_5936_out0 = v$IN_2566_out0[23:1];
assign v$SEL1_5968_out0 = v$IN_2576_out0[23:1];
assign v$SEL5_7988_out0 = v$SHIFT$AMOUNT_4980_out0[4:4];
assign v$SEL5_7992_out0 = v$SHIFT$AMOUNT_4984_out0[4:4];
assign v$DIFF_8303_out0 = v$MUX13_6905_out0;
assign v$DIFF_8304_out0 = v$MUX13_6906_out0;
assign v$SEL6_9304_out0 = v$SHIFT$AMOUNT_4980_out0[6:6];
assign v$SEL6_9308_out0 = v$SHIFT$AMOUNT_4984_out0[6:6];
assign v$SEL1_10680_out0 = v$IN_2566_out0[22:0];
assign v$SEL1_10712_out0 = v$IN_2576_out0[22:0];
assign v$N_11398_out0 = v$SEL25_9020_out0;
assign v$N_11399_out0 = v$SEL25_9021_out0;
assign v$N_11400_out0 = v$SEL25_9022_out0;
assign v$N_11401_out0 = v$SEL25_9023_out0;
assign v$SEL8_11646_out0 = v$SHIFT$AMOUNT_4980_out0[7:7];
assign v$SEL8_11650_out0 = v$SHIFT$AMOUNT_4984_out0[7:7];
assign v$NUPPER_12173_out0 = v$SEL26_3242_out0;
assign v$NUPPER_12174_out0 = v$SEL26_3243_out0;
assign v$NUPPER_12175_out0 = v$SEL26_3244_out0;
assign v$NUPPER_12176_out0 = v$SEL26_3245_out0;
assign v$UART$DOUT_12260_out0 = v$RAMDOutOut_1911_out0;
assign v$UART$DOUT_12261_out0 = v$RAMDOutOut_1912_out0;
assign v$SEL2_13056_out0 = v$SHIFT$AMOUNT_4980_out0[1:1];
assign v$SEL2_13060_out0 = v$SHIFT$AMOUNT_4984_out0[1:1];
assign v$DIFF_244_out0 = v$DIFF_8303_out0;
assign v$DIFF_245_out0 = v$DIFF_8304_out0;
assign v$EN_561_out0 = v$SEL5_7988_out0;
assign v$EN_562_out0 = v$SEL4_3330_out0;
assign v$EN_571_out0 = v$SEL5_7992_out0;
assign v$EN_572_out0 = v$SEL4_3334_out0;
assign v$EQ3_991_out0 = v$N_11398_out0 == 5'h2;
assign v$EQ3_992_out0 = v$N_11399_out0 == 5'h2;
assign v$EQ3_993_out0 = v$N_11400_out0 == 5'h2;
assign v$EQ3_994_out0 = v$N_11401_out0 == 5'h2;
assign v$MUX3_1101_out0 = v$G8_1039_out0 ? v$_8880_out0 : v$MUX1_4670_out0;
assign v$MUX3_1105_out0 = v$G8_1043_out0 ? v$_8884_out0 : v$MUX1_4674_out0;
assign v$EQ24_1445_out0 = v$N_11398_out0 == 5'h17;
assign v$EQ24_1446_out0 = v$N_11399_out0 == 5'h17;
assign v$EQ24_1447_out0 = v$N_11400_out0 == 5'h17;
assign v$EQ24_1448_out0 = v$N_11401_out0 == 5'h17;
assign v$EQ22_1599_out0 = v$N_11398_out0 == 5'h15;
assign v$EQ22_1600_out0 = v$N_11399_out0 == 5'h15;
assign v$EQ22_1601_out0 = v$N_11400_out0 == 5'h15;
assign v$EQ22_1602_out0 = v$N_11401_out0 == 5'h15;
assign v$EQ23_1913_out0 = v$N_11398_out0 == 5'h16;
assign v$EQ23_1914_out0 = v$N_11399_out0 == 5'h16;
assign v$EQ23_1915_out0 = v$N_11400_out0 == 5'h16;
assign v$EQ23_1916_out0 = v$N_11401_out0 == 5'h16;
assign v$EQ5_2013_out0 = v$N_11398_out0 == 5'h4;
assign v$EQ5_2014_out0 = v$N_11399_out0 == 5'h4;
assign v$EQ5_2015_out0 = v$N_11400_out0 == 5'h4;
assign v$EQ5_2016_out0 = v$N_11401_out0 == 5'h4;
assign v$EQ21_2017_out0 = v$N_11398_out0 == 5'h14;
assign v$EQ21_2018_out0 = v$N_11399_out0 == 5'h14;
assign v$EQ21_2019_out0 = v$N_11400_out0 == 5'h14;
assign v$EQ21_2020_out0 = v$N_11401_out0 == 5'h14;
assign v$EQ7_2788_out0 = v$N_11398_out0 == 5'h6;
assign v$EQ7_2789_out0 = v$N_11399_out0 == 5'h6;
assign v$EQ7_2790_out0 = v$N_11400_out0 == 5'h6;
assign v$EQ7_2791_out0 = v$N_11401_out0 == 5'h6;
assign v$_2922_out0 = { v$C2_98_out0,v$SEL1_10680_out0 };
assign v$_2954_out0 = { v$C2_130_out0,v$SEL1_10712_out0 };
assign v$EN_3165_out0 = v$SEL3_437_out0;
assign v$EN_3171_out0 = v$SEL3_441_out0;
assign v$EN_3585_out0 = v$SEL1_1191_out0;
assign v$EN_3595_out0 = v$SEL1_1195_out0;
assign v$EQ14_3647_out0 = v$N_11398_out0 == 5'hd;
assign v$EQ14_3648_out0 = v$N_11399_out0 == 5'hd;
assign v$EQ14_3649_out0 = v$N_11400_out0 == 5'hd;
assign v$EQ14_3650_out0 = v$N_11401_out0 == 5'hd;
assign v$A_3663_out0 = v$OP1_2798_out0;
assign v$A_3664_out0 = v$OP1_2799_out0;
assign v$EQ6_3671_out0 = v$N_11398_out0 == 5'h5;
assign v$EQ6_3672_out0 = v$N_11399_out0 == 5'h5;
assign v$EQ6_3673_out0 = v$N_11400_out0 == 5'h5;
assign v$EQ6_3674_out0 = v$N_11401_out0 == 5'h5;
assign v$EQ19_3689_out0 = v$N_11398_out0 == 5'h12;
assign v$EQ19_3690_out0 = v$N_11399_out0 == 5'h12;
assign v$EQ19_3691_out0 = v$N_11400_out0 == 5'h12;
assign v$EQ19_3692_out0 = v$N_11401_out0 == 5'h12;
assign v$EQ17_3906_out0 = v$N_11398_out0 == 5'h10;
assign v$EQ17_3907_out0 = v$N_11399_out0 == 5'h10;
assign v$EQ17_3908_out0 = v$N_11400_out0 == 5'h10;
assign v$EQ17_3909_out0 = v$N_11401_out0 == 5'h10;
assign v$EQ10_3914_out0 = v$N_11398_out0 == 5'h8;
assign v$EQ10_3915_out0 = v$N_11399_out0 == 5'h8;
assign v$EQ10_3916_out0 = v$N_11400_out0 == 5'h8;
assign v$EQ10_3917_out0 = v$N_11401_out0 == 5'h8;
assign v$EQ11_4157_out0 = v$N_11398_out0 == 5'ha;
assign v$EQ11_4158_out0 = v$N_11399_out0 == 5'ha;
assign v$EQ11_4159_out0 = v$N_11400_out0 == 5'ha;
assign v$EQ11_4160_out0 = v$N_11401_out0 == 5'ha;
assign v$SEL28_4925_out0 = v$NUPPER_12173_out0[1:1];
assign v$SEL28_4926_out0 = v$NUPPER_12174_out0[1:1];
assign v$SEL28_4927_out0 = v$NUPPER_12175_out0[1:1];
assign v$SEL28_4928_out0 = v$NUPPER_12176_out0[1:1];
assign v$EN_5389_out0 = v$SEL2_13056_out0;
assign v$EN_5395_out0 = v$SEL2_13060_out0;
assign v$RAMDOUT_5424_out0 = v$UART$DOUT_12260_out0;
assign v$RAMDOUT_5425_out0 = v$UART$DOUT_12261_out0;
assign v$EQ16_5760_out0 = v$N_11398_out0 == 5'hf;
assign v$EQ16_5761_out0 = v$N_11399_out0 == 5'hf;
assign v$EQ16_5762_out0 = v$N_11400_out0 == 5'hf;
assign v$EQ16_5763_out0 = v$N_11401_out0 == 5'hf;
assign v$_6229_out0 = { v$SEL1_5936_out0,v$C1_3965_out0 };
assign v$_6261_out0 = { v$SEL1_5968_out0,v$C1_3997_out0 };
assign v$EQ13_6491_out0 = v$N_11398_out0 == 5'hc;
assign v$EQ13_6492_out0 = v$N_11399_out0 == 5'hc;
assign v$EQ13_6493_out0 = v$N_11400_out0 == 5'hc;
assign v$EQ13_6494_out0 = v$N_11401_out0 == 5'hc;
assign v$EQ20_6666_out0 = v$N_11398_out0 == 5'h13;
assign v$EQ20_6667_out0 = v$N_11399_out0 == 5'h13;
assign v$EQ20_6668_out0 = v$N_11400_out0 == 5'h13;
assign v$EQ20_6669_out0 = v$N_11401_out0 == 5'h13;
assign v$EQ18_8460_out0 = v$N_11398_out0 == 5'h11;
assign v$EQ18_8461_out0 = v$N_11399_out0 == 5'h11;
assign v$EQ18_8462_out0 = v$N_11400_out0 == 5'h11;
assign v$EQ18_8463_out0 = v$N_11401_out0 == 5'h11;
assign v$EQ1_8984_out0 = v$N_11398_out0 == 5'h0;
assign v$EQ1_8985_out0 = v$N_11399_out0 == 5'h0;
assign v$EQ1_8986_out0 = v$N_11400_out0 == 5'h0;
assign v$EQ1_8987_out0 = v$N_11401_out0 == 5'h0;
assign v$EQ9_9300_out0 = v$N_11398_out0 == 5'h9;
assign v$EQ9_9301_out0 = v$N_11399_out0 == 5'h9;
assign v$EQ9_9302_out0 = v$N_11400_out0 == 5'h9;
assign v$EQ9_9303_out0 = v$N_11401_out0 == 5'h9;
assign v$EQ12_9356_out0 = v$N_11398_out0 == 5'hb;
assign v$EQ12_9357_out0 = v$N_11399_out0 == 5'hb;
assign v$EQ12_9358_out0 = v$N_11400_out0 == 5'hb;
assign v$EQ12_9359_out0 = v$N_11401_out0 == 5'hb;
assign v$EQ2_9605_out0 = v$N_11398_out0 == 5'h1;
assign v$EQ2_9606_out0 = v$N_11399_out0 == 5'h1;
assign v$EQ2_9607_out0 = v$N_11400_out0 == 5'h1;
assign v$EQ2_9608_out0 = v$N_11401_out0 == 5'h1;
assign v$EQ8_9797_out0 = v$N_11398_out0 == 5'h7;
assign v$EQ8_9798_out0 = v$N_11399_out0 == 5'h7;
assign v$EQ8_9799_out0 = v$N_11400_out0 == 5'h7;
assign v$EQ8_9800_out0 = v$N_11401_out0 == 5'h7;
assign v$EQ15_11158_out0 = v$N_11398_out0 == 5'he;
assign v$EQ15_11159_out0 = v$N_11399_out0 == 5'he;
assign v$EQ15_11160_out0 = v$N_11400_out0 == 5'he;
assign v$EQ15_11161_out0 = v$N_11401_out0 == 5'he;
assign v$G1_11209_out0 = v$SEL7_4357_out0 || v$SEL6_9304_out0;
assign v$G1_11213_out0 = v$SEL7_4361_out0 || v$SEL6_9308_out0;
assign v$SEL27_11434_out0 = v$NUPPER_12173_out0[0:0];
assign v$SEL27_11435_out0 = v$NUPPER_12174_out0[0:0];
assign v$SEL27_11436_out0 = v$NUPPER_12175_out0[0:0];
assign v$SEL27_11437_out0 = v$NUPPER_12176_out0[0:0];
assign v$SEL29_11666_out0 = v$NUPPER_12173_out0[2:2];
assign v$SEL29_11667_out0 = v$NUPPER_12174_out0[2:2];
assign v$SEL29_11668_out0 = v$NUPPER_12175_out0[2:2];
assign v$SEL29_11669_out0 = v$NUPPER_12176_out0[2:2];
assign v$G2_12962_out0 = v$HIGHER$SAME_6366_out0 && v$LOWER$OUT_4434_out0;
assign v$G2_12963_out0 = v$HIGHER$SAME_6367_out0 && v$LOWER$OUT_4435_out0;
assign v$G2_12964_out0 = v$HIGHER$SAME_6368_out0 && v$LOWER$OUT_4436_out0;
assign v$G2_12965_out0 = v$HIGHER$SAME_6369_out0 && v$LOWER$OUT_4437_out0;
assign v$EQ4_13241_out0 = v$N_11398_out0 == 5'h3;
assign v$EQ4_13242_out0 = v$N_11399_out0 == 5'h3;
assign v$EQ4_13243_out0 = v$N_11400_out0 == 5'h3;
assign v$EQ4_13244_out0 = v$N_11401_out0 == 5'h3;
assign v$RAMDOUT_66_out0 = v$RAMDOUT_5424_out0;
assign v$RAMDOUT_67_out0 = v$RAMDOUT_5425_out0;
assign v$MUX1_1285_out0 = v$LEFT$SHIT_1797_out0 ? v$_2922_out0 : v$_6229_out0;
assign v$MUX1_1317_out0 = v$LEFT$SHIT_1829_out0 ? v$_2954_out0 : v$_6261_out0;
assign v$DIFF_1587_out0 = v$DIFF_244_out0;
assign v$DIFF_1588_out0 = v$DIFF_245_out0;
assign v$OUT_1902_out0 = v$MUX3_1101_out0;
assign v$OUT_1906_out0 = v$MUX3_1105_out0;
assign v$G1_6037_out0 = v$SEL27_11434_out0 || v$SEL28_4925_out0;
assign v$G1_6038_out0 = v$SEL27_11435_out0 || v$SEL28_4926_out0;
assign v$G1_6039_out0 = v$SEL27_11436_out0 || v$SEL28_4927_out0;
assign v$G1_6040_out0 = v$SEL27_11437_out0 || v$SEL28_4928_out0;
assign v$G3_8684_out0 = v$HIGHER$OUT_5318_out0 || v$G2_12962_out0;
assign v$G3_8685_out0 = v$HIGHER$OUT_5319_out0 || v$G2_12963_out0;
assign v$G3_8686_out0 = v$HIGHER$OUT_5320_out0 || v$G2_12964_out0;
assign v$G3_8687_out0 = v$HIGHER$OUT_5321_out0 || v$G2_12965_out0;
assign v$A_10147_out0 = v$A_3663_out0;
assign v$A_10148_out0 = v$A_3664_out0;
assign v$G2_12220_out0 = v$G1_11209_out0 || v$SEL8_11646_out0;
assign v$G2_12224_out0 = v$G1_11213_out0 || v$SEL8_11650_out0;
assign v$RAMDOUT_3669_out0 = v$RAMDOUT_66_out0;
assign v$RAMDOUT_3670_out0 = v$RAMDOUT_67_out0;
assign v$MULTIPLIER_4366_out0 = v$A_10147_out0;
assign v$MULTIPLIER_4367_out0 = v$A_10147_out0;
assign v$MULTIPLIER_4368_out0 = v$A_10147_out0;
assign v$MULTIPLIER_4369_out0 = v$A_10147_out0;
assign v$MULTIPLIER_4370_out0 = v$A_10147_out0;
assign v$MULTIPLIER_4371_out0 = v$A_10147_out0;
assign v$MULTIPLIER_4372_out0 = v$A_10147_out0;
assign v$MULTIPLIER_4373_out0 = v$A_10147_out0;
assign v$MULTIPLIER_4374_out0 = v$A_10147_out0;
assign v$MULTIPLIER_4375_out0 = v$A_10147_out0;
assign v$MULTIPLIER_4376_out0 = v$A_10147_out0;
assign v$MULTIPLIER_4377_out0 = v$A_10147_out0;
assign v$MULTIPLIER_4378_out0 = v$A_10148_out0;
assign v$MULTIPLIER_4379_out0 = v$A_10148_out0;
assign v$MULTIPLIER_4380_out0 = v$A_10148_out0;
assign v$MULTIPLIER_4381_out0 = v$A_10148_out0;
assign v$MULTIPLIER_4382_out0 = v$A_10148_out0;
assign v$MULTIPLIER_4383_out0 = v$A_10148_out0;
assign v$MULTIPLIER_4384_out0 = v$A_10148_out0;
assign v$MULTIPLIER_4385_out0 = v$A_10148_out0;
assign v$MULTIPLIER_4386_out0 = v$A_10148_out0;
assign v$MULTIPLIER_4387_out0 = v$A_10148_out0;
assign v$MULTIPLIER_4388_out0 = v$A_10148_out0;
assign v$MULTIPLIER_4389_out0 = v$A_10148_out0;
assign v$SHIFT$AMOUNT_4981_out0 = v$DIFF_1587_out0;
assign v$SHIFT$AMOUNT_4982_out0 = v$DIFF_1587_out0;
assign v$SHIFT$AMOUNT_4985_out0 = v$DIFF_1588_out0;
assign v$SHIFT$AMOUNT_4986_out0 = v$DIFF_1588_out0;
assign v$OUT_6185_out0 = v$G3_8684_out0;
assign v$OUT_6186_out0 = v$G3_8685_out0;
assign v$OUT_6187_out0 = v$G3_8686_out0;
assign v$OUT_6188_out0 = v$G3_8687_out0;
assign v$G2_7692_out0 = v$G1_6037_out0 || v$SEL29_11666_out0;
assign v$G2_7693_out0 = v$G1_6038_out0 || v$SEL29_11667_out0;
assign v$G2_7694_out0 = v$G1_6039_out0 || v$SEL29_11668_out0;
assign v$G2_7695_out0 = v$G1_6040_out0 || v$SEL29_11669_out0;
assign v$OUT_9893_out0 = v$OUT_1902_out0;
assign v$OUT_9894_out0 = v$OUT_1906_out0;
assign v$MUX2_13217_out0 = v$EN_3585_out0 ? v$MUX1_1285_out0 : v$IN_2566_out0;
assign v$MUX2_13227_out0 = v$EN_3595_out0 ? v$MUX1_1317_out0 : v$IN_2576_out0;
assign v$SEL3_438_out0 = v$SHIFT$AMOUNT_4981_out0[2:2];
assign v$SEL3_439_out0 = v$SHIFT$AMOUNT_4982_out0[2:2];
assign v$SEL3_442_out0 = v$SHIFT$AMOUNT_4985_out0[2:2];
assign v$SEL3_443_out0 = v$SHIFT$AMOUNT_4986_out0[2:2];
assign v$SEL1_1192_out0 = v$SHIFT$AMOUNT_4981_out0[0:0];
assign v$SEL1_1193_out0 = v$SHIFT$AMOUNT_4982_out0[0:0];
assign v$SEL1_1196_out0 = v$SHIFT$AMOUNT_4985_out0[0:0];
assign v$SEL1_1197_out0 = v$SHIFT$AMOUNT_4986_out0[0:0];
assign v$G3_3149_out0 = v$OUT_6186_out0 && v$SAME$H_6167_out0;
assign v$G3_3150_out0 = v$OUT_6188_out0 && v$SAME$H_6168_out0;
assign v$SEL4_3331_out0 = v$SHIFT$AMOUNT_4981_out0[3:3];
assign v$SEL4_3332_out0 = v$SHIFT$AMOUNT_4982_out0[3:3];
assign v$SEL4_3335_out0 = v$SHIFT$AMOUNT_4985_out0[3:3];
assign v$SEL4_3336_out0 = v$SHIFT$AMOUNT_4986_out0[3:3];
assign v$SEL7_4358_out0 = v$SHIFT$AMOUNT_4981_out0[5:5];
assign v$SEL7_4359_out0 = v$SHIFT$AMOUNT_4982_out0[5:5];
assign v$SEL7_4362_out0 = v$SHIFT$AMOUNT_4985_out0[5:5];
assign v$SEL7_4363_out0 = v$SHIFT$AMOUNT_4986_out0[5:5];
assign v$OP2_6767_out0 = v$OUT_9893_out0;
assign v$OP2_6768_out0 = v$OUT_9894_out0;
assign v$SEL1_7324_out0 = v$MULTIPLIER_4366_out0[12:12];
assign v$SEL1_7325_out0 = v$MULTIPLIER_4367_out0[1:1];
assign v$SEL1_7326_out0 = v$MULTIPLIER_4368_out0[8:8];
assign v$SEL1_7327_out0 = v$MULTIPLIER_4369_out0[10:10];
assign v$SEL1_7328_out0 = v$MULTIPLIER_4370_out0[9:9];
assign v$SEL1_7329_out0 = v$MULTIPLIER_4371_out0[11:11];
assign v$SEL1_7330_out0 = v$MULTIPLIER_4372_out0[7:7];
assign v$SEL1_7331_out0 = v$MULTIPLIER_4373_out0[2:2];
assign v$SEL1_7332_out0 = v$MULTIPLIER_4374_out0[6:6];
assign v$SEL1_7333_out0 = v$MULTIPLIER_4375_out0[3:3];
assign v$SEL1_7334_out0 = v$MULTIPLIER_4376_out0[4:4];
assign v$SEL1_7335_out0 = v$MULTIPLIER_4377_out0[5:5];
assign v$SEL1_7336_out0 = v$MULTIPLIER_4378_out0[12:12];
assign v$SEL1_7337_out0 = v$MULTIPLIER_4379_out0[1:1];
assign v$SEL1_7338_out0 = v$MULTIPLIER_4380_out0[8:8];
assign v$SEL1_7339_out0 = v$MULTIPLIER_4381_out0[10:10];
assign v$SEL1_7340_out0 = v$MULTIPLIER_4382_out0[9:9];
assign v$SEL1_7341_out0 = v$MULTIPLIER_4383_out0[11:11];
assign v$SEL1_7342_out0 = v$MULTIPLIER_4384_out0[7:7];
assign v$SEL1_7343_out0 = v$MULTIPLIER_4385_out0[2:2];
assign v$SEL1_7344_out0 = v$MULTIPLIER_4386_out0[6:6];
assign v$SEL1_7345_out0 = v$MULTIPLIER_4387_out0[3:3];
assign v$SEL1_7346_out0 = v$MULTIPLIER_4388_out0[4:4];
assign v$SEL1_7347_out0 = v$MULTIPLIER_4389_out0[5:5];
assign v$SEL2_7442_out0 = v$MULTIPLIER_4367_out0[13:13];
assign v$SEL2_7443_out0 = v$MULTIPLIER_4368_out0[20:20];
assign v$SEL2_7444_out0 = v$MULTIPLIER_4369_out0[22:22];
assign v$SEL2_7445_out0 = v$MULTIPLIER_4370_out0[21:21];
assign v$SEL2_7446_out0 = v$MULTIPLIER_4371_out0[23:23];
assign v$SEL2_7447_out0 = v$MULTIPLIER_4372_out0[19:19];
assign v$SEL2_7448_out0 = v$MULTIPLIER_4373_out0[14:14];
assign v$SEL2_7449_out0 = v$MULTIPLIER_4374_out0[18:18];
assign v$SEL2_7450_out0 = v$MULTIPLIER_4375_out0[15:15];
assign v$SEL2_7451_out0 = v$MULTIPLIER_4376_out0[16:16];
assign v$SEL2_7452_out0 = v$MULTIPLIER_4377_out0[17:17];
assign v$SEL2_7453_out0 = v$MULTIPLIER_4379_out0[13:13];
assign v$SEL2_7454_out0 = v$MULTIPLIER_4380_out0[20:20];
assign v$SEL2_7455_out0 = v$MULTIPLIER_4381_out0[22:22];
assign v$SEL2_7456_out0 = v$MULTIPLIER_4382_out0[21:21];
assign v$SEL2_7457_out0 = v$MULTIPLIER_4383_out0[23:23];
assign v$SEL2_7458_out0 = v$MULTIPLIER_4384_out0[19:19];
assign v$SEL2_7459_out0 = v$MULTIPLIER_4385_out0[14:14];
assign v$SEL2_7460_out0 = v$MULTIPLIER_4386_out0[18:18];
assign v$SEL2_7461_out0 = v$MULTIPLIER_4387_out0[15:15];
assign v$SEL2_7462_out0 = v$MULTIPLIER_4388_out0[16:16];
assign v$SEL2_7463_out0 = v$MULTIPLIER_4389_out0[17:17];
assign v$MUX2_7752_out0 = v$G24_12707_out0 ? v$RAMDOUT_3669_out0 : v$RMN_4169_out0;
assign v$MUX2_7753_out0 = v$G24_12708_out0 ? v$RAMDOUT_3670_out0 : v$RMN_4170_out0;
assign v$SEL5_7989_out0 = v$SHIFT$AMOUNT_4981_out0[4:4];
assign v$SEL5_7990_out0 = v$SHIFT$AMOUNT_4982_out0[4:4];
assign v$SEL5_7993_out0 = v$SHIFT$AMOUNT_4985_out0[4:4];
assign v$SEL5_7994_out0 = v$SHIFT$AMOUNT_4986_out0[4:4];
assign v$SEL6_9305_out0 = v$SHIFT$AMOUNT_4981_out0[6:6];
assign v$SEL6_9306_out0 = v$SHIFT$AMOUNT_4982_out0[6:6];
assign v$SEL6_9309_out0 = v$SHIFT$AMOUNT_4985_out0[6:6];
assign v$SEL6_9310_out0 = v$SHIFT$AMOUNT_4986_out0[6:6];
assign v$OUT_10236_out0 = v$MUX2_13217_out0;
assign v$OUT_10268_out0 = v$MUX2_13227_out0;
assign v$SEL8_11647_out0 = v$SHIFT$AMOUNT_4981_out0[7:7];
assign v$SEL8_11648_out0 = v$SHIFT$AMOUNT_4982_out0[7:7];
assign v$SEL8_11651_out0 = v$SHIFT$AMOUNT_4985_out0[7:7];
assign v$SEL8_11652_out0 = v$SHIFT$AMOUNT_4986_out0[7:7];
assign v$SEL2_13057_out0 = v$SHIFT$AMOUNT_4981_out0[1:1];
assign v$SEL2_13058_out0 = v$SHIFT$AMOUNT_4982_out0[1:1];
assign v$SEL2_13061_out0 = v$SHIFT$AMOUNT_4985_out0[1:1];
assign v$SEL2_13062_out0 = v$SHIFT$AMOUNT_4986_out0[1:1];
assign v$EN_565_out0 = v$SEL5_7989_out0;
assign v$EN_566_out0 = v$SEL4_3331_out0;
assign v$EN_567_out0 = v$SEL5_7990_out0;
assign v$EN_568_out0 = v$SEL4_3332_out0;
assign v$EN_575_out0 = v$SEL5_7993_out0;
assign v$EN_576_out0 = v$SEL4_3335_out0;
assign v$EN_577_out0 = v$SEL5_7994_out0;
assign v$EN_578_out0 = v$SEL4_3336_out0;
assign v$MULTIPLYING$BIT_1607_out0 = v$SEL1_7324_out0;
assign v$MULTIPLYING$BIT_1619_out0 = v$SEL1_7336_out0;
assign v$EN_3168_out0 = v$SEL3_438_out0;
assign v$EN_3169_out0 = v$SEL3_439_out0;
assign v$EN_3174_out0 = v$SEL3_442_out0;
assign v$EN_3175_out0 = v$SEL3_443_out0;
assign v$IN_3525_out0 = v$OUT_10236_out0;
assign v$IN_3557_out0 = v$OUT_10268_out0;
assign v$EN_3592_out0 = v$SEL1_1192_out0;
assign v$EN_3593_out0 = v$SEL1_1193_out0;
assign v$EN_3602_out0 = v$SEL1_1196_out0;
assign v$EN_3603_out0 = v$SEL1_1197_out0;
assign v$EN_5392_out0 = v$SEL2_13057_out0;
assign v$EN_5393_out0 = v$SEL2_13058_out0;
assign v$EN_5398_out0 = v$SEL2_13061_out0;
assign v$EN_5399_out0 = v$SEL2_13062_out0;
assign v$OP2_10356_out0 = v$OP2_6767_out0;
assign v$OP2_10357_out0 = v$OP2_6768_out0;
assign v$G1_10855_out0 = v$G3_3149_out0 || v$OUT_6185_out0;
assign v$G1_10856_out0 = v$G3_3150_out0 || v$OUT_6187_out0;
assign v$G1_11210_out0 = v$SEL7_4358_out0 || v$SEL6_9305_out0;
assign v$G1_11211_out0 = v$SEL7_4359_out0 || v$SEL6_9306_out0;
assign v$G1_11214_out0 = v$SEL7_4362_out0 || v$SEL6_9309_out0;
assign v$G1_11215_out0 = v$SEL7_4363_out0 || v$SEL6_9310_out0;
assign v$MUX1_12005_out0 = v$EXEC1_5456_out0 ? v$SEL1_7325_out0 : v$SEL2_7442_out0;
assign v$MUX1_12006_out0 = v$EXEC1_5457_out0 ? v$SEL1_7326_out0 : v$SEL2_7443_out0;
assign v$MUX1_12007_out0 = v$EXEC1_5458_out0 ? v$SEL1_7327_out0 : v$SEL2_7444_out0;
assign v$MUX1_12008_out0 = v$EXEC1_5459_out0 ? v$SEL1_7328_out0 : v$SEL2_7445_out0;
assign v$MUX1_12009_out0 = v$EXEC1_5460_out0 ? v$SEL1_7329_out0 : v$SEL2_7446_out0;
assign v$MUX1_12010_out0 = v$EXEC1_5461_out0 ? v$SEL1_7330_out0 : v$SEL2_7447_out0;
assign v$MUX1_12011_out0 = v$EXEC1_5462_out0 ? v$SEL1_7331_out0 : v$SEL2_7448_out0;
assign v$MUX1_12012_out0 = v$EXEC1_5463_out0 ? v$SEL1_7332_out0 : v$SEL2_7449_out0;
assign v$MUX1_12013_out0 = v$EXEC1_5464_out0 ? v$SEL1_7333_out0 : v$SEL2_7450_out0;
assign v$MUX1_12014_out0 = v$EXEC1_5465_out0 ? v$SEL1_7334_out0 : v$SEL2_7451_out0;
assign v$MUX1_12015_out0 = v$EXEC1_5466_out0 ? v$SEL1_7335_out0 : v$SEL2_7452_out0;
assign v$MUX1_12016_out0 = v$EXEC1_5467_out0 ? v$SEL1_7337_out0 : v$SEL2_7453_out0;
assign v$MUX1_12017_out0 = v$EXEC1_5468_out0 ? v$SEL1_7338_out0 : v$SEL2_7454_out0;
assign v$MUX1_12018_out0 = v$EXEC1_5469_out0 ? v$SEL1_7339_out0 : v$SEL2_7455_out0;
assign v$MUX1_12019_out0 = v$EXEC1_5470_out0 ? v$SEL1_7340_out0 : v$SEL2_7456_out0;
assign v$MUX1_12020_out0 = v$EXEC1_5471_out0 ? v$SEL1_7341_out0 : v$SEL2_7457_out0;
assign v$MUX1_12021_out0 = v$EXEC1_5472_out0 ? v$SEL1_7342_out0 : v$SEL2_7458_out0;
assign v$MUX1_12022_out0 = v$EXEC1_5473_out0 ? v$SEL1_7343_out0 : v$SEL2_7459_out0;
assign v$MUX1_12023_out0 = v$EXEC1_5474_out0 ? v$SEL1_7344_out0 : v$SEL2_7460_out0;
assign v$MUX1_12024_out0 = v$EXEC1_5475_out0 ? v$SEL1_7345_out0 : v$SEL2_7461_out0;
assign v$MUX1_12025_out0 = v$EXEC1_5476_out0 ? v$SEL1_7346_out0 : v$SEL2_7462_out0;
assign v$MUX1_12026_out0 = v$EXEC1_5477_out0 ? v$SEL1_7347_out0 : v$SEL2_7463_out0;
assign v$REGDIN_13076_out0 = v$MUX2_7752_out0;
assign v$REGDIN_13077_out0 = v$MUX2_7753_out0;
assign v$MULTIPLYING$BIT_1608_out0 = v$MUX1_12005_out0;
assign v$MULTIPLYING$BIT_1609_out0 = v$MUX1_12006_out0;
assign v$MULTIPLYING$BIT_1610_out0 = v$MUX1_12007_out0;
assign v$MULTIPLYING$BIT_1611_out0 = v$MUX1_12008_out0;
assign v$MULTIPLYING$BIT_1612_out0 = v$MUX1_12009_out0;
assign v$MULTIPLYING$BIT_1613_out0 = v$MUX1_12010_out0;
assign v$MULTIPLYING$BIT_1614_out0 = v$MUX1_12011_out0;
assign v$MULTIPLYING$BIT_1615_out0 = v$MUX1_12012_out0;
assign v$MULTIPLYING$BIT_1616_out0 = v$MUX1_12013_out0;
assign v$MULTIPLYING$BIT_1617_out0 = v$MUX1_12014_out0;
assign v$MULTIPLYING$BIT_1618_out0 = v$MUX1_12015_out0;
assign v$MULTIPLYING$BIT_1620_out0 = v$MUX1_12016_out0;
assign v$MULTIPLYING$BIT_1621_out0 = v$MUX1_12017_out0;
assign v$MULTIPLYING$BIT_1622_out0 = v$MUX1_12018_out0;
assign v$MULTIPLYING$BIT_1623_out0 = v$MUX1_12019_out0;
assign v$MULTIPLYING$BIT_1624_out0 = v$MUX1_12020_out0;
assign v$MULTIPLYING$BIT_1625_out0 = v$MUX1_12021_out0;
assign v$MULTIPLYING$BIT_1626_out0 = v$MUX1_12022_out0;
assign v$MULTIPLYING$BIT_1627_out0 = v$MUX1_12023_out0;
assign v$MULTIPLYING$BIT_1628_out0 = v$MUX1_12024_out0;
assign v$MULTIPLYING$BIT_1629_out0 = v$MUX1_12025_out0;
assign v$MULTIPLYING$BIT_1630_out0 = v$MUX1_12026_out0;
assign v$OUT_2549_out0 = v$G1_10855_out0;
assign v$OUT_2550_out0 = v$G1_10856_out0;
assign v$OP2_5118_out0 = v$OP2_10356_out0;
assign v$OP2_5119_out0 = v$OP2_10357_out0;
assign v$IN_7582_out0 = v$IN_3525_out0;
assign v$IN_7588_out0 = v$IN_3557_out0;
assign v$REGDIN_11576_out0 = v$REGDIN_13076_out0;
assign v$REGDIN_11577_out0 = v$REGDIN_13077_out0;
assign v$G2_12221_out0 = v$G1_11210_out0 || v$SEL8_11647_out0;
assign v$G2_12222_out0 = v$G1_11211_out0 || v$SEL8_11648_out0;
assign v$G2_12225_out0 = v$G1_11214_out0 || v$SEL8_11651_out0;
assign v$G2_12226_out0 = v$G1_11215_out0 || v$SEL8_11652_out0;
assign v$SEL1_5938_out0 = v$IN_7582_out0[23:2];
assign v$SEL1_5970_out0 = v$IN_7588_out0[23:2];
assign v$XOR1_6518_out0 = v$OP2_5118_out0 ^ v$MUX1_12538_out0;
assign v$XOR1_6519_out0 = v$OP2_5119_out0 ^ v$MUX1_12539_out0;
assign v$B_7540_out0 = v$OP2_5118_out0;
assign v$B_7541_out0 = v$OP2_5119_out0;
assign v$SEL1_10682_out0 = v$IN_7582_out0[21:0];
assign v$SEL1_10714_out0 = v$IN_7588_out0[21:0];
assign v$A$MANTISA$LARGER_11207_out0 = v$OUT_2549_out0;
assign v$A$MANTISA$LARGER_11208_out0 = v$OUT_2550_out0;
assign v$_2924_out0 = { v$C2_100_out0,v$SEL1_10682_out0 };
assign v$_2956_out0 = { v$C2_132_out0,v$SEL1_10714_out0 };
assign v$_6231_out0 = { v$SEL1_5938_out0,v$C1_3967_out0 };
assign v$_6263_out0 = { v$SEL1_5970_out0,v$C1_3999_out0 };
assign {v$A1_6425_out1,v$A1_6425_out0 } = v$OP1_3661_out0 + v$XOR1_6518_out0 + v$MUX2_8006_out0;
assign {v$A1_6426_out1,v$A1_6426_out0 } = v$OP1_3662_out0 + v$XOR1_6519_out0 + v$MUX2_8007_out0;
assign v$B_6722_out0 = v$B_7540_out0;
assign v$B_6723_out0 = v$B_7541_out0;
assign v$G7_13277_out0 = v$A$MANTISA$LARGER_11207_out0 && v$EXP$SAME_408_out0;
assign v$G7_13278_out0 = v$A$MANTISA$LARGER_11208_out0 && v$EXP$SAME_409_out0;
assign v$MUX1_1287_out0 = v$LEFT$SHIT_1799_out0 ? v$_2924_out0 : v$_6231_out0;
assign v$MUX1_1319_out0 = v$LEFT$SHIT_1831_out0 ? v$_2956_out0 : v$_6263_out0;
assign v$ADDEROUT_2206_out0 = v$A1_6425_out0;
assign v$ADDEROUT_2207_out0 = v$A1_6426_out0;
assign v$_3609_out0 = v$B_6722_out0[7:4];
assign v$_3610_out0 = v$B_6723_out0[7:4];
assign v$_4355_out0 = v$B_6722_out0[11:8];
assign v$_4356_out0 = v$B_6723_out0[11:8];
assign v$G9_11973_out0 = v$A$EXP$LARGER_12968_out0 || v$G7_13277_out0;
assign v$G9_11974_out0 = v$A$EXP$LARGER_12969_out0 || v$G7_13278_out0;
assign v$_12972_out0 = v$B_6722_out0[15:12];
assign v$_12973_out0 = v$B_6723_out0[15:12];
assign v$_13249_out0 = v$B_6722_out0[3:0];
assign v$_13250_out0 = v$B_6723_out0[3:0];
assign v$_50_out0 = v$_13249_out0[1:0];
assign v$_50_out1 = v$_13249_out0[3:2];
assign v$_51_out0 = v$_13250_out0[1:0];
assign v$_51_out1 = v$_13250_out0[3:2];
assign v$_199_out0 = v$_3609_out0[1:0];
assign v$_199_out1 = v$_3609_out0[3:2];
assign v$_200_out0 = v$_3610_out0[1:0];
assign v$_200_out1 = v$_3610_out0[3:2];
assign v$_705_out0 = v$_12972_out0[1:0];
assign v$_705_out1 = v$_12972_out0[3:2];
assign v$_706_out0 = v$_12973_out0[1:0];
assign v$_706_out1 = v$_12973_out0[3:2];
assign v$MUX2_1393_out0 = v$EN_5389_out0 ? v$MUX1_1287_out0 : v$IN_7582_out0;
assign v$MUX2_1399_out0 = v$EN_5395_out0 ? v$MUX1_1319_out0 : v$IN_7588_out0;
assign v$_5044_out0 = v$_4355_out0[1:0];
assign v$_5044_out1 = v$_4355_out0[3:2];
assign v$_5045_out0 = v$_4356_out0[1:0];
assign v$_5045_out1 = v$_4356_out0[3:2];
assign v$IS$A$LARGER_11880_out0 = v$G9_11973_out0;
assign v$IS$A$LARGER_11881_out0 = v$G9_11974_out0;
assign v$G8_211_out0 = v$IS$A$LARGER_11880_out0 || v$IS$SUB_3087_out0;
assign v$G8_212_out0 = v$IS$A$LARGER_11881_out0 || v$IS$SUB_3088_out0;
assign v$MUX11_487_out0 = v$IS$A$LARGER_11880_out0 ? v$SEL5_260_out0 : v$G1_10445_out0;
assign v$MUX11_488_out0 = v$IS$A$LARGER_11881_out0 ? v$SEL5_261_out0 : v$G1_10446_out0;
assign v$_3433_out0 = v$_50_out1[0:0];
assign v$_3433_out1 = v$_50_out1[1:1];
assign v$_3434_out0 = v$_51_out1[0:0];
assign v$_3434_out1 = v$_51_out1[1:1];
assign v$MUX15_4768_out0 = v$IS$A$LARGER_11880_out0 ? v$A_1951_out0 : v$B_12546_out0;
assign v$MUX15_4769_out0 = v$IS$A$LARGER_11881_out0 ? v$A_1952_out0 : v$B_12547_out0;
assign v$IS$A$LARGER_4806_out0 = v$IS$A$LARGER_11880_out0;
assign v$IS$A$LARGER_4807_out0 = v$IS$A$LARGER_11881_out0;
assign v$_4988_out0 = v$_199_out1[0:0];
assign v$_4988_out1 = v$_199_out1[1:1];
assign v$_4989_out0 = v$_200_out1[0:0];
assign v$_4989_out1 = v$_200_out1[1:1];
assign v$_6308_out0 = v$_199_out0[0:0];
assign v$_6308_out1 = v$_199_out0[1:1];
assign v$_6309_out0 = v$_200_out0[0:0];
assign v$_6309_out1 = v$_200_out0[1:1];
assign v$_6349_out0 = v$_5044_out0[0:0];
assign v$_6349_out1 = v$_5044_out0[1:1];
assign v$_6350_out0 = v$_5045_out0[0:0];
assign v$_6350_out1 = v$_5045_out0[1:1];
assign v$_10014_out0 = v$_50_out0[0:0];
assign v$_10014_out1 = v$_50_out0[1:1];
assign v$_10015_out0 = v$_51_out0[0:0];
assign v$_10015_out1 = v$_51_out0[1:1];
assign v$OUT_10238_out0 = v$MUX2_1393_out0;
assign v$OUT_10270_out0 = v$MUX2_1399_out0;
assign v$_10493_out0 = v$_705_out0[0:0];
assign v$_10493_out1 = v$_705_out0[1:1];
assign v$_10494_out0 = v$_706_out0[0:0];
assign v$_10494_out1 = v$_706_out0[1:1];
assign v$_10627_out0 = v$_705_out1[0:0];
assign v$_10627_out1 = v$_705_out1[1:1];
assign v$_10628_out0 = v$_706_out1[0:0];
assign v$_10628_out1 = v$_706_out1[1:1];
assign v$G2_10819_out0 = v$IS$A$LARGER_11880_out0 && v$IS$SUB_3087_out0;
assign v$G2_10820_out0 = v$IS$A$LARGER_11881_out0 && v$IS$SUB_3088_out0;
assign v$_11302_out0 = v$_5044_out1[0:0];
assign v$_11302_out1 = v$_5044_out1[1:1];
assign v$_11303_out0 = v$_5045_out1[0:0];
assign v$_11303_out1 = v$_5045_out1[1:1];
assign v$MUX16_13179_out0 = v$IS$A$LARGER_11880_out0 ? v$A_1951_out0 : v$B_12546_out0;
assign v$MUX16_13180_out0 = v$IS$A$LARGER_11881_out0 ? v$A_1952_out0 : v$B_12547_out0;
assign v$G14_867_out0 = v$_11630_out1 && v$_10493_out1;
assign v$G14_868_out0 = v$_11631_out1 && v$_10494_out1;
assign v$G13_883_out0 = v$_11630_out0 && v$_10493_out0;
assign v$G13_884_out0 = v$_11631_out0 && v$_10494_out0;
assign v$G5_1162_out0 = v$_2736_out0 && v$_6308_out0;
assign v$G5_1163_out0 = v$_2737_out0 && v$_6309_out0;
assign v$G6_1174_out0 = v$_2736_out1 && v$_6308_out1;
assign v$G6_1175_out0 = v$_2737_out1 && v$_6309_out1;
assign v$G9_2141_out0 = v$_266_out0 && v$_6349_out0;
assign v$G9_2142_out0 = v$_267_out0 && v$_6350_out0;
assign v$A$IS$OP1_3397_out0 = v$G8_211_out0;
assign v$A$IS$OP1_3398_out0 = v$G8_212_out0;
assign v$IN_3524_out0 = v$OUT_10238_out0;
assign v$IN_3556_out0 = v$OUT_10270_out0;
assign v$SEL17_3633_out0 = v$MUX16_13179_out0[14:7];
assign v$SEL17_3634_out0 = v$MUX16_13180_out0[14:7];
assign v$G11_5694_out0 = v$_3284_out0 && v$_11302_out0;
assign v$G11_5695_out0 = v$_3285_out0 && v$_11303_out0;
assign v$G2_6316_out0 = v$_7294_out1 && v$_10014_out1;
assign v$G2_6317_out0 = v$_7295_out1 && v$_10015_out1;
assign v$G8_6322_out0 = v$_6815_out1 && v$_4988_out1;
assign v$G8_6323_out0 = v$_6816_out1 && v$_4989_out1;
assign v$IS$A$LARGER_6990_out0 = v$IS$A$LARGER_4806_out0;
assign v$IS$A$LARGER_6991_out0 = v$IS$A$LARGER_4807_out0;
assign v$G4_7665_out0 = v$G2_10819_out0 && v$G5_11019_out0;
assign v$G4_7666_out0 = v$G2_10820_out0 && v$G5_11020_out0;
assign v$SUBTRACTION$SIGN_7667_out0 = v$MUX11_487_out0;
assign v$SUBTRACTION$SIGN_7668_out0 = v$MUX11_488_out0;
assign v$G1_7899_out0 = v$_7294_out0 && v$_10014_out0;
assign v$G1_7900_out0 = v$_7295_out0 && v$_10015_out0;
assign v$G7_7976_out0 = v$_6815_out0 && v$_4988_out0;
assign v$G7_7977_out0 = v$_6816_out0 && v$_4989_out0;
assign v$G3_8587_out0 = v$_3651_out0 && v$_3433_out0;
assign v$G3_8588_out0 = v$_3652_out0 && v$_3434_out0;
assign v$G12_9318_out0 = v$_3284_out1 && v$_11302_out1;
assign v$G12_9319_out0 = v$_3285_out1 && v$_11303_out1;
assign v$G4_9889_out0 = v$_3651_out1 && v$_3433_out1;
assign v$G4_9890_out0 = v$_3652_out1 && v$_3434_out1;
assign v$G15_9960_out0 = v$_1868_out0 && v$_10627_out0;
assign v$G15_9961_out0 = v$_1869_out0 && v$_10628_out0;
assign v$SEL3_12563_out0 = v$MUX15_4768_out0[14:7];
assign v$SEL3_12564_out0 = v$MUX15_4769_out0[14:7];
assign v$SEL18_12974_out0 = v$MUX16_13179_out0[14:10];
assign v$SEL18_12975_out0 = v$MUX16_13180_out0[14:10];
assign v$G10_13153_out0 = v$_266_out1 && v$_6349_out1;
assign v$G10_13154_out0 = v$_267_out1 && v$_6350_out1;
assign v$G16_13408_out0 = v$_1868_out1 && v$_10627_out1;
assign v$G16_13409_out0 = v$_1869_out1 && v$_10628_out1;
assign v$MUX9_1381_out0 = v$A$IS$OP1_3397_out0 ? v$B$MANTISA_10857_out0 : v$A$MANTISA_2469_out0;
assign v$MUX9_1382_out0 = v$A$IS$OP1_3398_out0 ? v$B$MANTISA_10858_out0 : v$A$MANTISA_2470_out0;
assign v$_1879_out0 = { v$G15_9960_out0,v$G16_13408_out0 };
assign v$_1880_out0 = { v$G15_9961_out0,v$G16_13409_out0 };
assign v$_6453_out0 = { v$G7_7976_out0,v$G8_6322_out0 };
assign v$_6454_out0 = { v$G7_7977_out0,v$G8_6323_out0 };
assign v$_7233_out0 = { v$G3_8587_out0,v$G4_9889_out0 };
assign v$_7234_out0 = { v$G3_8588_out0,v$G4_9890_out0 };
assign v$SINGLE$PRECISION$EXPONENT_7284_out0 = v$SEL3_12563_out0;
assign v$SINGLE$PRECISION$EXPONENT_7285_out0 = v$SEL3_12564_out0;
assign v$MUX3_8454_out0 = v$A$IS$OP1_3397_out0 ? v$A$MANTISA_2469_out0 : v$B$MANTISA_10857_out0;
assign v$MUX3_8455_out0 = v$A$IS$OP1_3398_out0 ? v$A$MANTISA_2470_out0 : v$B$MANTISA_10858_out0;
assign v$EXPONENT_9232_out0 = v$SEL17_3633_out0;
assign v$EXPONENT_9233_out0 = v$SEL17_3634_out0;
assign v$_9554_out0 = { v$G1_7899_out0,v$G2_6316_out0 };
assign v$_9555_out0 = { v$G1_7900_out0,v$G2_6317_out0 };
assign v$_9609_out0 = { v$G5_1162_out0,v$G6_1174_out0 };
assign v$_9610_out0 = { v$G5_1163_out0,v$G6_1175_out0 };
assign v$IN_10872_out0 = v$IN_3524_out0;
assign v$IN_10878_out0 = v$IN_3556_out0;
assign v$G1_11011_out0 = ! v$IS$A$LARGER_6990_out0;
assign v$G1_11012_out0 = ! v$IS$A$LARGER_6991_out0;
assign v$_11188_out0 = { v$G11_5694_out0,v$G12_9318_out0 };
assign v$_11189_out0 = { v$G11_5695_out0,v$G12_9319_out0 };
assign v$EXPONENT_11194_out0 = v$SEL18_12974_out0;
assign v$EXPONENT_11195_out0 = v$SEL18_12975_out0;
assign v$_11823_out0 = { v$G9_2141_out0,v$G10_13153_out0 };
assign v$_11824_out0 = { v$G9_2142_out0,v$G10_13154_out0 };
assign v$MUX4_12532_out0 = v$G4_7665_out0 ? v$A_1951_out0 : v$B_12546_out0;
assign v$MUX4_12533_out0 = v$G4_7666_out0 ? v$A_1952_out0 : v$B_12547_out0;
assign v$_13213_out0 = { v$G13_883_out0,v$G14_867_out0 };
assign v$_13214_out0 = { v$G13_884_out0,v$G14_868_out0 };
assign v$_223_out0 = { v$_13213_out0,v$_1879_out0 };
assign v$_224_out0 = { v$_13214_out0,v$_1880_out0 };
assign v$EXPONENT_583_out0 = v$SINGLE$PRECISION$EXPONENT_7284_out0;
assign v$EXPONENT_584_out0 = v$SINGLE$PRECISION$EXPONENT_7285_out0;
assign v$_2419_out0 = { v$_11823_out0,v$_11188_out0 };
assign v$_2420_out0 = { v$_11824_out0,v$_11189_out0 };
assign v$SEL1_5937_out0 = v$IN_10872_out0[23:4];
assign v$SEL1_5969_out0 = v$IN_10878_out0[23:4];
assign v$OP1$MANTISA_6355_out0 = v$MUX3_8454_out0;
assign v$OP1$MANTISA_6356_out0 = v$MUX3_8455_out0;
assign v$SEL1_6461_out0 = v$MUX4_12532_out0[14:10];
assign v$SEL1_6462_out0 = v$MUX4_12533_out0[14:10];
assign v$OP2$MANTISA_6520_out0 = v$MUX9_1381_out0;
assign v$OP2$MANTISA_6521_out0 = v$MUX9_1382_out0;
assign v$_8636_out0 = { v$_9609_out0,v$_6453_out0 };
assign v$_8637_out0 = { v$_9610_out0,v$_6454_out0 };
assign v$SEL1_10681_out0 = v$IN_10872_out0[19:0];
assign v$SEL1_10713_out0 = v$IN_10878_out0[19:0];
assign v$G2_11580_out0 = v$IS$SUB_8690_out0 && v$G1_11011_out0;
assign v$G2_11581_out0 = v$IS$SUB_8691_out0 && v$G1_11012_out0;
assign v$_11935_out0 = { v$_9554_out0,v$_7233_out0 };
assign v$_11936_out0 = { v$_9555_out0,v$_7234_out0 };
assign v$C0_190_out0 = v$_11935_out0;
assign v$C0_191_out0 = v$_11936_out0;
assign v$OP2$MANTISA_1558_out0 = v$OP2$MANTISA_6520_out0;
assign v$OP2$MANTISA_1559_out0 = v$OP2$MANTISA_6521_out0;
assign v$C12_1981_out0 = v$_223_out0;
assign v$C12_1982_out0 = v$_224_out0;
assign v$OP1$MANTISA_2497_out0 = v$OP1$MANTISA_6355_out0;
assign v$OP1$MANTISA_2498_out0 = v$OP1$MANTISA_6356_out0;
assign v$_2923_out0 = { v$C2_99_out0,v$SEL1_10681_out0 };
assign v$_2955_out0 = { v$C2_131_out0,v$SEL1_10713_out0 };
assign v$NEED$SHIFT$OP1_3226_out0 = v$G2_11580_out0;
assign v$NEED$SHIFT$OP1_3227_out0 = v$G2_11581_out0;
assign v$HALF$PRECISION$EXPONENT_4401_out0 = v$SEL1_6461_out0;
assign v$HALF$PRECISION$EXPONENT_4402_out0 = v$SEL1_6462_out0;
assign v$C8_5798_out0 = v$_2419_out0;
assign v$C8_5799_out0 = v$_2420_out0;
assign v$_6230_out0 = { v$SEL1_5937_out0,v$C1_3966_out0 };
assign v$_6262_out0 = { v$SEL1_5969_out0,v$C1_3998_out0 };
assign v$C4_7090_out0 = v$_8636_out0;
assign v$C4_7091_out0 = v$_8637_out0;
assign v$MUX1_1286_out0 = v$LEFT$SHIT_1798_out0 ? v$_2923_out0 : v$_6230_out0;
assign v$MUX1_1318_out0 = v$LEFT$SHIT_1830_out0 ? v$_2955_out0 : v$_6262_out0;
assign v$OP2$MANTISA_2212_out0 = v$OP2$MANTISA_1558_out0;
assign v$OP2$MANTISA_2213_out0 = v$OP2$MANTISA_1559_out0;
assign v$_2402_out0 = { v$C0_190_out0,v$C4_7090_out0 };
assign v$_2403_out0 = { v$C0_191_out0,v$C4_7091_out0 };
assign v$_6291_out0 = { v$C8_5798_out0,v$C12_1981_out0 };
assign v$_6292_out0 = { v$C8_5799_out0,v$C12_1982_out0 };
assign v$OP1$MANTISA_7606_out0 = v$OP1$MANTISA_2497_out0;
assign v$OP1$MANTISA_7607_out0 = v$OP1$MANTISA_2498_out0;
assign v$EXPONENT_11500_out0 = v$HALF$PRECISION$EXPONENT_4401_out0;
assign v$EXPONENT_11501_out0 = v$HALF$PRECISION$EXPONENT_4402_out0;
assign v$IN_8775_out0 = v$OP2$MANTISA_2212_out0;
assign v$IN_8776_out0 = v$OP1$MANTISA_7606_out0;
assign v$IN_8779_out0 = v$OP2$MANTISA_2213_out0;
assign v$IN_8780_out0 = v$OP1$MANTISA_7607_out0;
assign v$MUX2_10555_out0 = v$EN_3165_out0 ? v$MUX1_1286_out0 : v$IN_10872_out0;
assign v$MUX2_10561_out0 = v$EN_3171_out0 ? v$MUX1_1318_out0 : v$IN_10878_out0;
assign v$_11479_out0 = { v$_2402_out0,v$_6291_out0 };
assign v$_11480_out0 = { v$_2403_out0,v$_6292_out0 };
assign v$IN_3540_out0 = v$IN_8775_out0;
assign v$IN_3545_out0 = v$IN_8776_out0;
assign v$IN_3572_out0 = v$IN_8779_out0;
assign v$IN_3577_out0 = v$IN_8780_out0;
assign v$OUT_10237_out0 = v$MUX2_10555_out0;
assign v$OUT_10269_out0 = v$MUX2_10561_out0;
assign v$C_12847_out0 = v$_11479_out0;
assign v$C_12848_out0 = v$_11480_out0;
assign v$IN_2573_out0 = v$IN_3540_out0;
assign v$IN_2574_out0 = v$IN_3545_out0;
assign v$IN_2583_out0 = v$IN_3572_out0;
assign v$IN_2584_out0 = v$IN_3577_out0;
assign v$IN_3522_out0 = v$OUT_10237_out0;
assign v$IN_3554_out0 = v$OUT_10269_out0;
assign v$ANDOUT_4975_out0 = v$C_12847_out0;
assign v$ANDOUT_4976_out0 = v$C_12848_out0;
assign v$MUX3_2588_out0 = v$G6_3951_out0 ? v$ANDOUT_4975_out0 : v$ADDEROUT_2206_out0;
assign v$MUX3_2589_out0 = v$G6_3952_out0 ? v$ANDOUT_4976_out0 : v$ADDEROUT_2207_out0;
assign v$IN_3412_out0 = v$IN_3522_out0;
assign v$IN_3422_out0 = v$IN_3554_out0;
assign v$SEL1_5953_out0 = v$IN_2573_out0[23:1];
assign v$SEL1_5958_out0 = v$IN_2574_out0[23:1];
assign v$SEL1_5985_out0 = v$IN_2583_out0[23:1];
assign v$SEL1_5990_out0 = v$IN_2584_out0[23:1];
assign v$SEL1_10697_out0 = v$IN_2573_out0[22:0];
assign v$SEL1_10702_out0 = v$IN_2574_out0[22:0];
assign v$SEL1_10729_out0 = v$IN_2583_out0[22:0];
assign v$SEL1_10734_out0 = v$IN_2584_out0[22:0];
assign v$_2939_out0 = { v$C2_115_out0,v$SEL1_10697_out0 };
assign v$_2944_out0 = { v$C2_120_out0,v$SEL1_10702_out0 };
assign v$_2971_out0 = { v$C2_147_out0,v$SEL1_10729_out0 };
assign v$_2976_out0 = { v$C2_152_out0,v$SEL1_10734_out0 };
assign v$MUX4_3947_out0 = v$EQ1_1429_out0 ? v$OP2_5118_out0 : v$MUX3_2588_out0;
assign v$MUX4_3948_out0 = v$EQ1_1430_out0 ? v$OP2_5119_out0 : v$MUX3_2589_out0;
assign v$SEL1_5935_out0 = v$IN_3412_out0[23:8];
assign v$SEL1_5967_out0 = v$IN_3422_out0[23:8];
assign v$_6246_out0 = { v$SEL1_5953_out0,v$C1_3982_out0 };
assign v$_6251_out0 = { v$SEL1_5958_out0,v$C1_3987_out0 };
assign v$_6278_out0 = { v$SEL1_5985_out0,v$C1_4014_out0 };
assign v$_6283_out0 = { v$SEL1_5990_out0,v$C1_4019_out0 };
assign v$SEL1_10679_out0 = v$IN_3412_out0[15:0];
assign v$SEL1_10711_out0 = v$IN_3422_out0[15:0];
assign v$MUX1_1302_out0 = v$LEFT$SHIT_1814_out0 ? v$_2939_out0 : v$_6246_out0;
assign v$MUX1_1307_out0 = v$LEFT$SHIT_1819_out0 ? v$_2944_out0 : v$_6251_out0;
assign v$MUX1_1334_out0 = v$LEFT$SHIT_1846_out0 ? v$_2971_out0 : v$_6278_out0;
assign v$MUX1_1339_out0 = v$LEFT$SHIT_1851_out0 ? v$_2976_out0 : v$_6283_out0;
assign v$_2921_out0 = { v$C2_97_out0,v$SEL1_10679_out0 };
assign v$_2953_out0 = { v$C2_129_out0,v$SEL1_10711_out0 };
assign v$_6228_out0 = { v$SEL1_5935_out0,v$C1_3964_out0 };
assign v$_6260_out0 = { v$SEL1_5967_out0,v$C1_3996_out0 };
assign v$ALUOUT_12827_out0 = v$MUX4_3947_out0;
assign v$ALUOUT_12828_out0 = v$MUX4_3948_out0;
assign v$MUX1_1284_out0 = v$LEFT$SHIT_1796_out0 ? v$_2921_out0 : v$_6228_out0;
assign v$MUX1_1316_out0 = v$LEFT$SHIT_1828_out0 ? v$_2953_out0 : v$_6260_out0;
assign v$ALUOUT_4692_out0 = v$ALUOUT_12827_out0;
assign v$ALUOUT_4693_out0 = v$ALUOUT_12828_out0;
assign v$MUX2_13224_out0 = v$EN_3592_out0 ? v$MUX1_1302_out0 : v$IN_2573_out0;
assign v$MUX2_13225_out0 = v$EN_3593_out0 ? v$MUX1_1307_out0 : v$IN_2574_out0;
assign v$MUX2_13234_out0 = v$EN_3602_out0 ? v$MUX1_1334_out0 : v$IN_2583_out0;
assign v$MUX2_13235_out0 = v$EN_3603_out0 ? v$MUX1_1339_out0 : v$IN_2584_out0;
assign v$MUX4_42_out0 = v$IR2$15_5012_out0 ? v$ALUOUT_4692_out0 : v$REGDIN_11576_out0;
assign v$MUX4_43_out0 = v$IR2$15_5013_out0 ? v$ALUOUT_4693_out0 : v$REGDIN_11577_out0;
assign v$MUX2_1406_out0 = v$EN_562_out0 ? v$MUX1_1284_out0 : v$IN_3412_out0;
assign v$MUX2_1416_out0 = v$EN_572_out0 ? v$MUX1_1316_out0 : v$IN_3422_out0;
assign v$OUT_10253_out0 = v$MUX2_13224_out0;
assign v$OUT_10258_out0 = v$MUX2_13225_out0;
assign v$OUT_10285_out0 = v$MUX2_13234_out0;
assign v$OUT_10290_out0 = v$MUX2_13235_out0;
assign v$ALUOUT_11622_out0 = v$ALUOUT_4692_out0;
assign v$ALUOUT_11623_out0 = v$ALUOUT_4693_out0;
assign v$IN_3542_out0 = v$OUT_10253_out0;
assign v$IN_3547_out0 = v$OUT_10258_out0;
assign v$IN_3574_out0 = v$OUT_10285_out0;
assign v$IN_3579_out0 = v$OUT_10290_out0;
assign v$ALUOUT_6795_out0 = v$ALUOUT_11622_out0;
assign v$ALUOUT_6796_out0 = v$ALUOUT_11623_out0;
assign v$OUT_10235_out0 = v$MUX2_1406_out0;
assign v$OUT_10267_out0 = v$MUX2_1416_out0;
assign v$IN_3521_out0 = v$OUT_10235_out0;
assign v$IN_3553_out0 = v$OUT_10267_out0;
assign v$_6015_out0 = v$ALUOUT_6795_out0[15:15];
assign v$_6016_out0 = v$ALUOUT_6796_out0[15:15];
assign v$IN_7585_out0 = v$IN_3542_out0;
assign v$IN_7586_out0 = v$IN_3547_out0;
assign v$IN_7591_out0 = v$IN_3574_out0;
assign v$IN_7592_out0 = v$IN_3579_out0;
assign v$EQ1_11412_out0 = v$ALUOUT_6795_out0 == 16'h0;
assign v$EQ1_11413_out0 = v$ALUOUT_6796_out0 == 16'h0;
assign v$IN_3411_out0 = v$IN_3521_out0;
assign v$IN_3421_out0 = v$IN_3553_out0;
assign v$SEL1_5955_out0 = v$IN_7585_out0[23:2];
assign v$SEL1_5960_out0 = v$IN_7586_out0[23:2];
assign v$SEL1_5987_out0 = v$IN_7591_out0[23:2];
assign v$SEL1_5992_out0 = v$IN_7592_out0[23:2];
assign v$G18_9163_out0 = v$_6015_out0 && v$IR2$VALID_8838_out0;
assign v$G18_9164_out0 = v$_6016_out0 && v$IR2$VALID_8839_out0;
assign v$G17_9354_out0 = v$EQ1_11412_out0 && v$IR2$VALID_8838_out0;
assign v$G17_9355_out0 = v$EQ1_11413_out0 && v$IR2$VALID_8839_out0;
assign v$SEL1_10699_out0 = v$IN_7585_out0[21:0];
assign v$SEL1_10704_out0 = v$IN_7586_out0[21:0];
assign v$SEL1_10731_out0 = v$IN_7591_out0[21:0];
assign v$SEL1_10736_out0 = v$IN_7592_out0[21:0];
assign v$MUX3_665_out0 = v$G18_9163_out0 ? v$G18_9163_out0 : v$REG2_7598_out0;
assign v$MUX3_666_out0 = v$G18_9164_out0 ? v$G18_9164_out0 : v$REG2_7599_out0;
assign v$_2941_out0 = { v$C2_117_out0,v$SEL1_10699_out0 };
assign v$_2946_out0 = { v$C2_122_out0,v$SEL1_10704_out0 };
assign v$_2973_out0 = { v$C2_149_out0,v$SEL1_10731_out0 };
assign v$_2978_out0 = { v$C2_154_out0,v$SEL1_10736_out0 };
assign v$SEL1_5934_out0 = v$IN_3411_out0[23:16];
assign v$SEL1_5966_out0 = v$IN_3421_out0[23:16];
assign v$_6248_out0 = { v$SEL1_5955_out0,v$C1_3984_out0 };
assign v$_6253_out0 = { v$SEL1_5960_out0,v$C1_3989_out0 };
assign v$_6280_out0 = { v$SEL1_5987_out0,v$C1_4016_out0 };
assign v$_6285_out0 = { v$SEL1_5992_out0,v$C1_4021_out0 };
assign v$MUX4_8278_out0 = v$G17_9354_out0 ? v$G17_9354_out0 : v$REG3_12548_out0;
assign v$MUX4_8279_out0 = v$G17_9355_out0 ? v$G17_9355_out0 : v$REG3_12549_out0;
assign v$SEL1_10678_out0 = v$IN_3411_out0[7:0];
assign v$SEL1_10710_out0 = v$IN_3421_out0[7:0];
assign v$MUX1_1304_out0 = v$LEFT$SHIT_1816_out0 ? v$_2941_out0 : v$_6248_out0;
assign v$MUX1_1309_out0 = v$LEFT$SHIT_1821_out0 ? v$_2946_out0 : v$_6253_out0;
assign v$MUX1_1336_out0 = v$LEFT$SHIT_1848_out0 ? v$_2973_out0 : v$_6280_out0;
assign v$MUX1_1341_out0 = v$LEFT$SHIT_1853_out0 ? v$_2978_out0 : v$_6285_out0;
assign v$EQ_2421_out0 = v$MUX4_8278_out0;
assign v$EQ_2422_out0 = v$MUX4_8279_out0;
assign v$_2920_out0 = { v$C2_96_out0,v$SEL1_10678_out0 };
assign v$_2952_out0 = { v$C2_128_out0,v$SEL1_10710_out0 };
assign v$_6227_out0 = { v$SEL1_5934_out0,v$C1_3963_out0 };
assign v$_6259_out0 = { v$SEL1_5966_out0,v$C1_3995_out0 };
assign v$MI_7903_out0 = v$MUX3_665_out0;
assign v$MI_7904_out0 = v$MUX3_666_out0;
assign v$EQ_360_out0 = v$EQ_2421_out0;
assign v$EQ_361_out0 = v$EQ_2422_out0;
assign v$MUX1_1283_out0 = v$LEFT$SHIT_1795_out0 ? v$_2920_out0 : v$_6227_out0;
assign v$MUX1_1315_out0 = v$LEFT$SHIT_1827_out0 ? v$_2952_out0 : v$_6259_out0;
assign v$MUX2_1396_out0 = v$EN_5392_out0 ? v$MUX1_1304_out0 : v$IN_7585_out0;
assign v$MUX2_1397_out0 = v$EN_5393_out0 ? v$MUX1_1309_out0 : v$IN_7586_out0;
assign v$MUX2_1402_out0 = v$EN_5398_out0 ? v$MUX1_1336_out0 : v$IN_7591_out0;
assign v$MUX2_1403_out0 = v$EN_5399_out0 ? v$MUX1_1341_out0 : v$IN_7592_out0;
assign v$MI_4239_out0 = v$MI_7903_out0;
assign v$MI_4240_out0 = v$MI_7904_out0;
assign v$MI_1351_out0 = v$MI_4239_out0;
assign v$MI_1352_out0 = v$MI_4240_out0;
assign v$MUX2_1405_out0 = v$EN_561_out0 ? v$MUX1_1283_out0 : v$IN_3411_out0;
assign v$MUX2_1415_out0 = v$EN_571_out0 ? v$MUX1_1315_out0 : v$IN_3421_out0;
assign v$EQ_4165_out0 = v$EQ_360_out0;
assign v$EQ_4166_out0 = v$EQ_361_out0;
assign v$OUT_10255_out0 = v$MUX2_1396_out0;
assign v$OUT_10260_out0 = v$MUX2_1397_out0;
assign v$OUT_10287_out0 = v$MUX2_1402_out0;
assign v$OUT_10292_out0 = v$MUX2_1403_out0;
assign v$EQ_2185_out0 = v$EQ_4165_out0;
assign v$EQ_2186_out0 = v$EQ_4166_out0;
assign v$IN_3541_out0 = v$OUT_10255_out0;
assign v$IN_3546_out0 = v$OUT_10260_out0;
assign v$IN_3573_out0 = v$OUT_10287_out0;
assign v$IN_3578_out0 = v$OUT_10292_out0;
assign v$MI_5906_out0 = v$MI_1351_out0;
assign v$MI_5907_out0 = v$MI_1352_out0;
assign v$OUT_10234_out0 = v$MUX2_1405_out0;
assign v$OUT_10266_out0 = v$MUX2_1415_out0;
assign v$MUX1_7471_out0 = v$G2_12220_out0 ? v$C1_3093_out0 : v$OUT_10234_out0;
assign v$MUX1_7475_out0 = v$G2_12224_out0 ? v$C1_3097_out0 : v$OUT_10266_out0;
assign v$MI_8107_out0 = v$MI_5906_out0;
assign v$MI_8108_out0 = v$MI_5907_out0;
assign v$EQ_8992_out0 = v$EQ_2185_out0;
assign v$EQ_8993_out0 = v$EQ_2186_out0;
assign v$IN_10875_out0 = v$IN_3541_out0;
assign v$IN_10876_out0 = v$IN_3546_out0;
assign v$IN_10881_out0 = v$IN_3573_out0;
assign v$IN_10882_out0 = v$IN_3578_out0;
assign v$SEL1_5954_out0 = v$IN_10875_out0[23:4];
assign v$SEL1_5959_out0 = v$IN_10876_out0[23:4];
assign v$SEL1_5986_out0 = v$IN_10881_out0[23:4];
assign v$SEL1_5991_out0 = v$IN_10882_out0[23:4];
assign v$OUT_6726_out0 = v$MUX1_7471_out0;
assign v$OUT_6730_out0 = v$MUX1_7475_out0;
assign v$MI_7673_out0 = v$MI_8107_out0;
assign v$MI_7674_out0 = v$MI_8108_out0;
assign v$EQ_9954_out0 = v$EQ_8992_out0;
assign v$EQ_9955_out0 = v$EQ_8993_out0;
assign v$SEL1_10698_out0 = v$IN_10875_out0[19:0];
assign v$SEL1_10703_out0 = v$IN_10876_out0[19:0];
assign v$SEL1_10730_out0 = v$IN_10881_out0[19:0];
assign v$SEL1_10735_out0 = v$IN_10882_out0[19:0];
assign v$G20_1501_out0 = v$G22_10639_out0 || v$EQ_9954_out0;
assign v$G20_1502_out0 = v$G22_10640_out0 || v$EQ_9955_out0;
assign v$_2940_out0 = { v$C2_116_out0,v$SEL1_10698_out0 };
assign v$_2945_out0 = { v$C2_121_out0,v$SEL1_10703_out0 };
assign v$_2972_out0 = { v$C2_148_out0,v$SEL1_10730_out0 };
assign v$_2977_out0 = { v$C2_153_out0,v$SEL1_10735_out0 };
assign v$_6247_out0 = { v$SEL1_5954_out0,v$C1_3983_out0 };
assign v$_6252_out0 = { v$SEL1_5959_out0,v$C1_3988_out0 };
assign v$_6279_out0 = { v$SEL1_5986_out0,v$C1_4015_out0 };
assign v$_6284_out0 = { v$SEL1_5991_out0,v$C1_4020_out0 };
assign v$SEL6_6954_out0 = v$OUT_6726_out0[23:13];
assign v$SEL6_6955_out0 = v$OUT_6730_out0[23:13];
assign v$G25_8408_out0 = v$JEQ_869_out0 && v$EQ_9954_out0;
assign v$G25_8409_out0 = v$JEQ_870_out0 && v$EQ_9955_out0;
assign v$G19_9396_out0 = v$JMI_8762_out0 && v$MI_7673_out0;
assign v$G19_9397_out0 = v$JMI_8763_out0 && v$MI_7674_out0;
assign v$G24_386_out0 = v$JLS_11527_out0 && v$G20_1501_out0;
assign v$G24_387_out0 = v$JLS_11528_out0 && v$G20_1502_out0;
assign v$MUX1_1303_out0 = v$LEFT$SHIT_1815_out0 ? v$_2940_out0 : v$_6247_out0;
assign v$MUX1_1308_out0 = v$LEFT$SHIT_1820_out0 ? v$_2945_out0 : v$_6252_out0;
assign v$MUX1_1335_out0 = v$LEFT$SHIT_1847_out0 ? v$_2972_out0 : v$_6279_out0;
assign v$MUX1_1340_out0 = v$LEFT$SHIT_1852_out0 ? v$_2977_out0 : v$_6284_out0;
assign v$_9986_out0 = { v$C5_6_out0,v$SEL6_6954_out0 };
assign v$_9987_out0 = { v$C5_7_out0,v$SEL6_6955_out0 };
assign v$G21_10619_out0 = v$G19_9396_out0 || v$G25_8408_out0;
assign v$G21_10620_out0 = v$G19_9397_out0 || v$G25_8409_out0;
assign v$G15_3722_out0 = v$JMP_2998_out0 || v$G21_10619_out0;
assign v$G15_3723_out0 = v$JMP_2999_out0 || v$G21_10620_out0;
assign v$MUX2_10558_out0 = v$EN_3168_out0 ? v$MUX1_1303_out0 : v$IN_10875_out0;
assign v$MUX2_10559_out0 = v$EN_3169_out0 ? v$MUX1_1308_out0 : v$IN_10876_out0;
assign v$MUX2_10564_out0 = v$EN_3174_out0 ? v$MUX1_1335_out0 : v$IN_10881_out0;
assign v$MUX2_10565_out0 = v$EN_3175_out0 ? v$MUX1_1340_out0 : v$IN_10882_out0;
assign v$MUX4_12976_out0 = v$IS$32$BITS_2837_out0 ? v$OUT_6726_out0 : v$_9986_out0;
assign v$MUX4_12977_out0 = v$IS$32$BITS_2838_out0 ? v$OUT_6730_out0 : v$_9987_out0;
assign v$OP2_2852_out0 = v$MUX4_12976_out0;
assign v$OP2_2853_out0 = v$MUX4_12977_out0;
assign v$OUT_10254_out0 = v$MUX2_10558_out0;
assign v$OUT_10259_out0 = v$MUX2_10559_out0;
assign v$OUT_10286_out0 = v$MUX2_10564_out0;
assign v$OUT_10291_out0 = v$MUX2_10565_out0;
assign v$G23_12511_out0 = v$G15_3722_out0 || v$G17_3706_out0;
assign v$G23_12512_out0 = v$G15_3723_out0 || v$G17_3707_out0;
assign v$G16_544_out0 = v$G23_12511_out0 || v$G24_386_out0;
assign v$G16_545_out0 = v$G23_12512_out0 || v$G24_387_out0;
assign v$IN_3539_out0 = v$OUT_10254_out0;
assign v$IN_3544_out0 = v$OUT_10259_out0;
assign v$IN_3571_out0 = v$OUT_10286_out0;
assign v$IN_3576_out0 = v$OUT_10291_out0;
assign v$B_5834_out0 = v$OP2_2852_out0;
assign v$B_5835_out0 = v$OP2_2853_out0;
assign v$B_1106_out0 = v$B_5834_out0;
assign v$B_1107_out0 = v$B_5835_out0;
assign v$IN_3416_out0 = v$IN_3539_out0;
assign v$IN_3418_out0 = v$IN_3544_out0;
assign v$IN_3426_out0 = v$IN_3571_out0;
assign v$IN_3428_out0 = v$IN_3576_out0;
assign v$TAKEJUMP_7106_out0 = v$G16_544_out0;
assign v$TAKEJUMP_7107_out0 = v$G16_545_out0;
assign v$SEL7_491_out0 = v$B_1106_out0[0:0];
assign v$SEL7_492_out0 = v$B_1107_out0[0:0];
assign v$OP2_2372_out0 = v$B_1106_out0;
assign v$OP2_2373_out0 = v$B_1106_out0;
assign v$OP2_2374_out0 = v$B_1106_out0;
assign v$OP2_2375_out0 = v$B_1106_out0;
assign v$OP2_2376_out0 = v$B_1106_out0;
assign v$OP2_2377_out0 = v$B_1106_out0;
assign v$OP2_2378_out0 = v$B_1106_out0;
assign v$OP2_2379_out0 = v$B_1106_out0;
assign v$OP2_2380_out0 = v$B_1106_out0;
assign v$OP2_2381_out0 = v$B_1106_out0;
assign v$OP2_2382_out0 = v$B_1106_out0;
assign v$OP2_2383_out0 = v$B_1106_out0;
assign v$OP2_2384_out0 = v$B_1107_out0;
assign v$OP2_2385_out0 = v$B_1107_out0;
assign v$OP2_2386_out0 = v$B_1107_out0;
assign v$OP2_2387_out0 = v$B_1107_out0;
assign v$OP2_2388_out0 = v$B_1107_out0;
assign v$OP2_2389_out0 = v$B_1107_out0;
assign v$OP2_2390_out0 = v$B_1107_out0;
assign v$OP2_2391_out0 = v$B_1107_out0;
assign v$OP2_2392_out0 = v$B_1107_out0;
assign v$OP2_2393_out0 = v$B_1107_out0;
assign v$OP2_2394_out0 = v$B_1107_out0;
assign v$OP2_2395_out0 = v$B_1107_out0;
assign v$SEL1_5952_out0 = v$IN_3416_out0[23:8];
assign v$SEL1_5957_out0 = v$IN_3418_out0[23:8];
assign v$SEL1_5984_out0 = v$IN_3426_out0[23:8];
assign v$SEL1_5989_out0 = v$IN_3428_out0[23:8];
assign v$G26_9193_out0 = v$G29_5378_out0 || v$TAKEJUMP_7106_out0;
assign v$G26_9194_out0 = v$G29_5379_out0 || v$TAKEJUMP_7107_out0;
assign v$SEL1_10696_out0 = v$IN_3416_out0[15:0];
assign v$SEL1_10701_out0 = v$IN_3418_out0[15:0];
assign v$SEL1_10728_out0 = v$IN_3426_out0[15:0];
assign v$SEL1_10733_out0 = v$IN_3428_out0[15:0];
assign v$_2938_out0 = { v$C2_114_out0,v$SEL1_10696_out0 };
assign v$_2943_out0 = { v$C2_119_out0,v$SEL1_10701_out0 };
assign v$_2970_out0 = { v$C2_146_out0,v$SEL1_10728_out0 };
assign v$_2975_out0 = { v$C2_151_out0,v$SEL1_10733_out0 };
assign v$MUX3_5173_out0 = v$SEL7_491_out0 ? v$A_10147_out0 : v$C2_5340_out0;
assign v$MUX3_5174_out0 = v$SEL7_492_out0 ? v$A_10148_out0 : v$C2_5341_out0;
assign v$_6245_out0 = { v$SEL1_5952_out0,v$C1_3981_out0 };
assign v$_6250_out0 = { v$SEL1_5957_out0,v$C1_3986_out0 };
assign v$_6277_out0 = { v$SEL1_5984_out0,v$C1_4013_out0 };
assign v$_6282_out0 = { v$SEL1_5989_out0,v$C1_4018_out0 };
assign v$OP2_6911_out0 = v$OP2_2372_out0;
assign v$OP2_6912_out0 = v$OP2_2373_out0;
assign v$OP2_6913_out0 = v$OP2_2374_out0;
assign v$OP2_6914_out0 = v$OP2_2375_out0;
assign v$OP2_6915_out0 = v$OP2_2376_out0;
assign v$OP2_6916_out0 = v$OP2_2377_out0;
assign v$OP2_6917_out0 = v$OP2_2378_out0;
assign v$OP2_6918_out0 = v$OP2_2379_out0;
assign v$OP2_6919_out0 = v$OP2_2380_out0;
assign v$OP2_6920_out0 = v$OP2_2381_out0;
assign v$OP2_6921_out0 = v$OP2_2382_out0;
assign v$OP2_6922_out0 = v$OP2_2383_out0;
assign v$OP2_6923_out0 = v$OP2_2384_out0;
assign v$OP2_6924_out0 = v$OP2_2385_out0;
assign v$OP2_6925_out0 = v$OP2_2386_out0;
assign v$OP2_6926_out0 = v$OP2_2387_out0;
assign v$OP2_6927_out0 = v$OP2_2388_out0;
assign v$OP2_6928_out0 = v$OP2_2389_out0;
assign v$OP2_6929_out0 = v$OP2_2390_out0;
assign v$OP2_6930_out0 = v$OP2_2391_out0;
assign v$OP2_6931_out0 = v$OP2_2392_out0;
assign v$OP2_6932_out0 = v$OP2_2393_out0;
assign v$OP2_6933_out0 = v$OP2_2394_out0;
assign v$OP2_6934_out0 = v$OP2_2395_out0;
assign v$MUX8_8058_out0 = v$G26_9193_out0 ? v$MUX5_12042_out0 : v$PCINTERRUPT_12603_out0;
assign v$MUX8_8059_out0 = v$G26_9194_out0 ? v$MUX5_12043_out0 : v$PCINTERRUPT_12604_out0;
assign v$MUX1_1301_out0 = v$LEFT$SHIT_1813_out0 ? v$_2938_out0 : v$_6245_out0;
assign v$MUX1_1306_out0 = v$LEFT$SHIT_1818_out0 ? v$_2943_out0 : v$_6250_out0;
assign v$MUX1_1333_out0 = v$LEFT$SHIT_1845_out0 ? v$_2970_out0 : v$_6277_out0;
assign v$MUX1_1338_out0 = v$LEFT$SHIT_1850_out0 ? v$_2975_out0 : v$_6282_out0;
assign v$MUX2_2435_out0 = v$ININTERRUPT_433_out0 ? v$MUX8_8058_out0 : v$PCNORMAL_8422_out0;
assign v$MUX2_2436_out0 = v$ININTERRUPT_434_out0 ? v$MUX8_8059_out0 : v$PCNORMAL_8423_out0;
assign v$MUX1_5806_out0 = v$MULTIPLYING$BIT_1607_out0 ? v$OP2_6911_out0 : v$C5_2672_out0;
assign v$MUX1_5807_out0 = v$MULTIPLYING$BIT_1608_out0 ? v$OP2_6912_out0 : v$C5_2673_out0;
assign v$MUX1_5808_out0 = v$MULTIPLYING$BIT_1609_out0 ? v$OP2_6913_out0 : v$C5_2674_out0;
assign v$MUX1_5809_out0 = v$MULTIPLYING$BIT_1610_out0 ? v$OP2_6914_out0 : v$C5_2675_out0;
assign v$MUX1_5810_out0 = v$MULTIPLYING$BIT_1611_out0 ? v$OP2_6915_out0 : v$C5_2676_out0;
assign v$MUX1_5811_out0 = v$MULTIPLYING$BIT_1612_out0 ? v$OP2_6916_out0 : v$C5_2677_out0;
assign v$MUX1_5812_out0 = v$MULTIPLYING$BIT_1613_out0 ? v$OP2_6917_out0 : v$C5_2678_out0;
assign v$MUX1_5813_out0 = v$MULTIPLYING$BIT_1614_out0 ? v$OP2_6918_out0 : v$C5_2679_out0;
assign v$MUX1_5814_out0 = v$MULTIPLYING$BIT_1615_out0 ? v$OP2_6919_out0 : v$C5_2680_out0;
assign v$MUX1_5815_out0 = v$MULTIPLYING$BIT_1616_out0 ? v$OP2_6920_out0 : v$C5_2681_out0;
assign v$MUX1_5816_out0 = v$MULTIPLYING$BIT_1617_out0 ? v$OP2_6921_out0 : v$C5_2682_out0;
assign v$MUX1_5817_out0 = v$MULTIPLYING$BIT_1618_out0 ? v$OP2_6922_out0 : v$C5_2683_out0;
assign v$MUX1_5818_out0 = v$MULTIPLYING$BIT_1619_out0 ? v$OP2_6923_out0 : v$C5_2684_out0;
assign v$MUX1_5819_out0 = v$MULTIPLYING$BIT_1620_out0 ? v$OP2_6924_out0 : v$C5_2685_out0;
assign v$MUX1_5820_out0 = v$MULTIPLYING$BIT_1621_out0 ? v$OP2_6925_out0 : v$C5_2686_out0;
assign v$MUX1_5821_out0 = v$MULTIPLYING$BIT_1622_out0 ? v$OP2_6926_out0 : v$C5_2687_out0;
assign v$MUX1_5822_out0 = v$MULTIPLYING$BIT_1623_out0 ? v$OP2_6927_out0 : v$C5_2688_out0;
assign v$MUX1_5823_out0 = v$MULTIPLYING$BIT_1624_out0 ? v$OP2_6928_out0 : v$C5_2689_out0;
assign v$MUX1_5824_out0 = v$MULTIPLYING$BIT_1625_out0 ? v$OP2_6929_out0 : v$C5_2690_out0;
assign v$MUX1_5825_out0 = v$MULTIPLYING$BIT_1626_out0 ? v$OP2_6930_out0 : v$C5_2691_out0;
assign v$MUX1_5826_out0 = v$MULTIPLYING$BIT_1627_out0 ? v$OP2_6931_out0 : v$C5_2692_out0;
assign v$MUX1_5827_out0 = v$MULTIPLYING$BIT_1628_out0 ? v$OP2_6932_out0 : v$C5_2693_out0;
assign v$MUX1_5828_out0 = v$MULTIPLYING$BIT_1629_out0 ? v$OP2_6933_out0 : v$C5_2694_out0;
assign v$MUX1_5829_out0 = v$MULTIPLYING$BIT_1630_out0 ? v$OP2_6934_out0 : v$C5_2695_out0;
assign v$MUX2_12807_out0 = v$EXEC1_13169_out0 ? v$MUX3_5173_out0 : v$SEL6_3784_out0;
assign v$MUX2_12808_out0 = v$EXEC1_13170_out0 ? v$MUX3_5174_out0 : v$SEL6_3785_out0;
assign v$MUX4_781_out0 = v$TAKEJUMP_7106_out0 ? v$N_13005_out0 : v$MUX2_2435_out0;
assign v$MUX4_782_out0 = v$TAKEJUMP_7107_out0 ? v$N_13006_out0 : v$MUX2_2436_out0;
assign v$SEL5_783_out0 = v$MUX2_12807_out0[0:0];
assign v$SEL5_784_out0 = v$MUX2_12808_out0[0:0];
assign v$MUX2_1410_out0 = v$EN_566_out0 ? v$MUX1_1301_out0 : v$IN_3416_out0;
assign v$MUX2_1412_out0 = v$EN_568_out0 ? v$MUX1_1306_out0 : v$IN_3418_out0;
assign v$MUX2_1420_out0 = v$EN_576_out0 ? v$MUX1_1333_out0 : v$IN_3426_out0;
assign v$MUX2_1422_out0 = v$EN_578_out0 ? v$MUX1_1338_out0 : v$IN_3428_out0;
assign v$OP1_9574_out0 = v$MUX2_12807_out0;
assign v$OP1_9586_out0 = v$MUX2_12808_out0;
assign v$PC_1881_out0 = v$MUX4_781_out0;
assign v$PC_1882_out0 = v$MUX4_782_out0;
assign v$OP1_2074_out0 = v$OP1_9574_out0;
assign v$OP1_2086_out0 = v$OP1_9586_out0;
assign v$SUM$0_8097_out0 = v$SEL5_783_out0;
assign v$SUM$0_8098_out0 = v$SEL5_784_out0;
assign v$OUT_10252_out0 = v$MUX2_1410_out0;
assign v$OUT_10257_out0 = v$MUX2_1412_out0;
assign v$OUT_10284_out0 = v$MUX2_1420_out0;
assign v$OUT_10289_out0 = v$MUX2_1422_out0;
assign v$NEXTINSTRUCTIONADDRESS_13095_out0 = v$MUX4_781_out0;
assign v$NEXTINSTRUCTIONADDRESS_13096_out0 = v$MUX4_782_out0;
assign v$IN_3538_out0 = v$OUT_10252_out0;
assign v$IN_3543_out0 = v$OUT_10257_out0;
assign v$IN_3570_out0 = v$OUT_10284_out0;
assign v$IN_3575_out0 = v$OUT_10289_out0;
assign v$PCNEXT_4654_out0 = v$NEXTINSTRUCTIONADDRESS_13095_out0;
assign v$PCNEXT_4655_out0 = v$NEXTINSTRUCTIONADDRESS_13096_out0;
assign {v$A1_10168_out1,v$A1_10168_out0 } = v$PC_1881_out0 + v$C1_11144_out0 + v$EN_6318_out0;
assign {v$A1_10169_out1,v$A1_10169_out0 } = v$PC_1882_out0 + v$C1_11145_out0 + v$EN_6319_out0;
assign v$SEL8_12466_out0 = v$OP1_2074_out0[23:1];
assign v$SEL8_12478_out0 = v$OP1_2086_out0[23:1];
assign v$PC$NEXT0_1086_out0 = v$PCNEXT_4654_out0;
assign v$PC$NEXT1_2199_out0 = v$PCNEXT_4655_out0;
assign v$IN_3415_out0 = v$IN_3538_out0;
assign v$IN_3417_out0 = v$IN_3543_out0;
assign v$IN_3425_out0 = v$IN_3570_out0;
assign v$IN_3427_out0 = v$IN_3575_out0;
assign v$IGNORE_3653_out0 = v$A1_10168_out1;
assign v$IGNORE_3654_out0 = v$A1_10169_out1;
assign v$SUM_9219_out0 = v$A1_10168_out0;
assign v$SUM_9220_out0 = v$A1_10169_out0;
assign v$_12756_out0 = { v$SEL8_12466_out0,v$CIN_11850_out0 };
assign v$_12768_out0 = { v$SEL8_12478_out0,v$CIN_11862_out0 };
assign v$SEL1_5951_out0 = v$IN_3415_out0[23:16];
assign v$SEL1_5956_out0 = v$IN_3417_out0[23:16];
assign v$SEL1_5983_out0 = v$IN_3425_out0[23:16];
assign v$SEL1_5988_out0 = v$IN_3427_out0[23:16];
assign v$ADDRESS_10499_out0 = v$PC$NEXT0_1086_out0;
assign v$ADDRESS_10500_out0 = v$PC$NEXT1_2199_out0;
assign {v$A1_10524_out1,v$A1_10524_out0 } = v$_12756_out0 + v$MUX1_5807_out0 + v$C6_7385_out0;
assign {v$A1_10536_out1,v$A1_10536_out0 } = v$_12768_out0 + v$MUX1_5819_out0 + v$C6_7397_out0;
assign v$SEL1_10695_out0 = v$IN_3415_out0[7:0];
assign v$SEL1_10700_out0 = v$IN_3417_out0[7:0];
assign v$SEL1_10727_out0 = v$IN_3425_out0[7:0];
assign v$SEL1_10732_out0 = v$IN_3427_out0[7:0];
assign v$_2937_out0 = { v$C2_113_out0,v$SEL1_10695_out0 };
assign v$_2942_out0 = { v$C2_118_out0,v$SEL1_10700_out0 };
assign v$_2969_out0 = { v$C2_145_out0,v$SEL1_10727_out0 };
assign v$_2974_out0 = { v$C2_150_out0,v$SEL1_10732_out0 };
assign v$COUT_5614_out0 = v$A1_10524_out1;
assign v$COUT_5626_out0 = v$A1_10536_out1;
assign v$_6244_out0 = { v$SEL1_5951_out0,v$C1_3980_out0 };
assign v$_6249_out0 = { v$SEL1_5956_out0,v$C1_3985_out0 };
assign v$_6276_out0 = { v$SEL1_5983_out0,v$C1_4012_out0 };
assign v$_6281_out0 = { v$SEL1_5988_out0,v$C1_4017_out0 };
assign v$SUM_10460_out0 = v$A1_10524_out0;
assign v$SUM_10472_out0 = v$A1_10536_out0;
assign v$MUX1_1300_out0 = v$LEFT$SHIT_1812_out0 ? v$_2937_out0 : v$_6244_out0;
assign v$MUX1_1305_out0 = v$LEFT$SHIT_1817_out0 ? v$_2942_out0 : v$_6249_out0;
assign v$MUX1_1332_out0 = v$LEFT$SHIT_1844_out0 ? v$_2969_out0 : v$_6276_out0;
assign v$MUX1_1337_out0 = v$LEFT$SHIT_1849_out0 ? v$_2974_out0 : v$_6281_out0;
assign v$SUM_2162_out0 = v$SUM_10460_out0;
assign v$SUM_2174_out0 = v$SUM_10472_out0;
assign v$COUT_7043_out0 = v$COUT_5614_out0;
assign v$COUT_7055_out0 = v$COUT_5626_out0;
assign v$MUX2_1409_out0 = v$EN_565_out0 ? v$MUX1_1300_out0 : v$IN_3415_out0;
assign v$MUX2_1411_out0 = v$EN_567_out0 ? v$MUX1_1305_out0 : v$IN_3417_out0;
assign v$MUX2_1419_out0 = v$EN_575_out0 ? v$MUX1_1332_out0 : v$IN_3425_out0;
assign v$MUX2_1421_out0 = v$EN_577_out0 ? v$MUX1_1337_out0 : v$IN_3427_out0;
assign v$SEL1_2216_out0 = v$SUM_2162_out0[0:0];
assign v$SEL1_2217_out0 = v$SUM_2174_out0[0:0];
assign v$CIN_2601_out0 = v$COUT_7043_out0;
assign v$CIN_2613_out0 = v$COUT_7055_out0;
assign v$OP1_9580_out0 = v$SUM_2162_out0;
assign v$OP1_9592_out0 = v$SUM_2174_out0;
assign v$OP1_2080_out0 = v$OP1_9580_out0;
assign v$OP1_2092_out0 = v$OP1_9592_out0;
assign v$SUM$1_6901_out0 = v$SEL1_2216_out0;
assign v$SUM$1_6902_out0 = v$SEL1_2217_out0;
assign v$OUT_10251_out0 = v$MUX2_1409_out0;
assign v$OUT_10256_out0 = v$MUX2_1411_out0;
assign v$OUT_10283_out0 = v$MUX2_1419_out0;
assign v$OUT_10288_out0 = v$MUX2_1421_out0;
assign v$CIN_11856_out0 = v$CIN_2601_out0;
assign v$CIN_11868_out0 = v$CIN_2613_out0;
assign v$MUX1_7472_out0 = v$G2_12221_out0 ? v$C1_3094_out0 : v$OUT_10251_out0;
assign v$MUX1_7473_out0 = v$G2_12222_out0 ? v$C1_3095_out0 : v$OUT_10256_out0;
assign v$MUX1_7476_out0 = v$G2_12225_out0 ? v$C1_3098_out0 : v$OUT_10283_out0;
assign v$MUX1_7477_out0 = v$G2_12226_out0 ? v$C1_3099_out0 : v$OUT_10288_out0;
assign v$SEL8_12472_out0 = v$OP1_2080_out0[23:1];
assign v$SEL8_12484_out0 = v$OP1_2092_out0[23:1];
assign v$OUT_6727_out0 = v$MUX1_7472_out0;
assign v$OUT_6728_out0 = v$MUX1_7473_out0;
assign v$OUT_6731_out0 = v$MUX1_7476_out0;
assign v$OUT_6732_out0 = v$MUX1_7477_out0;
assign v$_12762_out0 = { v$SEL8_12472_out0,v$CIN_11856_out0 };
assign v$_12774_out0 = { v$SEL8_12484_out0,v$CIN_11868_out0 };
assign v$MUX4_3912_out0 = v$NEED$SHIFT$OP1_3226_out0 ? v$OUT_6728_out0 : v$OP1$MANTISA_7606_out0;
assign v$MUX4_3913_out0 = v$NEED$SHIFT$OP1_3227_out0 ? v$OUT_6732_out0 : v$OP1$MANTISA_7607_out0;
assign v$MUX1_9571_out0 = v$NEED$SHIFT$OP1_3226_out0 ? v$OP2$MANTISA_2212_out0 : v$OUT_6727_out0;
assign v$MUX1_9572_out0 = v$NEED$SHIFT$OP1_3227_out0 ? v$OP2$MANTISA_2213_out0 : v$OUT_6731_out0;
assign {v$A1_10530_out1,v$A1_10530_out0 } = v$_12762_out0 + v$MUX1_5813_out0 + v$C6_7391_out0;
assign {v$A1_10542_out1,v$A1_10542_out0 } = v$_12774_out0 + v$MUX1_5825_out0 + v$C6_7403_out0;
assign v$XOR2_5376_out0 = v$MUX1_9571_out0 ^ v$MUX3_2479_out0;
assign v$XOR2_5377_out0 = v$MUX1_9572_out0 ^ v$MUX3_2480_out0;
assign v$COUT_5620_out0 = v$A1_10530_out1;
assign v$COUT_5632_out0 = v$A1_10542_out1;
assign v$SUM_10466_out0 = v$A1_10530_out0;
assign v$SUM_10478_out0 = v$A1_10542_out0;
assign v$SUM_2168_out0 = v$SUM_10466_out0;
assign v$SUM_2180_out0 = v$SUM_10478_out0;
assign v$COUT_7049_out0 = v$COUT_5620_out0;
assign v$COUT_7061_out0 = v$COUT_5632_out0;
assign {v$A2_8371_out1,v$A2_8371_out0 } = v$MUX4_3912_out0 + v$XOR2_5376_out0 + v$IS$SUB_8690_out0;
assign {v$A2_8372_out1,v$A2_8372_out0 } = v$MUX4_3913_out0 + v$XOR2_5377_out0 + v$IS$SUB_8691_out0;
assign v$SUM_1056_out0 = v$A2_8371_out0;
assign v$SUM_1057_out0 = v$A2_8372_out0;
assign v$CIN_2603_out0 = v$COUT_7049_out0;
assign v$CIN_2615_out0 = v$COUT_7061_out0;
assign v$OP1_9582_out0 = v$SUM_2168_out0;
assign v$OP1_9594_out0 = v$SUM_2180_out0;
assign v$SEL1_9750_out0 = v$A2_8371_out0[23:1];
assign v$SEL1_9751_out0 = v$A2_8372_out0[23:1];
assign v$SEL2_9793_out0 = v$SUM_2168_out0[0:0];
assign v$SEL2_9794_out0 = v$SUM_2180_out0[0:0];
assign v$OVERFLOW_10307_out0 = v$A2_8371_out1;
assign v$OVERFLOW_10308_out0 = v$A2_8372_out1;
assign v$OVERFLOW_355_out0 = v$OVERFLOW_10307_out0;
assign v$OVERFLOW_356_out0 = v$OVERFLOW_10308_out0;
assign v$_735_out0 = { v$SEL1_9750_out0,v$C4_2467_out0 };
assign v$_736_out0 = { v$SEL1_9751_out0,v$C4_2468_out0 };
assign v$OP1_2082_out0 = v$OP1_9582_out0;
assign v$OP1_2094_out0 = v$OP1_9594_out0;
assign v$XOR1_3645_out0 = v$SUM_1056_out0 ^ v$C9_10581_out0;
assign v$XOR1_3646_out0 = v$SUM_1057_out0 ^ v$C9_10582_out0;
assign v$SUM$2_6320_out0 = v$SEL2_9793_out0;
assign v$SUM$2_6321_out0 = v$SEL2_9794_out0;
assign v$CIN_11858_out0 = v$CIN_2603_out0;
assign v$CIN_11870_out0 = v$CIN_2615_out0;
assign {v$A1_229_out1,v$A1_229_out0 } = v$XOR1_3645_out0 + v$C7_10012_out0 + v$C6_8186_out0;
assign {v$A1_230_out1,v$A1_230_out0 } = v$XOR1_3646_out0 + v$C7_10013_out0 + v$C6_8187_out0;
assign v$MUX7_1979_out0 = v$OVERFLOW_10307_out0 ? v$_735_out0 : v$SUM_1056_out0;
assign v$MUX7_1980_out0 = v$OVERFLOW_10308_out0 ? v$_736_out0 : v$SUM_1057_out0;
assign v$OVERFLOW_2338_out0 = v$OVERFLOW_355_out0;
assign v$OVERFLOW_2339_out0 = v$OVERFLOW_356_out0;
assign v$SEL8_12474_out0 = v$OP1_2082_out0[23:1];
assign v$SEL8_12486_out0 = v$OP1_2094_out0[23:1];
assign v$TWOS$COMPLEMENT$ADDER$COUT_2137_out0 = v$A1_229_out1;
assign v$TWOS$COMPLEMENT$ADDER$COUT_2138_out0 = v$A1_230_out1;
assign v$MUX5_4229_out0 = v$IS$A$LARGER_6990_out0 ? v$SUM_1056_out0 : v$A1_229_out0;
assign v$MUX5_4230_out0 = v$IS$A$LARGER_6991_out0 ? v$SUM_1057_out0 : v$A1_230_out0;
assign v$SEL3_9646_out0 = v$MUX7_1979_out0[22:0];
assign v$SEL3_9647_out0 = v$MUX7_1980_out0[22:0];
assign v$_12764_out0 = { v$SEL8_12474_out0,v$CIN_11858_out0 };
assign v$_12776_out0 = { v$SEL8_12486_out0,v$CIN_11870_out0 };
assign v$OVERFLOW_13127_out0 = v$OVERFLOW_2338_out0;
assign v$OVERFLOW_13128_out0 = v$OVERFLOW_2339_out0;
assign v$OVERFLOW_13177_out0 = v$OVERFLOW_2338_out0;
assign v$OVERFLOW_13178_out0 = v$OVERFLOW_2339_out0;
assign v$LZD$INPUT_6076_out0 = v$MUX5_4229_out0;
assign v$LZD$INPUT_6077_out0 = v$MUX5_4230_out0;
assign {v$A1_7602_out1,v$A1_7602_out0 } = v$C1_5006_out0 + v$EXPONENT_11194_out0 + v$OVERFLOW_13177_out0;
assign {v$A1_7603_out1,v$A1_7603_out0 } = v$C1_5007_out0 + v$EXPONENT_11195_out0 + v$OVERFLOW_13178_out0;
assign {v$A1_10532_out1,v$A1_10532_out0 } = v$_12764_out0 + v$MUX1_5815_out0 + v$C6_7393_out0;
assign {v$A1_10544_out1,v$A1_10544_out0 } = v$_12776_out0 + v$MUX1_5827_out0 + v$C6_7405_out0;
assign {v$A1_11001_out1,v$A1_11001_out0 } = v$C1_9390_out0 + v$EXPONENT_9232_out0 + v$OVERFLOW_13127_out0;
assign {v$A1_11002_out1,v$A1_11002_out0 } = v$C1_9391_out0 + v$EXPONENT_9233_out0 + v$OVERFLOW_13128_out0;
assign v$OUT_164_out0 = v$A1_7602_out0;
assign v$OUT_165_out0 = v$A1_7603_out0;
assign v$NOT$USED_1667_out0 = v$A1_7602_out1;
assign v$NOT$USED_1668_out0 = v$A1_7603_out1;
assign v$NOT$USED_3696_out0 = v$A1_11001_out1;
assign v$NOT$USED_3697_out0 = v$A1_11002_out1;
assign v$COUT_5622_out0 = v$A1_10532_out1;
assign v$COUT_5634_out0 = v$A1_10544_out1;
assign v$IN_8777_out0 = v$LZD$INPUT_6076_out0;
assign v$IN_8781_out0 = v$LZD$INPUT_6077_out0;
assign v$OUT_10129_out0 = v$A1_11001_out0;
assign v$OUT_10130_out0 = v$A1_11002_out0;
assign v$SUM_10468_out0 = v$A1_10532_out0;
assign v$SUM_10480_out0 = v$A1_10544_out0;
assign v$IN_12747_out0 = v$LZD$INPUT_6076_out0;
assign v$IN_12748_out0 = v$LZD$INPUT_6077_out0;
assign v$SEL1_282_out0 = v$IN_12747_out0[23:16];
assign v$SEL1_283_out0 = v$IN_12748_out0[23:16];
assign v$SUM_2170_out0 = v$SUM_10468_out0;
assign v$SUM_2182_out0 = v$SUM_10480_out0;
assign v$IN_3550_out0 = v$IN_8777_out0;
assign v$IN_3582_out0 = v$IN_8781_out0;
assign v$COUT_7051_out0 = v$COUT_5622_out0;
assign v$COUT_7063_out0 = v$COUT_5634_out0;
assign v$SEL2_12179_out0 = v$IN_12747_out0[15:8];
assign v$SEL2_12180_out0 = v$IN_12748_out0[15:8];
assign v$SEL1_12232_out0 = v$IN_12747_out0[7:0];
assign v$SEL1_12233_out0 = v$IN_12748_out0[7:0];
assign v$SEL3_887_out0 = v$SUM_2170_out0[0:0];
assign v$SEL3_888_out0 = v$SUM_2182_out0[0:0];
assign v$IN_2575_out0 = v$IN_3550_out0;
assign v$IN_2585_out0 = v$IN_3582_out0;
assign v$CIN_2604_out0 = v$COUT_7051_out0;
assign v$CIN_2616_out0 = v$COUT_7063_out0;
assign v$OP1_9583_out0 = v$SUM_2170_out0;
assign v$OP1_9595_out0 = v$SUM_2182_out0;
assign v$IN_10194_out0 = v$SEL1_282_out0;
assign v$IN_10195_out0 = v$SEL2_12179_out0;
assign v$IN_10196_out0 = v$SEL1_12232_out0;
assign v$IN_10197_out0 = v$SEL1_283_out0;
assign v$IN_10198_out0 = v$SEL2_12180_out0;
assign v$IN_10199_out0 = v$SEL1_12233_out0;
assign v$SEL2_1785_out0 = v$IN_10194_out0[7:4];
assign v$SEL2_1786_out0 = v$IN_10195_out0[7:4];
assign v$SEL2_1787_out0 = v$IN_10196_out0[7:4];
assign v$SEL2_1788_out0 = v$IN_10197_out0[7:4];
assign v$SEL2_1789_out0 = v$IN_10198_out0[7:4];
assign v$SEL2_1790_out0 = v$IN_10199_out0[7:4];
assign v$OP1_2083_out0 = v$OP1_9583_out0;
assign v$OP1_2095_out0 = v$OP1_9595_out0;
assign v$SUM$3_5420_out0 = v$SEL3_887_out0;
assign v$SUM$3_5421_out0 = v$SEL3_888_out0;
assign v$SEL1_5963_out0 = v$IN_2575_out0[23:1];
assign v$SEL1_5995_out0 = v$IN_2585_out0[23:1];
assign v$SEL1_10707_out0 = v$IN_2575_out0[22:0];
assign v$SEL1_10739_out0 = v$IN_2585_out0[22:0];
assign v$SEL1_11535_out0 = v$IN_10194_out0[3:0];
assign v$SEL1_11536_out0 = v$IN_10195_out0[3:0];
assign v$SEL1_11537_out0 = v$IN_10196_out0[3:0];
assign v$SEL1_11538_out0 = v$IN_10197_out0[3:0];
assign v$SEL1_11539_out0 = v$IN_10198_out0[3:0];
assign v$SEL1_11540_out0 = v$IN_10199_out0[3:0];
assign v$CIN_11859_out0 = v$CIN_2604_out0;
assign v$CIN_11871_out0 = v$CIN_2616_out0;
assign v$_2949_out0 = { v$C2_125_out0,v$SEL1_10707_out0 };
assign v$_2981_out0 = { v$C2_157_out0,v$SEL1_10739_out0 };
assign v$_6256_out0 = { v$SEL1_5963_out0,v$C1_3992_out0 };
assign v$_6288_out0 = { v$SEL1_5995_out0,v$C1_4024_out0 };
assign v$IN_10382_out0 = v$SEL1_11535_out0;
assign v$IN_10383_out0 = v$SEL2_1785_out0;
assign v$IN_10384_out0 = v$SEL1_11536_out0;
assign v$IN_10385_out0 = v$SEL2_1786_out0;
assign v$IN_10386_out0 = v$SEL1_11537_out0;
assign v$IN_10387_out0 = v$SEL2_1787_out0;
assign v$IN_10412_out0 = v$SEL1_11538_out0;
assign v$IN_10413_out0 = v$SEL2_1788_out0;
assign v$IN_10414_out0 = v$SEL1_11539_out0;
assign v$IN_10415_out0 = v$SEL2_1789_out0;
assign v$IN_10416_out0 = v$SEL1_11540_out0;
assign v$IN_10417_out0 = v$SEL2_1790_out0;
assign v$SEL8_12475_out0 = v$OP1_2083_out0[23:1];
assign v$SEL8_12487_out0 = v$OP1_2095_out0[23:1];
assign v$SEL3_1241_out0 = v$IN_10382_out0[2:2];
assign v$SEL3_1242_out0 = v$IN_10383_out0[2:2];
assign v$SEL3_1243_out0 = v$IN_10384_out0[2:2];
assign v$SEL3_1244_out0 = v$IN_10385_out0[2:2];
assign v$SEL3_1245_out0 = v$IN_10386_out0[2:2];
assign v$SEL3_1246_out0 = v$IN_10387_out0[2:2];
assign v$SEL3_1271_out0 = v$IN_10412_out0[2:2];
assign v$SEL3_1272_out0 = v$IN_10413_out0[2:2];
assign v$SEL3_1273_out0 = v$IN_10414_out0[2:2];
assign v$SEL3_1274_out0 = v$IN_10415_out0[2:2];
assign v$SEL3_1275_out0 = v$IN_10416_out0[2:2];
assign v$SEL3_1276_out0 = v$IN_10417_out0[2:2];
assign v$MUX1_1312_out0 = v$LEFT$SHIT_1824_out0 ? v$_2949_out0 : v$_6256_out0;
assign v$MUX1_1344_out0 = v$LEFT$SHIT_1856_out0 ? v$_2981_out0 : v$_6288_out0;
assign v$SEL4_4105_out0 = v$IN_10382_out0[3:3];
assign v$SEL4_4106_out0 = v$IN_10383_out0[3:3];
assign v$SEL4_4107_out0 = v$IN_10384_out0[3:3];
assign v$SEL4_4108_out0 = v$IN_10385_out0[3:3];
assign v$SEL4_4109_out0 = v$IN_10386_out0[3:3];
assign v$SEL4_4110_out0 = v$IN_10387_out0[3:3];
assign v$SEL4_4135_out0 = v$IN_10412_out0[3:3];
assign v$SEL4_4136_out0 = v$IN_10413_out0[3:3];
assign v$SEL4_4137_out0 = v$IN_10414_out0[3:3];
assign v$SEL4_4138_out0 = v$IN_10415_out0[3:3];
assign v$SEL4_4139_out0 = v$IN_10416_out0[3:3];
assign v$SEL4_4140_out0 = v$IN_10417_out0[3:3];
assign v$SEL2_5225_out0 = v$IN_10382_out0[1:1];
assign v$SEL2_5226_out0 = v$IN_10383_out0[1:1];
assign v$SEL2_5227_out0 = v$IN_10384_out0[1:1];
assign v$SEL2_5228_out0 = v$IN_10385_out0[1:1];
assign v$SEL2_5229_out0 = v$IN_10386_out0[1:1];
assign v$SEL2_5230_out0 = v$IN_10387_out0[1:1];
assign v$SEL2_5255_out0 = v$IN_10412_out0[1:1];
assign v$SEL2_5256_out0 = v$IN_10413_out0[1:1];
assign v$SEL2_5257_out0 = v$IN_10414_out0[1:1];
assign v$SEL2_5258_out0 = v$IN_10415_out0[1:1];
assign v$SEL2_5259_out0 = v$IN_10416_out0[1:1];
assign v$SEL2_5260_out0 = v$IN_10417_out0[1:1];
assign v$SEL1_9049_out0 = v$IN_10382_out0[0:0];
assign v$SEL1_9050_out0 = v$IN_10383_out0[0:0];
assign v$SEL1_9051_out0 = v$IN_10384_out0[0:0];
assign v$SEL1_9052_out0 = v$IN_10385_out0[0:0];
assign v$SEL1_9053_out0 = v$IN_10386_out0[0:0];
assign v$SEL1_9054_out0 = v$IN_10387_out0[0:0];
assign v$SEL1_9079_out0 = v$IN_10412_out0[0:0];
assign v$SEL1_9080_out0 = v$IN_10413_out0[0:0];
assign v$SEL1_9081_out0 = v$IN_10414_out0[0:0];
assign v$SEL1_9082_out0 = v$IN_10415_out0[0:0];
assign v$SEL1_9083_out0 = v$IN_10416_out0[0:0];
assign v$SEL1_9084_out0 = v$IN_10417_out0[0:0];
assign v$_12765_out0 = { v$SEL8_12475_out0,v$CIN_11859_out0 };
assign v$_12777_out0 = { v$SEL8_12487_out0,v$CIN_11871_out0 };
assign v$G10_629_out0 = !(v$SEL1_9049_out0 || v$SEL2_5225_out0);
assign v$G10_630_out0 = !(v$SEL1_9050_out0 || v$SEL2_5226_out0);
assign v$G10_631_out0 = !(v$SEL1_9051_out0 || v$SEL2_5227_out0);
assign v$G10_632_out0 = !(v$SEL1_9052_out0 || v$SEL2_5228_out0);
assign v$G10_633_out0 = !(v$SEL1_9053_out0 || v$SEL2_5229_out0);
assign v$G10_634_out0 = !(v$SEL1_9054_out0 || v$SEL2_5230_out0);
assign v$G10_659_out0 = !(v$SEL1_9079_out0 || v$SEL2_5255_out0);
assign v$G10_660_out0 = !(v$SEL1_9080_out0 || v$SEL2_5256_out0);
assign v$G10_661_out0 = !(v$SEL1_9081_out0 || v$SEL2_5257_out0);
assign v$G10_662_out0 = !(v$SEL1_9082_out0 || v$SEL2_5258_out0);
assign v$G10_663_out0 = !(v$SEL1_9083_out0 || v$SEL2_5259_out0);
assign v$G10_664_out0 = !(v$SEL1_9084_out0 || v$SEL2_5260_out0);
assign v$G6_2280_out0 = ! v$SEL2_5225_out0;
assign v$G6_2281_out0 = ! v$SEL2_5226_out0;
assign v$G6_2282_out0 = ! v$SEL2_5227_out0;
assign v$G6_2283_out0 = ! v$SEL2_5228_out0;
assign v$G6_2284_out0 = ! v$SEL2_5229_out0;
assign v$G6_2285_out0 = ! v$SEL2_5230_out0;
assign v$G6_2310_out0 = ! v$SEL2_5255_out0;
assign v$G6_2311_out0 = ! v$SEL2_5256_out0;
assign v$G6_2312_out0 = ! v$SEL2_5257_out0;
assign v$G6_2313_out0 = ! v$SEL2_5258_out0;
assign v$G6_2314_out0 = ! v$SEL2_5259_out0;
assign v$G6_2315_out0 = ! v$SEL2_5260_out0;
assign v$G5_3870_out0 = ! v$SEL4_4105_out0;
assign v$G5_3871_out0 = ! v$SEL4_4106_out0;
assign v$G5_3872_out0 = ! v$SEL4_4107_out0;
assign v$G5_3873_out0 = ! v$SEL4_4108_out0;
assign v$G5_3874_out0 = ! v$SEL4_4109_out0;
assign v$G5_3875_out0 = ! v$SEL4_4110_out0;
assign v$G5_3900_out0 = ! v$SEL4_4135_out0;
assign v$G5_3901_out0 = ! v$SEL4_4136_out0;
assign v$G5_3902_out0 = ! v$SEL4_4137_out0;
assign v$G5_3903_out0 = ! v$SEL4_4138_out0;
assign v$G5_3904_out0 = ! v$SEL4_4139_out0;
assign v$G5_3905_out0 = ! v$SEL4_4140_out0;
assign v$G11_6105_out0 = !(v$SEL3_1241_out0 || v$SEL4_4105_out0);
assign v$G11_6106_out0 = !(v$SEL3_1242_out0 || v$SEL4_4106_out0);
assign v$G11_6107_out0 = !(v$SEL3_1243_out0 || v$SEL4_4107_out0);
assign v$G11_6108_out0 = !(v$SEL3_1244_out0 || v$SEL4_4108_out0);
assign v$G11_6109_out0 = !(v$SEL3_1245_out0 || v$SEL4_4109_out0);
assign v$G11_6110_out0 = !(v$SEL3_1246_out0 || v$SEL4_4110_out0);
assign v$G11_6135_out0 = !(v$SEL3_1271_out0 || v$SEL4_4135_out0);
assign v$G11_6136_out0 = !(v$SEL3_1272_out0 || v$SEL4_4136_out0);
assign v$G11_6137_out0 = !(v$SEL3_1273_out0 || v$SEL4_4137_out0);
assign v$G11_6138_out0 = !(v$SEL3_1274_out0 || v$SEL4_4138_out0);
assign v$G11_6139_out0 = !(v$SEL3_1275_out0 || v$SEL4_4139_out0);
assign v$G11_6140_out0 = !(v$SEL3_1276_out0 || v$SEL4_4140_out0);
assign v$G8_7786_out0 = ! v$SEL3_1241_out0;
assign v$G8_7787_out0 = ! v$SEL3_1242_out0;
assign v$G8_7788_out0 = ! v$SEL3_1243_out0;
assign v$G8_7789_out0 = ! v$SEL3_1244_out0;
assign v$G8_7790_out0 = ! v$SEL3_1245_out0;
assign v$G8_7791_out0 = ! v$SEL3_1246_out0;
assign v$G8_7816_out0 = ! v$SEL3_1271_out0;
assign v$G8_7817_out0 = ! v$SEL3_1272_out0;
assign v$G8_7818_out0 = ! v$SEL3_1273_out0;
assign v$G8_7819_out0 = ! v$SEL3_1274_out0;
assign v$G8_7820_out0 = ! v$SEL3_1275_out0;
assign v$G8_7821_out0 = ! v$SEL3_1276_out0;
assign {v$A1_10533_out1,v$A1_10533_out0 } = v$_12765_out0 + v$MUX1_5816_out0 + v$C6_7394_out0;
assign {v$A1_10545_out1,v$A1_10545_out0 } = v$_12777_out0 + v$MUX1_5828_out0 + v$C6_7406_out0;
assign v$COUT_5623_out0 = v$A1_10533_out1;
assign v$COUT_5635_out0 = v$A1_10545_out1;
assign v$G3_8329_out0 = v$G10_629_out0 && v$G11_6105_out0;
assign v$G3_8330_out0 = v$G10_630_out0 && v$G11_6106_out0;
assign v$G3_8331_out0 = v$G10_631_out0 && v$G11_6107_out0;
assign v$G3_8332_out0 = v$G10_632_out0 && v$G11_6108_out0;
assign v$G3_8333_out0 = v$G10_633_out0 && v$G11_6109_out0;
assign v$G3_8334_out0 = v$G10_634_out0 && v$G11_6110_out0;
assign v$G3_8359_out0 = v$G10_659_out0 && v$G11_6135_out0;
assign v$G3_8360_out0 = v$G10_660_out0 && v$G11_6136_out0;
assign v$G3_8361_out0 = v$G10_661_out0 && v$G11_6137_out0;
assign v$G3_8362_out0 = v$G10_662_out0 && v$G11_6138_out0;
assign v$G3_8363_out0 = v$G10_663_out0 && v$G11_6139_out0;
assign v$G3_8364_out0 = v$G10_664_out0 && v$G11_6140_out0;
assign v$SUM_10469_out0 = v$A1_10533_out0;
assign v$SUM_10481_out0 = v$A1_10545_out0;
assign v$G9_12419_out0 = v$G8_7786_out0 && v$G5_3870_out0;
assign v$G9_12420_out0 = v$G8_7787_out0 && v$G5_3871_out0;
assign v$G9_12421_out0 = v$G8_7788_out0 && v$G5_3872_out0;
assign v$G9_12422_out0 = v$G8_7789_out0 && v$G5_3873_out0;
assign v$G9_12423_out0 = v$G8_7790_out0 && v$G5_3874_out0;
assign v$G9_12424_out0 = v$G8_7791_out0 && v$G5_3875_out0;
assign v$G9_12449_out0 = v$G8_7816_out0 && v$G5_3900_out0;
assign v$G9_12450_out0 = v$G8_7817_out0 && v$G5_3901_out0;
assign v$G9_12451_out0 = v$G8_7818_out0 && v$G5_3902_out0;
assign v$G9_12452_out0 = v$G8_7819_out0 && v$G5_3903_out0;
assign v$G9_12453_out0 = v$G8_7820_out0 && v$G5_3904_out0;
assign v$G9_12454_out0 = v$G8_7821_out0 && v$G5_3905_out0;
assign v$G7_12889_out0 = v$G6_2280_out0 || v$SEL3_1241_out0;
assign v$G7_12890_out0 = v$G6_2281_out0 || v$SEL3_1242_out0;
assign v$G7_12891_out0 = v$G6_2282_out0 || v$SEL3_1243_out0;
assign v$G7_12892_out0 = v$G6_2283_out0 || v$SEL3_1244_out0;
assign v$G7_12893_out0 = v$G6_2284_out0 || v$SEL3_1245_out0;
assign v$G7_12894_out0 = v$G6_2285_out0 || v$SEL3_1246_out0;
assign v$G7_12919_out0 = v$G6_2310_out0 || v$SEL3_1271_out0;
assign v$G7_12920_out0 = v$G6_2311_out0 || v$SEL3_1272_out0;
assign v$G7_12921_out0 = v$G6_2312_out0 || v$SEL3_1273_out0;
assign v$G7_12922_out0 = v$G6_2313_out0 || v$SEL3_1274_out0;
assign v$G7_12923_out0 = v$G6_2314_out0 || v$SEL3_1275_out0;
assign v$G7_12924_out0 = v$G6_2315_out0 || v$SEL3_1276_out0;
assign v$SUM_2171_out0 = v$SUM_10469_out0;
assign v$SUM_2183_out0 = v$SUM_10481_out0;
assign v$COUT_7052_out0 = v$COUT_5623_out0;
assign v$COUT_7064_out0 = v$COUT_5635_out0;
assign v$Z_8212_out0 = v$G3_8329_out0;
assign v$Z_8213_out0 = v$G3_8330_out0;
assign v$Z_8214_out0 = v$G3_8331_out0;
assign v$Z_8215_out0 = v$G3_8332_out0;
assign v$Z_8216_out0 = v$G3_8333_out0;
assign v$Z_8217_out0 = v$G3_8334_out0;
assign v$Z_8242_out0 = v$G3_8359_out0;
assign v$Z_8243_out0 = v$G3_8360_out0;
assign v$Z_8244_out0 = v$G3_8361_out0;
assign v$Z_8245_out0 = v$G3_8362_out0;
assign v$Z_8246_out0 = v$G3_8363_out0;
assign v$Z_8247_out0 = v$G3_8364_out0;
assign v$G4_12342_out0 = v$G7_12889_out0 && v$G5_3870_out0;
assign v$G4_12343_out0 = v$G7_12890_out0 && v$G5_3871_out0;
assign v$G4_12344_out0 = v$G7_12891_out0 && v$G5_3872_out0;
assign v$G4_12345_out0 = v$G7_12892_out0 && v$G5_3873_out0;
assign v$G4_12346_out0 = v$G7_12893_out0 && v$G5_3874_out0;
assign v$G4_12347_out0 = v$G7_12894_out0 && v$G5_3875_out0;
assign v$G4_12372_out0 = v$G7_12919_out0 && v$G5_3900_out0;
assign v$G4_12373_out0 = v$G7_12920_out0 && v$G5_3901_out0;
assign v$G4_12374_out0 = v$G7_12921_out0 && v$G5_3902_out0;
assign v$G4_12375_out0 = v$G7_12922_out0 && v$G5_3903_out0;
assign v$G4_12376_out0 = v$G7_12923_out0 && v$G5_3904_out0;
assign v$G4_12377_out0 = v$G7_12924_out0 && v$G5_3905_out0;
assign v$Z2_168_out0 = v$Z_8212_out0;
assign v$Z2_169_out0 = v$Z_8214_out0;
assign v$Z2_170_out0 = v$Z_8216_out0;
assign v$Z2_171_out0 = v$Z_8242_out0;
assign v$Z2_172_out0 = v$Z_8244_out0;
assign v$Z2_173_out0 = v$Z_8246_out0;
assign v$SEL4_475_out0 = v$SUM_2171_out0[0:0];
assign v$SEL4_476_out0 = v$SUM_2183_out0[0:0];
assign v$CIN_2605_out0 = v$COUT_7052_out0;
assign v$CIN_2617_out0 = v$COUT_7064_out0;
assign v$Z1_3792_out0 = v$Z_8213_out0;
assign v$Z1_3793_out0 = v$Z_8215_out0;
assign v$Z1_3794_out0 = v$Z_8217_out0;
assign v$Z1_3795_out0 = v$Z_8243_out0;
assign v$Z1_3796_out0 = v$Z_8245_out0;
assign v$Z1_3797_out0 = v$Z_8247_out0;
assign v$_4291_out0 = { v$G4_12342_out0,v$G9_12419_out0 };
assign v$_4292_out0 = { v$G4_12343_out0,v$G9_12420_out0 };
assign v$_4293_out0 = { v$G4_12344_out0,v$G9_12421_out0 };
assign v$_4294_out0 = { v$G4_12345_out0,v$G9_12422_out0 };
assign v$_4295_out0 = { v$G4_12346_out0,v$G9_12423_out0 };
assign v$_4296_out0 = { v$G4_12347_out0,v$G9_12424_out0 };
assign v$_4321_out0 = { v$G4_12372_out0,v$G9_12449_out0 };
assign v$_4322_out0 = { v$G4_12373_out0,v$G9_12450_out0 };
assign v$_4323_out0 = { v$G4_12374_out0,v$G9_12451_out0 };
assign v$_4324_out0 = { v$G4_12375_out0,v$G9_12452_out0 };
assign v$_4325_out0 = { v$G4_12376_out0,v$G9_12453_out0 };
assign v$_4326_out0 = { v$G4_12377_out0,v$G9_12454_out0 };
assign v$OP1_9584_out0 = v$SUM_2171_out0;
assign v$OP1_9596_out0 = v$SUM_2183_out0;
assign v$OP1_2084_out0 = v$OP1_9584_out0;
assign v$OP1_2096_out0 = v$OP1_9596_out0;
assign v$Y_4498_out0 = v$_4291_out0;
assign v$Y_4499_out0 = v$_4292_out0;
assign v$Y_4500_out0 = v$_4293_out0;
assign v$Y_4501_out0 = v$_4294_out0;
assign v$Y_4502_out0 = v$_4295_out0;
assign v$Y_4503_out0 = v$_4296_out0;
assign v$Y_4528_out0 = v$_4321_out0;
assign v$Y_4529_out0 = v$_4322_out0;
assign v$Y_4530_out0 = v$_4323_out0;
assign v$Y_4531_out0 = v$_4324_out0;
assign v$Y_4532_out0 = v$_4325_out0;
assign v$Y_4533_out0 = v$_4326_out0;
assign v$G1_9970_out0 = v$Z1_3792_out0 && v$Z2_168_out0;
assign v$G1_9971_out0 = v$Z1_3793_out0 && v$Z2_169_out0;
assign v$G1_9972_out0 = v$Z1_3794_out0 && v$Z2_170_out0;
assign v$G1_9973_out0 = v$Z1_3795_out0 && v$Z2_171_out0;
assign v$G1_9974_out0 = v$Z1_3796_out0 && v$Z2_172_out0;
assign v$G1_9975_out0 = v$Z1_3797_out0 && v$Z2_173_out0;
assign v$SUM$4_10567_out0 = v$SEL4_475_out0;
assign v$SUM$4_10568_out0 = v$SEL4_476_out0;
assign v$CIN_11860_out0 = v$CIN_2605_out0;
assign v$CIN_11872_out0 = v$CIN_2617_out0;
assign v$_3712_out0 = { v$Y_4499_out0,v$C1_12492_out0 };
assign v$_3713_out0 = { v$Y_4501_out0,v$C1_12493_out0 };
assign v$_3714_out0 = { v$Y_4503_out0,v$C1_12494_out0 };
assign v$_3715_out0 = { v$Y_4529_out0,v$C1_12495_out0 };
assign v$_3716_out0 = { v$Y_4531_out0,v$C1_12496_out0 };
assign v$_3717_out0 = { v$Y_4533_out0,v$C1_12497_out0 };
assign v$_5652_out0 = { v$Y_4498_out0,v$C2_5163_out0 };
assign v$_5653_out0 = { v$Y_4500_out0,v$C2_5164_out0 };
assign v$_5654_out0 = { v$Y_4502_out0,v$C2_5165_out0 };
assign v$_5655_out0 = { v$Y_4528_out0,v$C2_5166_out0 };
assign v$_5656_out0 = { v$Y_4530_out0,v$C2_5167_out0 };
assign v$_5657_out0 = { v$Y_4532_out0,v$C2_5168_out0 };
assign v$Z_6883_out0 = v$G1_9970_out0;
assign v$Z_6884_out0 = v$G1_9971_out0;
assign v$Z_6885_out0 = v$G1_9972_out0;
assign v$Z_6886_out0 = v$G1_9973_out0;
assign v$Z_6887_out0 = v$G1_9974_out0;
assign v$Z_6888_out0 = v$G1_9975_out0;
assign v$SEL8_12476_out0 = v$OP1_2084_out0[23:1];
assign v$SEL8_12488_out0 = v$OP1_2096_out0[23:1];
assign v$Z2_1177_out0 = v$Z_6884_out0;
assign v$Z2_1178_out0 = v$Z_6887_out0;
assign v$Z3_7758_out0 = v$Z_6883_out0;
assign v$Z3_7759_out0 = v$Z_6886_out0;
assign v$MUX1_10052_out0 = v$Z1_3792_out0 ? v$_5652_out0 : v$_3712_out0;
assign v$MUX1_10053_out0 = v$Z1_3793_out0 ? v$_5653_out0 : v$_3713_out0;
assign v$MUX1_10054_out0 = v$Z1_3794_out0 ? v$_5654_out0 : v$_3714_out0;
assign v$MUX1_10055_out0 = v$Z1_3795_out0 ? v$_5655_out0 : v$_3715_out0;
assign v$MUX1_10056_out0 = v$Z1_3796_out0 ? v$_5656_out0 : v$_3716_out0;
assign v$MUX1_10057_out0 = v$Z1_3797_out0 ? v$_5657_out0 : v$_3717_out0;
assign v$Z1_12534_out0 = v$Z_6885_out0;
assign v$Z1_12535_out0 = v$Z_6888_out0;
assign v$_12766_out0 = { v$SEL8_12476_out0,v$CIN_11860_out0 };
assign v$_12778_out0 = { v$SEL8_12488_out0,v$CIN_11872_out0 };
assign v$Y_5296_out0 = v$MUX1_10052_out0;
assign v$Y_5297_out0 = v$MUX1_10053_out0;
assign v$Y_5298_out0 = v$MUX1_10054_out0;
assign v$Y_5299_out0 = v$MUX1_10055_out0;
assign v$Y_5300_out0 = v$MUX1_10056_out0;
assign v$Y_5301_out0 = v$MUX1_10057_out0;
assign {v$A1_10534_out1,v$A1_10534_out0 } = v$_12766_out0 + v$MUX1_5817_out0 + v$C6_7395_out0;
assign {v$A1_10546_out1,v$A1_10546_out0 } = v$_12778_out0 + v$MUX1_5829_out0 + v$C6_7407_out0;
assign v$G2_11082_out0 = v$Z2_1177_out0 && v$Z3_7758_out0;
assign v$G2_11083_out0 = v$Z2_1178_out0 && v$Z3_7759_out0;
assign v$_555_out0 = { v$Y_5298_out0,v$C1_5267_out0 };
assign v$_556_out0 = { v$Y_5301_out0,v$C1_5268_out0 };
assign v$_1577_out0 = { v$Y_5297_out0,v$C2_8960_out0 };
assign v$_1578_out0 = { v$Y_5300_out0,v$C2_8961_out0 };
assign v$_2021_out0 = { v$Y_5296_out0,v$C4_11432_out0 };
assign v$_2022_out0 = { v$Y_5299_out0,v$C4_11433_out0 };
assign v$COUT_5624_out0 = v$A1_10534_out1;
assign v$COUT_5636_out0 = v$A1_10546_out1;
assign v$SUM_10470_out0 = v$A1_10534_out0;
assign v$SUM_10482_out0 = v$A1_10546_out0;
assign v$G1_12074_out0 = v$Z1_12534_out0 && v$G2_11082_out0;
assign v$G1_12075_out0 = v$Z1_12535_out0 && v$G2_11083_out0;
assign v$SUM_2172_out0 = v$SUM_10470_out0;
assign v$SUM_2184_out0 = v$SUM_10482_out0;
assign v$COUT_7053_out0 = v$COUT_5624_out0;
assign v$COUT_7065_out0 = v$COUT_5636_out0;
assign v$Z_9121_out0 = v$G1_12074_out0;
assign v$Z_9122_out0 = v$G1_12075_out0;
assign v$MUX1_10603_out0 = v$Z2_1177_out0 ? v$_555_out0 : v$_1577_out0;
assign v$MUX1_10604_out0 = v$Z2_1178_out0 ? v$_556_out0 : v$_1578_out0;
assign v$CIN_2602_out0 = v$COUT_7053_out0;
assign v$CIN_2614_out0 = v$COUT_7065_out0;
assign v$SEL9_3639_out0 = v$SUM_2172_out0[0:0];
assign v$SEL9_3640_out0 = v$SUM_2184_out0[0:0];
assign v$MUX2_9114_out0 = v$Z3_7758_out0 ? v$MUX1_10603_out0 : v$_2021_out0;
assign v$MUX2_9115_out0 = v$Z3_7759_out0 ? v$MUX1_10604_out0 : v$_2022_out0;
assign v$OP1_9581_out0 = v$SUM_2172_out0;
assign v$OP1_9593_out0 = v$SUM_2184_out0;
assign v$IS$SUM$0_10892_out0 = v$Z_9121_out0;
assign v$IS$SUM$0_10893_out0 = v$Z_9122_out0;
assign v$OP1_2081_out0 = v$OP1_9581_out0;
assign v$OP1_2093_out0 = v$OP1_9593_out0;
assign v$SUM$5_5344_out0 = v$SEL9_3639_out0;
assign v$SUM$5_5345_out0 = v$SEL9_3640_out0;
assign v$OUT_6175_out0 = v$MUX2_9114_out0;
assign v$OUT_6176_out0 = v$MUX2_9115_out0;
assign v$IS$SUM$0_10944_out0 = v$IS$SUM$0_10892_out0;
assign v$IS$SUM$0_10945_out0 = v$IS$SUM$0_10893_out0;
assign v$CIN_11857_out0 = v$CIN_2602_out0;
assign v$CIN_11869_out0 = v$CIN_2614_out0;
assign v$IS$SUM$0_402_out0 = v$IS$SUM$0_10944_out0;
assign v$IS$SUM$0_403_out0 = v$IS$SUM$0_10945_out0;
assign v$_6907_out0 = { v$OUT_6175_out0,v$C10_9110_out0 };
assign v$_6908_out0 = { v$OUT_6176_out0,v$C10_9111_out0 };
assign v$SEL8_12473_out0 = v$OP1_2081_out0[23:1];
assign v$SEL8_12485_out0 = v$OP1_2093_out0[23:1];
assign v$NORMALIZATION$SHIFT_1957_out0 = v$_6907_out0;
assign v$NORMALIZATION$SHIFT_1958_out0 = v$_6908_out0;
assign v$_12763_out0 = { v$SEL8_12473_out0,v$CIN_11857_out0 };
assign v$_12775_out0 = { v$SEL8_12485_out0,v$CIN_11869_out0 };
assign v$NORMALIZATION$SHIFT_459_out0 = v$NORMALIZATION$SHIFT_1957_out0;
assign v$NORMALIZATION$SHIFT_460_out0 = v$NORMALIZATION$SHIFT_1958_out0;
assign v$SHIFT$AMOUNT_4983_out0 = v$NORMALIZATION$SHIFT_1957_out0;
assign v$SHIFT$AMOUNT_4987_out0 = v$NORMALIZATION$SHIFT_1958_out0;
assign {v$A1_10531_out1,v$A1_10531_out0 } = v$_12763_out0 + v$MUX1_5814_out0 + v$C6_7392_out0;
assign {v$A1_10543_out1,v$A1_10543_out0 } = v$_12775_out0 + v$MUX1_5826_out0 + v$C6_7404_out0;
assign v$SEL3_440_out0 = v$SHIFT$AMOUNT_4983_out0[2:2];
assign v$SEL3_444_out0 = v$SHIFT$AMOUNT_4987_out0[2:2];
assign v$SEL1_1194_out0 = v$SHIFT$AMOUNT_4983_out0[0:0];
assign v$SEL1_1198_out0 = v$SHIFT$AMOUNT_4987_out0[0:0];
assign v$SEL4_3333_out0 = v$SHIFT$AMOUNT_4983_out0[3:3];
assign v$SEL4_3337_out0 = v$SHIFT$AMOUNT_4987_out0[3:3];
assign v$SEL7_4360_out0 = v$SHIFT$AMOUNT_4983_out0[5:5];
assign v$SEL7_4364_out0 = v$SHIFT$AMOUNT_4987_out0[5:5];
assign v$COUT_5621_out0 = v$A1_10531_out1;
assign v$COUT_5633_out0 = v$A1_10543_out1;
assign v$SEL5_7991_out0 = v$SHIFT$AMOUNT_4983_out0[4:4];
assign v$SEL5_7995_out0 = v$SHIFT$AMOUNT_4987_out0[4:4];
assign v$SEL6_9307_out0 = v$SHIFT$AMOUNT_4983_out0[6:6];
assign v$SEL6_9311_out0 = v$SHIFT$AMOUNT_4987_out0[6:6];
assign v$SUM_10467_out0 = v$A1_10531_out0;
assign v$SUM_10479_out0 = v$A1_10543_out0;
assign v$SEL8_11649_out0 = v$SHIFT$AMOUNT_4983_out0[7:7];
assign v$SEL8_11653_out0 = v$SHIFT$AMOUNT_4987_out0[7:7];
assign v$SEL2_13059_out0 = v$SHIFT$AMOUNT_4983_out0[1:1];
assign v$SEL2_13063_out0 = v$SHIFT$AMOUNT_4987_out0[1:1];
assign v$NORMALIZATION$SHIFT_13257_out0 = v$NORMALIZATION$SHIFT_459_out0;
assign v$NORMALIZATION$SHIFT_13258_out0 = v$NORMALIZATION$SHIFT_460_out0;
assign v$EN_569_out0 = v$SEL5_7991_out0;
assign v$EN_570_out0 = v$SEL4_3333_out0;
assign v$EN_579_out0 = v$SEL5_7995_out0;
assign v$EN_580_out0 = v$SEL4_3337_out0;
assign v$SUM_2169_out0 = v$SUM_10467_out0;
assign v$SUM_2181_out0 = v$SUM_10479_out0;
assign v$EN_3170_out0 = v$SEL3_440_out0;
assign v$EN_3176_out0 = v$SEL3_444_out0;
assign v$EN_3594_out0 = v$SEL1_1194_out0;
assign v$EN_3604_out0 = v$SEL1_1198_out0;
assign v$EN_5394_out0 = v$SEL2_13059_out0;
assign v$EN_5400_out0 = v$SEL2_13063_out0;
assign v$SEL14_6339_out0 = v$NORMALIZATION$SHIFT_13257_out0[4:0];
assign v$SEL14_6340_out0 = v$NORMALIZATION$SHIFT_13258_out0[4:0];
assign v$COUT_7050_out0 = v$COUT_5621_out0;
assign v$COUT_7062_out0 = v$COUT_5633_out0;
assign v$NORMALIZATION$SHIFT_7068_out0 = v$NORMALIZATION$SHIFT_13257_out0;
assign v$NORMALIZATION$SHIFT_7069_out0 = v$NORMALIZATION$SHIFT_13258_out0;
assign v$G1_11212_out0 = v$SEL7_4360_out0 || v$SEL6_9307_out0;
assign v$G1_11216_out0 = v$SEL7_4364_out0 || v$SEL6_9311_out0;
assign v$SEL10_989_out0 = v$SUM_2169_out0[0:0];
assign v$SEL10_990_out0 = v$SUM_2181_out0[0:0];
assign v$CIN_2600_out0 = v$COUT_7050_out0;
assign v$CIN_2612_out0 = v$COUT_7062_out0;
assign v$NORMALIZATION$SHIFT_3052_out0 = v$SEL14_6339_out0;
assign v$NORMALIZATION$SHIFT_3053_out0 = v$SEL14_6340_out0;
assign v$OP1_9579_out0 = v$SUM_2169_out0;
assign v$OP1_9591_out0 = v$SUM_2181_out0;
assign v$XOR1_9935_out0 = v$NORMALIZATION$SHIFT_7068_out0 ^ v$C1_767_out0;
assign v$XOR1_9936_out0 = v$NORMALIZATION$SHIFT_7069_out0 ^ v$C1_768_out0;
assign v$G2_12223_out0 = v$G1_11212_out0 || v$SEL8_11649_out0;
assign v$G2_12227_out0 = v$G1_11216_out0 || v$SEL8_11653_out0;
assign v$MUX2_13226_out0 = v$EN_3594_out0 ? v$MUX1_1312_out0 : v$IN_2575_out0;
assign v$MUX2_13236_out0 = v$EN_3604_out0 ? v$MUX1_1344_out0 : v$IN_2585_out0;
assign {v$A1_362_out1,v$A1_362_out0 } = v$EXPONENT_583_out0 + v$XOR1_9935_out0 + v$C2_1736_out0;
assign {v$A1_363_out1,v$A1_363_out0 } = v$EXPONENT_584_out0 + v$XOR1_9936_out0 + v$C2_1737_out0;
assign v$OP1_2079_out0 = v$OP1_9579_out0;
assign v$OP1_2091_out0 = v$OP1_9591_out0;
assign v$XOR1_7199_out0 = v$NORMALIZATION$SHIFT_3052_out0 ^ v$C1_10982_out0;
assign v$XOR1_7200_out0 = v$NORMALIZATION$SHIFT_3053_out0 ^ v$C1_10983_out0;
assign v$SUM$6_8556_out0 = v$SEL10_989_out0;
assign v$SUM$6_8557_out0 = v$SEL10_990_out0;
assign v$OUT_10263_out0 = v$MUX2_13226_out0;
assign v$OUT_10295_out0 = v$MUX2_13236_out0;
assign v$CIN_11855_out0 = v$CIN_2600_out0;
assign v$CIN_11867_out0 = v$CIN_2612_out0;
assign v$IN_3552_out0 = v$OUT_10263_out0;
assign v$IN_3584_out0 = v$OUT_10295_out0;
assign {v$A1_5275_out1,v$A1_5275_out0 } = v$EXPONENT_11500_out0 + v$XOR1_7199_out0 + v$C2_693_out0;
assign {v$A1_5276_out1,v$A1_5276_out0 } = v$EXPONENT_11501_out0 + v$XOR1_7200_out0 + v$C2_694_out0;
assign v$IGNORE_7524_out0 = v$A1_362_out1;
assign v$IGNORE_7525_out0 = v$A1_363_out1;
assign v$OUT_11281_out0 = v$A1_362_out0;
assign v$OUT_11282_out0 = v$A1_363_out0;
assign v$SEL8_12471_out0 = v$OP1_2079_out0[23:1];
assign v$SEL8_12483_out0 = v$OP1_2091_out0[23:1];
assign v$OUT_4211_out0 = v$A1_5275_out0;
assign v$OUT_4212_out0 = v$A1_5276_out0;
assign v$IN_7587_out0 = v$IN_3552_out0;
assign v$IN_7593_out0 = v$IN_3584_out0;
assign v$IGNORE_11642_out0 = v$A1_5275_out1;
assign v$IGNORE_11643_out0 = v$A1_5276_out1;
assign v$_12761_out0 = { v$SEL8_12471_out0,v$CIN_11855_out0 };
assign v$_12773_out0 = { v$SEL8_12483_out0,v$CIN_11867_out0 };
assign v$SEL1_5965_out0 = v$IN_7587_out0[23:2];
assign v$SEL1_5997_out0 = v$IN_7593_out0[23:2];
assign {v$A1_10529_out1,v$A1_10529_out0 } = v$_12761_out0 + v$MUX1_5812_out0 + v$C6_7390_out0;
assign {v$A1_10541_out1,v$A1_10541_out0 } = v$_12773_out0 + v$MUX1_5824_out0 + v$C6_7402_out0;
assign v$SEL1_10709_out0 = v$IN_7587_out0[21:0];
assign v$SEL1_10741_out0 = v$IN_7593_out0[21:0];
assign v$_2951_out0 = { v$C2_127_out0,v$SEL1_10709_out0 };
assign v$_2983_out0 = { v$C2_159_out0,v$SEL1_10741_out0 };
assign v$COUT_5619_out0 = v$A1_10529_out1;
assign v$COUT_5631_out0 = v$A1_10541_out1;
assign v$_6258_out0 = { v$SEL1_5965_out0,v$C1_3994_out0 };
assign v$_6290_out0 = { v$SEL1_5997_out0,v$C1_4026_out0 };
assign v$SUM_10465_out0 = v$A1_10529_out0;
assign v$SUM_10477_out0 = v$A1_10541_out0;
assign v$MUX1_1314_out0 = v$LEFT$SHIT_1826_out0 ? v$_2951_out0 : v$_6258_out0;
assign v$MUX1_1346_out0 = v$LEFT$SHIT_1858_out0 ? v$_2983_out0 : v$_6290_out0;
assign v$SUM_2167_out0 = v$SUM_10465_out0;
assign v$SUM_2179_out0 = v$SUM_10477_out0;
assign v$COUT_7048_out0 = v$COUT_5619_out0;
assign v$COUT_7060_out0 = v$COUT_5631_out0;
assign v$SEL11_729_out0 = v$SUM_2167_out0[0:0];
assign v$SEL11_730_out0 = v$SUM_2179_out0[0:0];
assign v$MUX2_1398_out0 = v$EN_5394_out0 ? v$MUX1_1314_out0 : v$IN_7587_out0;
assign v$MUX2_1404_out0 = v$EN_5400_out0 ? v$MUX1_1346_out0 : v$IN_7593_out0;
assign v$CIN_2596_out0 = v$COUT_7048_out0;
assign v$CIN_2608_out0 = v$COUT_7060_out0;
assign v$OP1_9575_out0 = v$SUM_2167_out0;
assign v$OP1_9587_out0 = v$SUM_2179_out0;
assign v$OP1_2075_out0 = v$OP1_9575_out0;
assign v$OP1_2087_out0 = v$OP1_9587_out0;
assign v$SUM$7_5287_out0 = v$SEL11_729_out0;
assign v$SUM$7_5288_out0 = v$SEL11_730_out0;
assign v$OUT_10265_out0 = v$MUX2_1398_out0;
assign v$OUT_10297_out0 = v$MUX2_1404_out0;
assign v$CIN_11851_out0 = v$CIN_2596_out0;
assign v$CIN_11863_out0 = v$CIN_2608_out0;
assign v$IN_3551_out0 = v$OUT_10265_out0;
assign v$IN_3583_out0 = v$OUT_10297_out0;
assign v$SEL8_12467_out0 = v$OP1_2075_out0[23:1];
assign v$SEL8_12479_out0 = v$OP1_2087_out0[23:1];
assign v$IN_10877_out0 = v$IN_3551_out0;
assign v$IN_10883_out0 = v$IN_3583_out0;
assign v$_12757_out0 = { v$SEL8_12467_out0,v$CIN_11851_out0 };
assign v$_12769_out0 = { v$SEL8_12479_out0,v$CIN_11863_out0 };
assign v$SEL1_5964_out0 = v$IN_10877_out0[23:4];
assign v$SEL1_5996_out0 = v$IN_10883_out0[23:4];
assign {v$A1_10525_out1,v$A1_10525_out0 } = v$_12757_out0 + v$MUX1_5808_out0 + v$C6_7386_out0;
assign {v$A1_10537_out1,v$A1_10537_out0 } = v$_12769_out0 + v$MUX1_5820_out0 + v$C6_7398_out0;
assign v$SEL1_10708_out0 = v$IN_10877_out0[19:0];
assign v$SEL1_10740_out0 = v$IN_10883_out0[19:0];
assign v$_2950_out0 = { v$C2_126_out0,v$SEL1_10708_out0 };
assign v$_2982_out0 = { v$C2_158_out0,v$SEL1_10740_out0 };
assign v$COUT_5615_out0 = v$A1_10525_out1;
assign v$COUT_5627_out0 = v$A1_10537_out1;
assign v$_6257_out0 = { v$SEL1_5964_out0,v$C1_3993_out0 };
assign v$_6289_out0 = { v$SEL1_5996_out0,v$C1_4025_out0 };
assign v$SUM_10461_out0 = v$A1_10525_out0;
assign v$SUM_10473_out0 = v$A1_10537_out0;
assign v$MUX1_1313_out0 = v$LEFT$SHIT_1825_out0 ? v$_2950_out0 : v$_6257_out0;
assign v$MUX1_1345_out0 = v$LEFT$SHIT_1857_out0 ? v$_2982_out0 : v$_6289_out0;
assign v$SUM_2163_out0 = v$SUM_10461_out0;
assign v$SUM_2175_out0 = v$SUM_10473_out0;
assign v$COUT_7044_out0 = v$COUT_5615_out0;
assign v$COUT_7056_out0 = v$COUT_5627_out0;
assign v$COUT$HALF_70_out0 = v$COUT_7044_out0;
assign v$COUT$HALF_71_out0 = v$COUT_7056_out0;
assign v$SUM$HALF_1659_out0 = v$SUM_2163_out0;
assign v$SUM$HALF_1660_out0 = v$SUM_2175_out0;
assign v$SEL13_2590_out0 = v$SUM_2163_out0[0:0];
assign v$SEL13_2591_out0 = v$SUM_2175_out0[0:0];
assign v$MUX2_10560_out0 = v$EN_3170_out0 ? v$MUX1_1313_out0 : v$IN_10877_out0;
assign v$MUX2_10566_out0 = v$EN_3176_out0 ? v$MUX1_1345_out0 : v$IN_10883_out0;
assign v$CIN_2598_out0 = v$COUT$HALF_70_out0;
assign v$CIN_2610_out0 = v$COUT$HALF_71_out0;
assign v$OP1_9577_out0 = v$SUM$HALF_1659_out0;
assign v$OP1_9589_out0 = v$SUM$HALF_1660_out0;
assign v$OUT_10264_out0 = v$MUX2_10560_out0;
assign v$OUT_10296_out0 = v$MUX2_10566_out0;
assign v$SUM$8_11009_out0 = v$SEL13_2590_out0;
assign v$SUM$8_11010_out0 = v$SEL13_2591_out0;
assign v$OP1_2077_out0 = v$OP1_9577_out0;
assign v$OP1_2089_out0 = v$OP1_9589_out0;
assign v$IN_3549_out0 = v$OUT_10264_out0;
assign v$IN_3581_out0 = v$OUT_10296_out0;
assign v$CIN_11853_out0 = v$CIN_2598_out0;
assign v$CIN_11865_out0 = v$CIN_2610_out0;
assign v$IN_3420_out0 = v$IN_3549_out0;
assign v$IN_3430_out0 = v$IN_3581_out0;
assign v$SEL8_12469_out0 = v$OP1_2077_out0[23:1];
assign v$SEL8_12481_out0 = v$OP1_2089_out0[23:1];
assign v$SEL1_5962_out0 = v$IN_3420_out0[23:8];
assign v$SEL1_5994_out0 = v$IN_3430_out0[23:8];
assign v$SEL1_10706_out0 = v$IN_3420_out0[15:0];
assign v$SEL1_10738_out0 = v$IN_3430_out0[15:0];
assign v$_12759_out0 = { v$SEL8_12469_out0,v$CIN_11853_out0 };
assign v$_12771_out0 = { v$SEL8_12481_out0,v$CIN_11865_out0 };
assign v$_2948_out0 = { v$C2_124_out0,v$SEL1_10706_out0 };
assign v$_2980_out0 = { v$C2_156_out0,v$SEL1_10738_out0 };
assign v$_6255_out0 = { v$SEL1_5962_out0,v$C1_3991_out0 };
assign v$_6287_out0 = { v$SEL1_5994_out0,v$C1_4023_out0 };
assign {v$A1_10527_out1,v$A1_10527_out0 } = v$_12759_out0 + v$MUX1_5810_out0 + v$C6_7388_out0;
assign {v$A1_10539_out1,v$A1_10539_out0 } = v$_12771_out0 + v$MUX1_5822_out0 + v$C6_7400_out0;
assign v$MUX1_1311_out0 = v$LEFT$SHIT_1823_out0 ? v$_2948_out0 : v$_6255_out0;
assign v$MUX1_1343_out0 = v$LEFT$SHIT_1855_out0 ? v$_2980_out0 : v$_6287_out0;
assign v$COUT_5617_out0 = v$A1_10527_out1;
assign v$COUT_5629_out0 = v$A1_10539_out1;
assign v$SUM_10463_out0 = v$A1_10527_out0;
assign v$SUM_10475_out0 = v$A1_10539_out0;
assign v$MUX2_1414_out0 = v$EN_570_out0 ? v$MUX1_1311_out0 : v$IN_3420_out0;
assign v$MUX2_1424_out0 = v$EN_580_out0 ? v$MUX1_1343_out0 : v$IN_3430_out0;
assign v$SUM_2165_out0 = v$SUM_10463_out0;
assign v$SUM_2177_out0 = v$SUM_10475_out0;
assign v$COUT_7046_out0 = v$COUT_5617_out0;
assign v$COUT_7058_out0 = v$COUT_5629_out0;
assign v$SEL12_741_out0 = v$SUM_2165_out0[0:0];
assign v$SEL12_742_out0 = v$SUM_2177_out0[0:0];
assign v$CIN_2597_out0 = v$COUT_7046_out0;
assign v$CIN_2609_out0 = v$COUT_7058_out0;
assign v$OP1_9576_out0 = v$SUM_2165_out0;
assign v$OP1_9588_out0 = v$SUM_2177_out0;
assign v$OUT_10262_out0 = v$MUX2_1414_out0;
assign v$OUT_10294_out0 = v$MUX2_1424_out0;
assign v$SUM$9_184_out0 = v$SEL12_741_out0;
assign v$SUM$9_185_out0 = v$SEL12_742_out0;
assign v$OP1_2076_out0 = v$OP1_9576_out0;
assign v$OP1_2088_out0 = v$OP1_9588_out0;
assign v$IN_3548_out0 = v$OUT_10262_out0;
assign v$IN_3580_out0 = v$OUT_10294_out0;
assign v$CIN_11852_out0 = v$CIN_2597_out0;
assign v$CIN_11864_out0 = v$CIN_2609_out0;
assign v$IN_3419_out0 = v$IN_3548_out0;
assign v$IN_3429_out0 = v$IN_3580_out0;
assign v$SEL8_12468_out0 = v$OP1_2076_out0[23:1];
assign v$SEL8_12480_out0 = v$OP1_2088_out0[23:1];
assign v$SEL1_5961_out0 = v$IN_3419_out0[23:16];
assign v$SEL1_5993_out0 = v$IN_3429_out0[23:16];
assign v$SEL1_10705_out0 = v$IN_3419_out0[7:0];
assign v$SEL1_10737_out0 = v$IN_3429_out0[7:0];
assign v$_12758_out0 = { v$SEL8_12468_out0,v$CIN_11852_out0 };
assign v$_12770_out0 = { v$SEL8_12480_out0,v$CIN_11864_out0 };
assign v$_2947_out0 = { v$C2_123_out0,v$SEL1_10705_out0 };
assign v$_2979_out0 = { v$C2_155_out0,v$SEL1_10737_out0 };
assign v$_6254_out0 = { v$SEL1_5961_out0,v$C1_3990_out0 };
assign v$_6286_out0 = { v$SEL1_5993_out0,v$C1_4022_out0 };
assign {v$A1_10526_out1,v$A1_10526_out0 } = v$_12758_out0 + v$MUX1_5809_out0 + v$C6_7387_out0;
assign {v$A1_10538_out1,v$A1_10538_out0 } = v$_12770_out0 + v$MUX1_5821_out0 + v$C6_7399_out0;
assign v$MUX1_1310_out0 = v$LEFT$SHIT_1822_out0 ? v$_2947_out0 : v$_6254_out0;
assign v$MUX1_1342_out0 = v$LEFT$SHIT_1854_out0 ? v$_2979_out0 : v$_6286_out0;
assign v$COUT_5616_out0 = v$A1_10526_out1;
assign v$COUT_5628_out0 = v$A1_10538_out1;
assign v$SUM_10462_out0 = v$A1_10526_out0;
assign v$SUM_10474_out0 = v$A1_10538_out0;
assign v$MUX2_1413_out0 = v$EN_569_out0 ? v$MUX1_1310_out0 : v$IN_3419_out0;
assign v$MUX2_1423_out0 = v$EN_579_out0 ? v$MUX1_1342_out0 : v$IN_3429_out0;
assign v$SUM_2164_out0 = v$SUM_10462_out0;
assign v$SUM_2176_out0 = v$SUM_10474_out0;
assign v$COUT_7045_out0 = v$COUT_5616_out0;
assign v$COUT_7057_out0 = v$COUT_5628_out0;
assign v$CIN_2599_out0 = v$COUT_7045_out0;
assign v$CIN_2611_out0 = v$COUT_7057_out0;
assign v$SEL14_3219_out0 = v$SUM_2164_out0[0:0];
assign v$SEL14_3220_out0 = v$SUM_2176_out0[0:0];
assign v$OP1_9578_out0 = v$SUM_2164_out0;
assign v$OP1_9590_out0 = v$SUM_2176_out0;
assign v$OUT_10261_out0 = v$MUX2_1413_out0;
assign v$OUT_10293_out0 = v$MUX2_1423_out0;
assign v$OP1_2078_out0 = v$OP1_9578_out0;
assign v$OP1_2090_out0 = v$OP1_9590_out0;
assign v$MUX1_7474_out0 = v$G2_12223_out0 ? v$C1_3096_out0 : v$OUT_10261_out0;
assign v$MUX1_7478_out0 = v$G2_12227_out0 ? v$C1_3100_out0 : v$OUT_10293_out0;
assign v$SUM$10_9699_out0 = v$SEL14_3219_out0;
assign v$SUM$10_9700_out0 = v$SEL14_3220_out0;
assign v$CIN_11854_out0 = v$CIN_2599_out0;
assign v$CIN_11866_out0 = v$CIN_2611_out0;
assign v$OUT_6729_out0 = v$MUX1_7474_out0;
assign v$OUT_6733_out0 = v$MUX1_7478_out0;
assign v$SEL8_12470_out0 = v$OP1_2078_out0[23:1];
assign v$SEL8_12482_out0 = v$OP1_2090_out0[23:1];
assign v$SEL2_4035_out0 = v$OUT_6729_out0[22:0];
assign v$SEL2_4036_out0 = v$OUT_6733_out0[22:0];
assign v$_12760_out0 = { v$SEL8_12470_out0,v$CIN_11854_out0 };
assign v$_12772_out0 = { v$SEL8_12482_out0,v$CIN_11866_out0 };
assign v$MUX2_1734_out0 = v$IS$SUM$0_10892_out0 ? v$C5_10888_out0 : v$SEL2_4035_out0;
assign v$MUX2_1735_out0 = v$IS$SUM$0_10893_out0 ? v$C5_10889_out0 : v$SEL2_4036_out0;
assign {v$A1_10528_out1,v$A1_10528_out0 } = v$_12760_out0 + v$MUX1_5811_out0 + v$C6_7389_out0;
assign {v$A1_10540_out1,v$A1_10540_out0 } = v$_12772_out0 + v$MUX1_5823_out0 + v$C6_7401_out0;
assign v$COUT_5618_out0 = v$A1_10528_out1;
assign v$COUT_5630_out0 = v$A1_10540_out1;
assign v$MUX6_8424_out0 = v$IS$SUB_8690_out0 ? v$MUX2_1734_out0 : v$SEL3_9646_out0;
assign v$MUX6_8425_out0 = v$IS$SUB_8691_out0 ? v$MUX2_1735_out0 : v$SEL3_9647_out0;
assign v$SUM_10464_out0 = v$A1_10528_out0;
assign v$SUM_10476_out0 = v$A1_10540_out0;
assign v$SUM_2166_out0 = v$SUM_10464_out0;
assign v$SUM_2178_out0 = v$SUM_10476_out0;
assign v$OUT1_6958_out0 = v$MUX6_8424_out0;
assign v$OUT1_6959_out0 = v$MUX6_8425_out0;
assign v$COUT_7047_out0 = v$COUT_5618_out0;
assign v$COUT_7059_out0 = v$COUT_5630_out0;
assign v$SUM_396_out0 = v$SUM_2166_out0;
assign v$SUM_397_out0 = v$SUM_2178_out0;
assign v$CIN_2594_out0 = v$COUT_7047_out0;
assign v$CIN_2606_out0 = v$COUT_7059_out0;
assign v$COUT_3407_out0 = v$COUT_7047_out0;
assign v$COUT_3408_out0 = v$COUT_7059_out0;
assign v$MANTISA$RESULT_4552_out0 = v$OUT1_6958_out0;
assign v$MANTISA$RESULT_4553_out0 = v$OUT1_6959_out0;
assign v$SEL15_6433_out0 = v$SUM_2166_out0[0:0];
assign v$SEL15_6434_out0 = v$SUM_2178_out0[0:0];
assign v$OP1_9573_out0 = v$SUM_2166_out0;
assign v$OP1_9585_out0 = v$SUM_2178_out0;
assign v$SEL10_1921_out0 = v$MANTISA$RESULT_4552_out0[22:13];
assign v$SEL10_1922_out0 = v$MANTISA$RESULT_4553_out0[22:13];
assign v$SEL7_1973_out0 = v$MANTISA$RESULT_4552_out0[22:13];
assign v$SEL7_1974_out0 = v$MANTISA$RESULT_4553_out0[22:13];
assign v$OP1_2073_out0 = v$OP1_9573_out0;
assign v$OP1_2085_out0 = v$OP1_9585_out0;
assign v$_4780_out0 = { v$MANTISA$RESULT_4552_out0,v$OUT_10129_out0 };
assign v$_4781_out0 = { v$MANTISA$RESULT_4553_out0,v$OUT_10130_out0 };
assign v$_6994_out0 = { v$SUM_396_out0,v$COUT_3407_out0 };
assign v$_6995_out0 = { v$SUM_397_out0,v$COUT_3408_out0 };
assign v$_10647_out0 = { v$MANTISA$RESULT_4552_out0,v$OUT_11281_out0 };
assign v$_10648_out0 = { v$MANTISA$RESULT_4553_out0,v$OUT_11282_out0 };
assign v$CIN_11849_out0 = v$CIN_2594_out0;
assign v$CIN_11861_out0 = v$CIN_2606_out0;
assign v$SUM$11_12086_out0 = v$SEL15_6433_out0;
assign v$SUM$11_12087_out0 = v$SEL15_6434_out0;
assign v$_3302_out0 = { v$SUM$11_12086_out0,v$_6994_out0 };
assign v$_3303_out0 = { v$SUM$11_12087_out0,v$_6995_out0 };
assign v$_7424_out0 = { v$SEL10_1921_out0,v$OUT_4211_out0 };
assign v$_7425_out0 = { v$SEL10_1922_out0,v$OUT_4212_out0 };
assign v$_10451_out0 = { v$SEL7_1973_out0,v$OUT_164_out0 };
assign v$_10452_out0 = { v$SEL7_1974_out0,v$OUT_165_out0 };
assign v$SEL8_12465_out0 = v$OP1_2073_out0[23:1];
assign v$SEL8_12477_out0 = v$OP1_2085_out0[23:1];
assign v$_52_out0 = { v$C9_1999_out0,v$_7424_out0 };
assign v$_53_out0 = { v$C9_2000_out0,v$_7425_out0 };
assign v$_7631_out0 = { v$C7_893_out0,v$_10451_out0 };
assign v$_7632_out0 = { v$C7_894_out0,v$_10452_out0 };
assign v$_9388_out0 = { v$SUM$10_9699_out0,v$_3302_out0 };
assign v$_9389_out0 = { v$SUM$10_9700_out0,v$_3303_out0 };
assign v$_12755_out0 = { v$SEL8_12465_out0,v$CIN_11849_out0 };
assign v$_12767_out0 = { v$SEL8_12477_out0,v$CIN_11861_out0 };
assign v$_6742_out0 = { v$SUM$9_184_out0,v$_9388_out0 };
assign v$_6743_out0 = { v$SUM$9_185_out0,v$_9389_out0 };
assign v$MUX12_10443_out0 = v$IS$32$BIT_7152_out0 ? v$_4780_out0 : v$_7631_out0;
assign v$MUX12_10444_out0 = v$IS$32$BIT_7153_out0 ? v$_4781_out0 : v$_7632_out0;
assign {v$A1_10523_out1,v$A1_10523_out0 } = v$_12755_out0 + v$MUX1_5806_out0 + v$C6_7384_out0;
assign {v$A1_10535_out1,v$A1_10535_out0 } = v$_12767_out0 + v$MUX1_5818_out0 + v$C6_7396_out0;
assign v$MUX6_12238_out0 = v$IS$32$BIT_7152_out0 ? v$_10647_out0 : v$_52_out0;
assign v$MUX6_12239_out0 = v$IS$32$BIT_7153_out0 ? v$_10648_out0 : v$_53_out0;
assign v$COUT_5613_out0 = v$A1_10523_out1;
assign v$COUT_5625_out0 = v$A1_10535_out1;
assign v$_10424_out0 = { v$SUM$8_11009_out0,v$_6742_out0 };
assign v$_10425_out0 = { v$SUM$8_11010_out0,v$_6743_out0 };
assign v$SUM_10459_out0 = v$A1_10523_out0;
assign v$SUM_10471_out0 = v$A1_10535_out0;
assign v$_11586_out0 = { v$MUX12_10443_out0,v$SEL13_12388_out0 };
assign v$_11587_out0 = { v$MUX12_10444_out0,v$SEL13_12389_out0 };
assign v$_11836_out0 = { v$MUX6_12238_out0,v$SUBTRACTION$SIGN_7667_out0 };
assign v$_11837_out0 = { v$MUX6_12239_out0,v$SUBTRACTION$SIGN_7668_out0 };
assign v$_1113_out0 = { v$SUM$7_5287_out0,v$_10424_out0 };
assign v$_1114_out0 = { v$SUM$7_5288_out0,v$_10425_out0 };
assign v$SUM_2161_out0 = v$SUM_10459_out0;
assign v$SUM_2173_out0 = v$SUM_10471_out0;
assign v$COUT_7042_out0 = v$COUT_5613_out0;
assign v$COUT_7054_out0 = v$COUT_5625_out0;
assign v$MUX1_9125_out0 = v$IS$SUB_3087_out0 ? v$_11836_out0 : v$_11586_out0;
assign v$MUX1_9126_out0 = v$IS$SUB_3088_out0 ? v$_11837_out0 : v$_11587_out0;
assign v$COUT$EXEC1_796_out0 = v$COUT_7042_out0;
assign v$COUT$EXEC1_797_out0 = v$COUT_7054_out0;
assign v$MUX7_3262_out0 = v$IS$SUM$0_402_out0 ? v$C5_2811_out0 : v$MUX1_9125_out0;
assign v$MUX7_3263_out0 = v$IS$SUM$0_403_out0 ? v$C5_2812_out0 : v$MUX1_9126_out0;
assign v$_8292_out0 = { v$SUM$6_8556_out0,v$_1113_out0 };
assign v$_8293_out0 = { v$SUM$6_8557_out0,v$_1114_out0 };
assign v$SUM$EXEC1_13195_out0 = v$SUM_2161_out0;
assign v$SUM$EXEC1_13196_out0 = v$SUM_2173_out0;
assign v$_3734_out0 = { v$SUM$5_5344_out0,v$_8292_out0 };
assign v$_3735_out0 = { v$SUM$5_5345_out0,v$_8293_out0 };
assign v$OUT1_12605_out0 = v$MUX7_3262_out0;
assign v$OUT1_12606_out0 = v$MUX7_3263_out0;
assign v$_12837_out0 = { v$SUM$11_12086_out0,v$SUM$EXEC1_13195_out0 };
assign v$_12838_out0 = { v$SUM$11_12087_out0,v$SUM$EXEC1_13196_out0 };
assign v$_6479_out0 = { v$SUM$4_10567_out0,v$_3734_out0 };
assign v$_6480_out0 = { v$SUM$4_10568_out0,v$_3735_out0 };
assign v$_7574_out0 = { v$SUM$10_9699_out0,v$_12837_out0 };
assign v$_7575_out0 = { v$SUM$10_9700_out0,v$_12838_out0 };
assign v$MUX2_11385_out0 = v$G2_2437_out0 ? v$OUT1_12605_out0 : v$C4_9419_out0;
assign v$MUX2_11386_out0 = v$G2_2438_out0 ? v$OUT1_12606_out0 : v$C4_9420_out0;
assign v$_5159_out0 = { v$SUM$9_184_out0,v$_7574_out0 };
assign v$_5160_out0 = { v$SUM$9_185_out0,v$_7575_out0 };
assign v$_11582_out0 = { v$SUM$3_5420_out0,v$_6479_out0 };
assign v$_11583_out0 = { v$SUM$3_5421_out0,v$_6480_out0 };
assign v$_2847_out0 = { v$SUM$8_11009_out0,v$_5159_out0 };
assign v$_2848_out0 = { v$SUM$8_11010_out0,v$_5160_out0 };
assign v$_11454_out0 = { v$SUM$2_6320_out0,v$_11582_out0 };
assign v$_11455_out0 = { v$SUM$2_6321_out0,v$_11583_out0 };
assign v$_8889_out0 = { v$SUM$1_6901_out0,v$_11454_out0 };
assign v$_8890_out0 = { v$SUM$1_6902_out0,v$_11455_out0 };
assign v$_11466_out0 = { v$SUM$7_5287_out0,v$_2847_out0 };
assign v$_11467_out0 = { v$SUM$7_5288_out0,v$_2848_out0 };
assign v$_1441_out0 = { v$SEL8_8402_out0,v$_8889_out0 };
assign v$_1442_out0 = { v$SEL8_8403_out0,v$_8890_out0 };
assign v$_12212_out0 = { v$SUM$6_8556_out0,v$_11466_out0 };
assign v$_12213_out0 = { v$SUM$6_8557_out0,v$_11467_out0 };
assign v$OUT_5704_out0 = v$_1441_out0;
assign v$OUT_5705_out0 = v$_1442_out0;
assign v$_5743_out0 = { v$SUM$5_5344_out0,v$_12212_out0 };
assign v$_5744_out0 = { v$SUM$5_5345_out0,v$_12213_out0 };
assign v$MULTIPLIER$OUT_6372_out0 = v$OUT_5704_out0;
assign v$MULTIPLIER$OUT_6373_out0 = v$OUT_5705_out0;
assign v$_11279_out0 = { v$SUM$4_10567_out0,v$_5743_out0 };
assign v$_11280_out0 = { v$SUM$4_10568_out0,v$_5744_out0 };
assign v$IN_7304_out0 = v$MULTIPLIER$OUT_6372_out0;
assign v$IN_7305_out0 = v$MULTIPLIER$OUT_6372_out0;
assign v$IN_7306_out0 = v$MULTIPLIER$OUT_6373_out0;
assign v$IN_7307_out0 = v$MULTIPLIER$OUT_6373_out0;
assign v$_8624_out0 = { v$SUM$3_5420_out0,v$_11279_out0 };
assign v$_8625_out0 = { v$SUM$3_5421_out0,v$_11280_out0 };
assign v$IN_7482_out0 = v$IN_7304_out0;
assign v$IN_7483_out0 = v$IN_7305_out0;
assign v$IN_7484_out0 = v$IN_7306_out0;
assign v$IN_7485_out0 = v$IN_7307_out0;
assign v$_11078_out0 = { v$SUM$2_6320_out0,v$_8624_out0 };
assign v$_11079_out0 = { v$SUM$2_6321_out0,v$_8625_out0 };
assign v$_1003_out0 = { v$SUM$1_6901_out0,v$_11078_out0 };
assign v$_1004_out0 = { v$SUM$1_6902_out0,v$_11079_out0 };
assign v$IN_5768_out0 = v$IN_7482_out0;
assign v$IN_5769_out0 = v$IN_7483_out0;
assign v$IN_5770_out0 = v$IN_7484_out0;
assign v$IN_5771_out0 = v$IN_7485_out0;
assign v$IN_9131_out0 = v$IN_7482_out0;
assign v$IN_9135_out0 = v$IN_7483_out0;
assign v$IN_9139_out0 = v$IN_7484_out0;
assign v$IN_9143_out0 = v$IN_7485_out0;
assign v$IN_12982_out0 = v$IN_7482_out0;
assign v$IN_12983_out0 = v$IN_7483_out0;
assign v$IN_12984_out0 = v$IN_7484_out0;
assign v$IN_12985_out0 = v$IN_7485_out0;
assign v$_809_out0 = { v$SUM$0_8097_out0,v$_1003_out0 };
assign v$_810_out0 = { v$SUM$0_8098_out0,v$_1004_out0 };
assign v$IN_2880_out0 = v$IN_5768_out0;
assign v$IN_2881_out0 = v$IN_5769_out0;
assign v$IN_2882_out0 = v$IN_5770_out0;
assign v$IN_2883_out0 = v$IN_5771_out0;
assign v$IN_3530_out0 = v$IN_12982_out0;
assign v$IN_3536_out0 = v$IN_12983_out0;
assign v$IN_3562_out0 = v$IN_12984_out0;
assign v$IN_3568_out0 = v$IN_12985_out0;
assign v$SEL3_4957_out0 = v$IN_9131_out0[47:32];
assign v$SEL3_4961_out0 = v$IN_9135_out0[47:32];
assign v$SEL3_4965_out0 = v$IN_9139_out0[47:32];
assign v$SEL3_4969_out0 = v$IN_9143_out0[47:32];
assign v$SEL2_9368_out0 = v$IN_9131_out0[31:16];
assign v$SEL2_9372_out0 = v$IN_9135_out0[31:16];
assign v$SEL2_9376_out0 = v$IN_9139_out0[31:16];
assign v$SEL2_9380_out0 = v$IN_9143_out0[31:16];
assign v$SEL1_11746_out0 = v$IN_9131_out0[15:0];
assign v$SEL1_11750_out0 = v$IN_9135_out0[15:0];
assign v$SEL1_11754_out0 = v$IN_9139_out0[15:0];
assign v$SEL1_11758_out0 = v$IN_9143_out0[15:0];
assign v$IN_2569_out0 = v$IN_3530_out0;
assign v$IN_2572_out0 = v$IN_3536_out0;
assign v$IN_2579_out0 = v$IN_3562_out0;
assign v$IN_2582_out0 = v$IN_3568_out0;
assign v$SEL15_3278_out0 = v$IN_2880_out0[33:33];
assign v$SEL15_3279_out0 = v$IN_2881_out0[33:33];
assign v$SEL15_3280_out0 = v$IN_2882_out0[33:33];
assign v$SEL15_3281_out0 = v$IN_2883_out0[33:33];
assign v$SEL13_4694_out0 = v$IN_2880_out0[35:35];
assign v$SEL13_4695_out0 = v$IN_2881_out0[35:35];
assign v$SEL13_4696_out0 = v$IN_2882_out0[35:35];
assign v$SEL13_4697_out0 = v$IN_2883_out0[35:35];
assign v$SEL1_4817_out0 = v$IN_2880_out0[47:47];
assign v$SEL1_4818_out0 = v$IN_2881_out0[47:47];
assign v$SEL1_4819_out0 = v$IN_2882_out0[47:47];
assign v$SEL1_4820_out0 = v$IN_2883_out0[47:47];
assign v$SEL11_4834_out0 = v$IN_2880_out0[37:37];
assign v$SEL11_4835_out0 = v$IN_2881_out0[37:37];
assign v$SEL11_4836_out0 = v$IN_2882_out0[37:37];
assign v$SEL11_4837_out0 = v$IN_2883_out0[37:37];
assign v$SEL4_4919_out0 = v$IN_2880_out0[44:44];
assign v$SEL4_4920_out0 = v$IN_2881_out0[44:44];
assign v$SEL4_4921_out0 = v$IN_2882_out0[44:44];
assign v$SEL4_4922_out0 = v$IN_2883_out0[44:44];
assign v$SEL22_4990_out0 = v$IN_2880_out0[26:26];
assign v$SEL22_4991_out0 = v$IN_2881_out0[26:26];
assign v$SEL22_4992_out0 = v$IN_2882_out0[26:26];
assign v$SEL22_4993_out0 = v$IN_2883_out0[26:26];
assign v$SEL23_5155_out0 = v$IN_2880_out0[25:25];
assign v$SEL23_5156_out0 = v$IN_2881_out0[25:25];
assign v$SEL23_5157_out0 = v$IN_2882_out0[25:25];
assign v$SEL23_5158_out0 = v$IN_2883_out0[25:25];
assign v$SEL20_5666_out0 = v$IN_2880_out0[28:28];
assign v$SEL20_5667_out0 = v$IN_2881_out0[28:28];
assign v$SEL20_5668_out0 = v$IN_2882_out0[28:28];
assign v$SEL20_5669_out0 = v$IN_2883_out0[28:28];
assign v$SEL10_6487_out0 = v$IN_2880_out0[40:40];
assign v$SEL10_6488_out0 = v$IN_2881_out0[40:40];
assign v$SEL10_6489_out0 = v$IN_2882_out0[40:40];
assign v$SEL10_6490_out0 = v$IN_2883_out0[40:40];
assign v$SEL9_6829_out0 = v$IN_2880_out0[38:38];
assign v$SEL9_6830_out0 = v$IN_2881_out0[38:38];
assign v$SEL9_6831_out0 = v$IN_2882_out0[38:38];
assign v$SEL9_6832_out0 = v$IN_2883_out0[38:38];
assign v$SEL21_7286_out0 = v$IN_2880_out0[27:27];
assign v$SEL21_7287_out0 = v$IN_2881_out0[27:27];
assign v$SEL21_7288_out0 = v$IN_2882_out0[27:27];
assign v$SEL21_7289_out0 = v$IN_2883_out0[27:27];
assign v$SEL18_7420_out0 = v$IN_2880_out0[30:30];
assign v$SEL18_7421_out0 = v$IN_2881_out0[30:30];
assign v$SEL18_7422_out0 = v$IN_2882_out0[30:30];
assign v$SEL18_7423_out0 = v$IN_2883_out0[30:30];
assign v$SEL3_7544_out0 = v$IN_2880_out0[45:45];
assign v$SEL3_7545_out0 = v$IN_2881_out0[45:45];
assign v$SEL3_7546_out0 = v$IN_2882_out0[45:45];
assign v$SEL3_7547_out0 = v$IN_2883_out0[45:45];
assign v$SEL6_8113_out0 = v$IN_2880_out0[42:42];
assign v$SEL6_8114_out0 = v$IN_2881_out0[42:42];
assign v$SEL6_8115_out0 = v$IN_2882_out0[42:42];
assign v$SEL6_8116_out0 = v$IN_2883_out0[42:42];
assign v$SEL19_8464_out0 = v$IN_2880_out0[29:29];
assign v$SEL19_8465_out0 = v$IN_2881_out0[29:29];
assign v$SEL19_8466_out0 = v$IN_2882_out0[29:29];
assign v$SEL19_8467_out0 = v$IN_2883_out0[29:29];
assign v$SEL2_8895_out0 = v$IN_2880_out0[46:46];
assign v$SEL2_8896_out0 = v$IN_2881_out0[46:46];
assign v$SEL2_8897_out0 = v$IN_2882_out0[46:46];
assign v$SEL2_8898_out0 = v$IN_2883_out0[46:46];
assign v$IN_9132_out0 = v$SEL1_11746_out0;
assign v$IN_9133_out0 = v$SEL2_9368_out0;
assign v$IN_9134_out0 = v$SEL3_4957_out0;
assign v$IN_9136_out0 = v$SEL1_11750_out0;
assign v$IN_9137_out0 = v$SEL2_9372_out0;
assign v$IN_9138_out0 = v$SEL3_4961_out0;
assign v$IN_9140_out0 = v$SEL1_11754_out0;
assign v$IN_9141_out0 = v$SEL2_9376_out0;
assign v$IN_9142_out0 = v$SEL3_4965_out0;
assign v$IN_9144_out0 = v$SEL1_11758_out0;
assign v$IN_9145_out0 = v$SEL2_9380_out0;
assign v$IN_9146_out0 = v$SEL3_4969_out0;
assign v$SEL12_9362_out0 = v$IN_2880_out0[36:36];
assign v$SEL12_9363_out0 = v$IN_2881_out0[36:36];
assign v$SEL12_9364_out0 = v$IN_2882_out0[36:36];
assign v$SEL12_9365_out0 = v$IN_2883_out0[36:36];
assign v$SEL7_9719_out0 = v$IN_2880_out0[41:41];
assign v$SEL7_9720_out0 = v$IN_2881_out0[41:41];
assign v$SEL7_9721_out0 = v$IN_2882_out0[41:41];
assign v$SEL7_9722_out0 = v$IN_2883_out0[41:41];
assign v$SEL5_10744_out0 = v$IN_2880_out0[43:43];
assign v$SEL5_10745_out0 = v$IN_2881_out0[43:43];
assign v$SEL5_10746_out0 = v$IN_2882_out0[43:43];
assign v$SEL5_10747_out0 = v$IN_2883_out0[43:43];
assign v$SEL17_11249_out0 = v$IN_2880_out0[31:31];
assign v$SEL17_11250_out0 = v$IN_2881_out0[31:31];
assign v$SEL17_11251_out0 = v$IN_2882_out0[31:31];
assign v$SEL17_11252_out0 = v$IN_2883_out0[31:31];
assign v$SEL14_11462_out0 = v$IN_2880_out0[34:34];
assign v$SEL14_11463_out0 = v$IN_2881_out0[34:34];
assign v$SEL14_11464_out0 = v$IN_2882_out0[34:34];
assign v$SEL14_11465_out0 = v$IN_2883_out0[34:34];
assign v$SEL16_11943_out0 = v$IN_2880_out0[32:32];
assign v$SEL16_11944_out0 = v$IN_2881_out0[32:32];
assign v$SEL16_11945_out0 = v$IN_2882_out0[32:32];
assign v$SEL16_11946_out0 = v$IN_2883_out0[32:32];
assign v$SEL24_11975_out0 = v$IN_2880_out0[24:24];
assign v$SEL24_11976_out0 = v$IN_2881_out0[24:24];
assign v$SEL24_11977_out0 = v$IN_2882_out0[24:24];
assign v$SEL24_11978_out0 = v$IN_2883_out0[24:24];
assign v$SEL8_12507_out0 = v$IN_2880_out0[39:39];
assign v$SEL8_12508_out0 = v$IN_2881_out0[39:39];
assign v$SEL8_12509_out0 = v$IN_2882_out0[39:39];
assign v$SEL8_12510_out0 = v$IN_2883_out0[39:39];
assign v$SEL4_2058_out0 = v$IN_9132_out0[15:12];
assign v$SEL4_2059_out0 = v$IN_9133_out0[15:12];
assign v$SEL4_2060_out0 = v$IN_9134_out0[15:12];
assign v$SEL4_2061_out0 = v$IN_9136_out0[15:12];
assign v$SEL4_2062_out0 = v$IN_9137_out0[15:12];
assign v$SEL4_2063_out0 = v$IN_9138_out0[15:12];
assign v$SEL4_2064_out0 = v$IN_9140_out0[15:12];
assign v$SEL4_2065_out0 = v$IN_9141_out0[15:12];
assign v$SEL4_2066_out0 = v$IN_9142_out0[15:12];
assign v$SEL4_2067_out0 = v$IN_9144_out0[15:12];
assign v$SEL4_2068_out0 = v$IN_9145_out0[15:12];
assign v$SEL4_2069_out0 = v$IN_9146_out0[15:12];
assign v$SEL3_4958_out0 = v$IN_9132_out0[11:8];
assign v$SEL3_4959_out0 = v$IN_9133_out0[11:8];
assign v$SEL3_4960_out0 = v$IN_9134_out0[11:8];
assign v$SEL3_4962_out0 = v$IN_9136_out0[11:8];
assign v$SEL3_4963_out0 = v$IN_9137_out0[11:8];
assign v$SEL3_4964_out0 = v$IN_9138_out0[11:8];
assign v$SEL3_4966_out0 = v$IN_9140_out0[11:8];
assign v$SEL3_4967_out0 = v$IN_9141_out0[11:8];
assign v$SEL3_4968_out0 = v$IN_9142_out0[11:8];
assign v$SEL3_4970_out0 = v$IN_9144_out0[11:8];
assign v$SEL3_4971_out0 = v$IN_9145_out0[11:8];
assign v$SEL3_4972_out0 = v$IN_9146_out0[11:8];
assign v$SEL1_5943_out0 = v$IN_2569_out0[47:1];
assign v$SEL1_5949_out0 = v$IN_2572_out0[47:1];
assign v$SEL1_5975_out0 = v$IN_2579_out0[47:1];
assign v$SEL1_5981_out0 = v$IN_2582_out0[47:1];
assign v$SEL2_9369_out0 = v$IN_9132_out0[7:4];
assign v$SEL2_9370_out0 = v$IN_9133_out0[7:4];
assign v$SEL2_9371_out0 = v$IN_9134_out0[7:4];
assign v$SEL2_9373_out0 = v$IN_9136_out0[7:4];
assign v$SEL2_9374_out0 = v$IN_9137_out0[7:4];
assign v$SEL2_9375_out0 = v$IN_9138_out0[7:4];
assign v$SEL2_9377_out0 = v$IN_9140_out0[7:4];
assign v$SEL2_9378_out0 = v$IN_9141_out0[7:4];
assign v$SEL2_9379_out0 = v$IN_9142_out0[7:4];
assign v$SEL2_9381_out0 = v$IN_9144_out0[7:4];
assign v$SEL2_9382_out0 = v$IN_9145_out0[7:4];
assign v$SEL2_9383_out0 = v$IN_9146_out0[7:4];
assign v$SEL1_10687_out0 = v$IN_2569_out0[46:0];
assign v$SEL1_10693_out0 = v$IN_2572_out0[46:0];
assign v$SEL1_10719_out0 = v$IN_2579_out0[46:0];
assign v$SEL1_10725_out0 = v$IN_2582_out0[46:0];
assign v$SEL1_11747_out0 = v$IN_9132_out0[3:0];
assign v$SEL1_11748_out0 = v$IN_9133_out0[3:0];
assign v$SEL1_11749_out0 = v$IN_9134_out0[3:0];
assign v$SEL1_11751_out0 = v$IN_9136_out0[3:0];
assign v$SEL1_11752_out0 = v$IN_9137_out0[3:0];
assign v$SEL1_11753_out0 = v$IN_9138_out0[3:0];
assign v$SEL1_11755_out0 = v$IN_9140_out0[3:0];
assign v$SEL1_11756_out0 = v$IN_9141_out0[3:0];
assign v$SEL1_11757_out0 = v$IN_9142_out0[3:0];
assign v$SEL1_11759_out0 = v$IN_9144_out0[3:0];
assign v$SEL1_11760_out0 = v$IN_9145_out0[3:0];
assign v$SEL1_11761_out0 = v$IN_9146_out0[3:0];
assign v$MUX24_12821_out0 = v$EQ24_1445_out0 ? v$SEL24_11975_out0 : v$C1_10973_out0;
assign v$MUX24_12822_out0 = v$EQ24_1446_out0 ? v$SEL24_11976_out0 : v$C1_10974_out0;
assign v$MUX24_12823_out0 = v$EQ24_1447_out0 ? v$SEL24_11977_out0 : v$C1_10975_out0;
assign v$MUX24_12824_out0 = v$EQ24_1448_out0 ? v$SEL24_11978_out0 : v$C1_10976_out0;
assign v$_2929_out0 = { v$C2_105_out0,v$SEL1_10687_out0 };
assign v$_2935_out0 = { v$C2_111_out0,v$SEL1_10693_out0 };
assign v$_2961_out0 = { v$C2_137_out0,v$SEL1_10719_out0 };
assign v$_2967_out0 = { v$C2_143_out0,v$SEL1_10725_out0 };
assign v$_6236_out0 = { v$SEL1_5943_out0,v$C1_3972_out0 };
assign v$_6242_out0 = { v$SEL1_5949_out0,v$C1_3978_out0 };
assign v$_6268_out0 = { v$SEL1_5975_out0,v$C1_4004_out0 };
assign v$_6274_out0 = { v$SEL1_5981_out0,v$C1_4010_out0 };
assign v$IN_10358_out0 = v$SEL3_4958_out0;
assign v$IN_10359_out0 = v$SEL1_11747_out0;
assign v$IN_10360_out0 = v$SEL2_9369_out0;
assign v$IN_10361_out0 = v$SEL4_2058_out0;
assign v$IN_10362_out0 = v$SEL3_4959_out0;
assign v$IN_10363_out0 = v$SEL1_11748_out0;
assign v$IN_10364_out0 = v$SEL2_9370_out0;
assign v$IN_10365_out0 = v$SEL4_2059_out0;
assign v$IN_10366_out0 = v$SEL3_4960_out0;
assign v$IN_10367_out0 = v$SEL1_11749_out0;
assign v$IN_10368_out0 = v$SEL2_9371_out0;
assign v$IN_10369_out0 = v$SEL4_2060_out0;
assign v$IN_10370_out0 = v$SEL3_4962_out0;
assign v$IN_10371_out0 = v$SEL1_11751_out0;
assign v$IN_10372_out0 = v$SEL2_9373_out0;
assign v$IN_10373_out0 = v$SEL4_2061_out0;
assign v$IN_10374_out0 = v$SEL3_4963_out0;
assign v$IN_10375_out0 = v$SEL1_11752_out0;
assign v$IN_10376_out0 = v$SEL2_9374_out0;
assign v$IN_10377_out0 = v$SEL4_2062_out0;
assign v$IN_10378_out0 = v$SEL3_4964_out0;
assign v$IN_10379_out0 = v$SEL1_11753_out0;
assign v$IN_10380_out0 = v$SEL2_9375_out0;
assign v$IN_10381_out0 = v$SEL4_2063_out0;
assign v$IN_10388_out0 = v$SEL3_4966_out0;
assign v$IN_10389_out0 = v$SEL1_11755_out0;
assign v$IN_10390_out0 = v$SEL2_9377_out0;
assign v$IN_10391_out0 = v$SEL4_2064_out0;
assign v$IN_10392_out0 = v$SEL3_4967_out0;
assign v$IN_10393_out0 = v$SEL1_11756_out0;
assign v$IN_10394_out0 = v$SEL2_9378_out0;
assign v$IN_10395_out0 = v$SEL4_2065_out0;
assign v$IN_10396_out0 = v$SEL3_4968_out0;
assign v$IN_10397_out0 = v$SEL1_11757_out0;
assign v$IN_10398_out0 = v$SEL2_9379_out0;
assign v$IN_10399_out0 = v$SEL4_2066_out0;
assign v$IN_10400_out0 = v$SEL3_4970_out0;
assign v$IN_10401_out0 = v$SEL1_11759_out0;
assign v$IN_10402_out0 = v$SEL2_9381_out0;
assign v$IN_10403_out0 = v$SEL4_2067_out0;
assign v$IN_10404_out0 = v$SEL3_4971_out0;
assign v$IN_10405_out0 = v$SEL1_11760_out0;
assign v$IN_10406_out0 = v$SEL2_9382_out0;
assign v$IN_10407_out0 = v$SEL4_2068_out0;
assign v$IN_10408_out0 = v$SEL3_4972_out0;
assign v$IN_10409_out0 = v$SEL1_11761_out0;
assign v$IN_10410_out0 = v$SEL2_9383_out0;
assign v$IN_10411_out0 = v$SEL4_2069_out0;
assign v$MUX23_11379_out0 = v$EQ23_1913_out0 ? v$SEL23_5155_out0 : v$MUX24_12821_out0;
assign v$MUX23_11380_out0 = v$EQ23_1914_out0 ? v$SEL23_5156_out0 : v$MUX24_12822_out0;
assign v$MUX23_11381_out0 = v$EQ23_1915_out0 ? v$SEL23_5157_out0 : v$MUX24_12823_out0;
assign v$MUX23_11382_out0 = v$EQ23_1916_out0 ? v$SEL23_5158_out0 : v$MUX24_12824_out0;
assign v$SEL3_1217_out0 = v$IN_10358_out0[2:2];
assign v$SEL3_1218_out0 = v$IN_10359_out0[2:2];
assign v$SEL3_1219_out0 = v$IN_10360_out0[2:2];
assign v$SEL3_1220_out0 = v$IN_10361_out0[2:2];
assign v$SEL3_1221_out0 = v$IN_10362_out0[2:2];
assign v$SEL3_1222_out0 = v$IN_10363_out0[2:2];
assign v$SEL3_1223_out0 = v$IN_10364_out0[2:2];
assign v$SEL3_1224_out0 = v$IN_10365_out0[2:2];
assign v$SEL3_1225_out0 = v$IN_10366_out0[2:2];
assign v$SEL3_1226_out0 = v$IN_10367_out0[2:2];
assign v$SEL3_1227_out0 = v$IN_10368_out0[2:2];
assign v$SEL3_1228_out0 = v$IN_10369_out0[2:2];
assign v$SEL3_1229_out0 = v$IN_10370_out0[2:2];
assign v$SEL3_1230_out0 = v$IN_10371_out0[2:2];
assign v$SEL3_1231_out0 = v$IN_10372_out0[2:2];
assign v$SEL3_1232_out0 = v$IN_10373_out0[2:2];
assign v$SEL3_1233_out0 = v$IN_10374_out0[2:2];
assign v$SEL3_1234_out0 = v$IN_10375_out0[2:2];
assign v$SEL3_1235_out0 = v$IN_10376_out0[2:2];
assign v$SEL3_1236_out0 = v$IN_10377_out0[2:2];
assign v$SEL3_1237_out0 = v$IN_10378_out0[2:2];
assign v$SEL3_1238_out0 = v$IN_10379_out0[2:2];
assign v$SEL3_1239_out0 = v$IN_10380_out0[2:2];
assign v$SEL3_1240_out0 = v$IN_10381_out0[2:2];
assign v$SEL3_1247_out0 = v$IN_10388_out0[2:2];
assign v$SEL3_1248_out0 = v$IN_10389_out0[2:2];
assign v$SEL3_1249_out0 = v$IN_10390_out0[2:2];
assign v$SEL3_1250_out0 = v$IN_10391_out0[2:2];
assign v$SEL3_1251_out0 = v$IN_10392_out0[2:2];
assign v$SEL3_1252_out0 = v$IN_10393_out0[2:2];
assign v$SEL3_1253_out0 = v$IN_10394_out0[2:2];
assign v$SEL3_1254_out0 = v$IN_10395_out0[2:2];
assign v$SEL3_1255_out0 = v$IN_10396_out0[2:2];
assign v$SEL3_1256_out0 = v$IN_10397_out0[2:2];
assign v$SEL3_1257_out0 = v$IN_10398_out0[2:2];
assign v$SEL3_1258_out0 = v$IN_10399_out0[2:2];
assign v$SEL3_1259_out0 = v$IN_10400_out0[2:2];
assign v$SEL3_1260_out0 = v$IN_10401_out0[2:2];
assign v$SEL3_1261_out0 = v$IN_10402_out0[2:2];
assign v$SEL3_1262_out0 = v$IN_10403_out0[2:2];
assign v$SEL3_1263_out0 = v$IN_10404_out0[2:2];
assign v$SEL3_1264_out0 = v$IN_10405_out0[2:2];
assign v$SEL3_1265_out0 = v$IN_10406_out0[2:2];
assign v$SEL3_1266_out0 = v$IN_10407_out0[2:2];
assign v$SEL3_1267_out0 = v$IN_10408_out0[2:2];
assign v$SEL3_1268_out0 = v$IN_10409_out0[2:2];
assign v$SEL3_1269_out0 = v$IN_10410_out0[2:2];
assign v$SEL3_1270_out0 = v$IN_10411_out0[2:2];
assign v$MUX1_1292_out0 = v$LEFT$SHIT_1804_out0 ? v$_2929_out0 : v$_6236_out0;
assign v$MUX1_1298_out0 = v$LEFT$SHIT_1810_out0 ? v$_2935_out0 : v$_6242_out0;
assign v$MUX1_1324_out0 = v$LEFT$SHIT_1836_out0 ? v$_2961_out0 : v$_6268_out0;
assign v$MUX1_1330_out0 = v$LEFT$SHIT_1842_out0 ? v$_2967_out0 : v$_6274_out0;
assign v$SEL4_4081_out0 = v$IN_10358_out0[3:3];
assign v$SEL4_4082_out0 = v$IN_10359_out0[3:3];
assign v$SEL4_4083_out0 = v$IN_10360_out0[3:3];
assign v$SEL4_4084_out0 = v$IN_10361_out0[3:3];
assign v$SEL4_4085_out0 = v$IN_10362_out0[3:3];
assign v$SEL4_4086_out0 = v$IN_10363_out0[3:3];
assign v$SEL4_4087_out0 = v$IN_10364_out0[3:3];
assign v$SEL4_4088_out0 = v$IN_10365_out0[3:3];
assign v$SEL4_4089_out0 = v$IN_10366_out0[3:3];
assign v$SEL4_4090_out0 = v$IN_10367_out0[3:3];
assign v$SEL4_4091_out0 = v$IN_10368_out0[3:3];
assign v$SEL4_4092_out0 = v$IN_10369_out0[3:3];
assign v$SEL4_4093_out0 = v$IN_10370_out0[3:3];
assign v$SEL4_4094_out0 = v$IN_10371_out0[3:3];
assign v$SEL4_4095_out0 = v$IN_10372_out0[3:3];
assign v$SEL4_4096_out0 = v$IN_10373_out0[3:3];
assign v$SEL4_4097_out0 = v$IN_10374_out0[3:3];
assign v$SEL4_4098_out0 = v$IN_10375_out0[3:3];
assign v$SEL4_4099_out0 = v$IN_10376_out0[3:3];
assign v$SEL4_4100_out0 = v$IN_10377_out0[3:3];
assign v$SEL4_4101_out0 = v$IN_10378_out0[3:3];
assign v$SEL4_4102_out0 = v$IN_10379_out0[3:3];
assign v$SEL4_4103_out0 = v$IN_10380_out0[3:3];
assign v$SEL4_4104_out0 = v$IN_10381_out0[3:3];
assign v$SEL4_4111_out0 = v$IN_10388_out0[3:3];
assign v$SEL4_4112_out0 = v$IN_10389_out0[3:3];
assign v$SEL4_4113_out0 = v$IN_10390_out0[3:3];
assign v$SEL4_4114_out0 = v$IN_10391_out0[3:3];
assign v$SEL4_4115_out0 = v$IN_10392_out0[3:3];
assign v$SEL4_4116_out0 = v$IN_10393_out0[3:3];
assign v$SEL4_4117_out0 = v$IN_10394_out0[3:3];
assign v$SEL4_4118_out0 = v$IN_10395_out0[3:3];
assign v$SEL4_4119_out0 = v$IN_10396_out0[3:3];
assign v$SEL4_4120_out0 = v$IN_10397_out0[3:3];
assign v$SEL4_4121_out0 = v$IN_10398_out0[3:3];
assign v$SEL4_4122_out0 = v$IN_10399_out0[3:3];
assign v$SEL4_4123_out0 = v$IN_10400_out0[3:3];
assign v$SEL4_4124_out0 = v$IN_10401_out0[3:3];
assign v$SEL4_4125_out0 = v$IN_10402_out0[3:3];
assign v$SEL4_4126_out0 = v$IN_10403_out0[3:3];
assign v$SEL4_4127_out0 = v$IN_10404_out0[3:3];
assign v$SEL4_4128_out0 = v$IN_10405_out0[3:3];
assign v$SEL4_4129_out0 = v$IN_10406_out0[3:3];
assign v$SEL4_4130_out0 = v$IN_10407_out0[3:3];
assign v$SEL4_4131_out0 = v$IN_10408_out0[3:3];
assign v$SEL4_4132_out0 = v$IN_10409_out0[3:3];
assign v$SEL4_4133_out0 = v$IN_10410_out0[3:3];
assign v$SEL4_4134_out0 = v$IN_10411_out0[3:3];
assign v$SEL2_5201_out0 = v$IN_10358_out0[1:1];
assign v$SEL2_5202_out0 = v$IN_10359_out0[1:1];
assign v$SEL2_5203_out0 = v$IN_10360_out0[1:1];
assign v$SEL2_5204_out0 = v$IN_10361_out0[1:1];
assign v$SEL2_5205_out0 = v$IN_10362_out0[1:1];
assign v$SEL2_5206_out0 = v$IN_10363_out0[1:1];
assign v$SEL2_5207_out0 = v$IN_10364_out0[1:1];
assign v$SEL2_5208_out0 = v$IN_10365_out0[1:1];
assign v$SEL2_5209_out0 = v$IN_10366_out0[1:1];
assign v$SEL2_5210_out0 = v$IN_10367_out0[1:1];
assign v$SEL2_5211_out0 = v$IN_10368_out0[1:1];
assign v$SEL2_5212_out0 = v$IN_10369_out0[1:1];
assign v$SEL2_5213_out0 = v$IN_10370_out0[1:1];
assign v$SEL2_5214_out0 = v$IN_10371_out0[1:1];
assign v$SEL2_5215_out0 = v$IN_10372_out0[1:1];
assign v$SEL2_5216_out0 = v$IN_10373_out0[1:1];
assign v$SEL2_5217_out0 = v$IN_10374_out0[1:1];
assign v$SEL2_5218_out0 = v$IN_10375_out0[1:1];
assign v$SEL2_5219_out0 = v$IN_10376_out0[1:1];
assign v$SEL2_5220_out0 = v$IN_10377_out0[1:1];
assign v$SEL2_5221_out0 = v$IN_10378_out0[1:1];
assign v$SEL2_5222_out0 = v$IN_10379_out0[1:1];
assign v$SEL2_5223_out0 = v$IN_10380_out0[1:1];
assign v$SEL2_5224_out0 = v$IN_10381_out0[1:1];
assign v$SEL2_5231_out0 = v$IN_10388_out0[1:1];
assign v$SEL2_5232_out0 = v$IN_10389_out0[1:1];
assign v$SEL2_5233_out0 = v$IN_10390_out0[1:1];
assign v$SEL2_5234_out0 = v$IN_10391_out0[1:1];
assign v$SEL2_5235_out0 = v$IN_10392_out0[1:1];
assign v$SEL2_5236_out0 = v$IN_10393_out0[1:1];
assign v$SEL2_5237_out0 = v$IN_10394_out0[1:1];
assign v$SEL2_5238_out0 = v$IN_10395_out0[1:1];
assign v$SEL2_5239_out0 = v$IN_10396_out0[1:1];
assign v$SEL2_5240_out0 = v$IN_10397_out0[1:1];
assign v$SEL2_5241_out0 = v$IN_10398_out0[1:1];
assign v$SEL2_5242_out0 = v$IN_10399_out0[1:1];
assign v$SEL2_5243_out0 = v$IN_10400_out0[1:1];
assign v$SEL2_5244_out0 = v$IN_10401_out0[1:1];
assign v$SEL2_5245_out0 = v$IN_10402_out0[1:1];
assign v$SEL2_5246_out0 = v$IN_10403_out0[1:1];
assign v$SEL2_5247_out0 = v$IN_10404_out0[1:1];
assign v$SEL2_5248_out0 = v$IN_10405_out0[1:1];
assign v$SEL2_5249_out0 = v$IN_10406_out0[1:1];
assign v$SEL2_5250_out0 = v$IN_10407_out0[1:1];
assign v$SEL2_5251_out0 = v$IN_10408_out0[1:1];
assign v$SEL2_5252_out0 = v$IN_10409_out0[1:1];
assign v$SEL2_5253_out0 = v$IN_10410_out0[1:1];
assign v$SEL2_5254_out0 = v$IN_10411_out0[1:1];
assign v$SEL1_9025_out0 = v$IN_10358_out0[0:0];
assign v$SEL1_9026_out0 = v$IN_10359_out0[0:0];
assign v$SEL1_9027_out0 = v$IN_10360_out0[0:0];
assign v$SEL1_9028_out0 = v$IN_10361_out0[0:0];
assign v$SEL1_9029_out0 = v$IN_10362_out0[0:0];
assign v$SEL1_9030_out0 = v$IN_10363_out0[0:0];
assign v$SEL1_9031_out0 = v$IN_10364_out0[0:0];
assign v$SEL1_9032_out0 = v$IN_10365_out0[0:0];
assign v$SEL1_9033_out0 = v$IN_10366_out0[0:0];
assign v$SEL1_9034_out0 = v$IN_10367_out0[0:0];
assign v$SEL1_9035_out0 = v$IN_10368_out0[0:0];
assign v$SEL1_9036_out0 = v$IN_10369_out0[0:0];
assign v$SEL1_9037_out0 = v$IN_10370_out0[0:0];
assign v$SEL1_9038_out0 = v$IN_10371_out0[0:0];
assign v$SEL1_9039_out0 = v$IN_10372_out0[0:0];
assign v$SEL1_9040_out0 = v$IN_10373_out0[0:0];
assign v$SEL1_9041_out0 = v$IN_10374_out0[0:0];
assign v$SEL1_9042_out0 = v$IN_10375_out0[0:0];
assign v$SEL1_9043_out0 = v$IN_10376_out0[0:0];
assign v$SEL1_9044_out0 = v$IN_10377_out0[0:0];
assign v$SEL1_9045_out0 = v$IN_10378_out0[0:0];
assign v$SEL1_9046_out0 = v$IN_10379_out0[0:0];
assign v$SEL1_9047_out0 = v$IN_10380_out0[0:0];
assign v$SEL1_9048_out0 = v$IN_10381_out0[0:0];
assign v$SEL1_9055_out0 = v$IN_10388_out0[0:0];
assign v$SEL1_9056_out0 = v$IN_10389_out0[0:0];
assign v$SEL1_9057_out0 = v$IN_10390_out0[0:0];
assign v$SEL1_9058_out0 = v$IN_10391_out0[0:0];
assign v$SEL1_9059_out0 = v$IN_10392_out0[0:0];
assign v$SEL1_9060_out0 = v$IN_10393_out0[0:0];
assign v$SEL1_9061_out0 = v$IN_10394_out0[0:0];
assign v$SEL1_9062_out0 = v$IN_10395_out0[0:0];
assign v$SEL1_9063_out0 = v$IN_10396_out0[0:0];
assign v$SEL1_9064_out0 = v$IN_10397_out0[0:0];
assign v$SEL1_9065_out0 = v$IN_10398_out0[0:0];
assign v$SEL1_9066_out0 = v$IN_10399_out0[0:0];
assign v$SEL1_9067_out0 = v$IN_10400_out0[0:0];
assign v$SEL1_9068_out0 = v$IN_10401_out0[0:0];
assign v$SEL1_9069_out0 = v$IN_10402_out0[0:0];
assign v$SEL1_9070_out0 = v$IN_10403_out0[0:0];
assign v$SEL1_9071_out0 = v$IN_10404_out0[0:0];
assign v$SEL1_9072_out0 = v$IN_10405_out0[0:0];
assign v$SEL1_9073_out0 = v$IN_10406_out0[0:0];
assign v$SEL1_9074_out0 = v$IN_10407_out0[0:0];
assign v$SEL1_9075_out0 = v$IN_10408_out0[0:0];
assign v$SEL1_9076_out0 = v$IN_10409_out0[0:0];
assign v$SEL1_9077_out0 = v$IN_10410_out0[0:0];
assign v$SEL1_9078_out0 = v$IN_10411_out0[0:0];
assign v$MUX22_11542_out0 = v$EQ22_1599_out0 ? v$SEL22_4990_out0 : v$MUX23_11379_out0;
assign v$MUX22_11543_out0 = v$EQ22_1600_out0 ? v$SEL22_4991_out0 : v$MUX23_11380_out0;
assign v$MUX22_11544_out0 = v$EQ22_1601_out0 ? v$SEL22_4992_out0 : v$MUX23_11381_out0;
assign v$MUX22_11545_out0 = v$EQ22_1602_out0 ? v$SEL22_4993_out0 : v$MUX23_11382_out0;
assign v$G10_605_out0 = !(v$SEL1_9025_out0 || v$SEL2_5201_out0);
assign v$G10_606_out0 = !(v$SEL1_9026_out0 || v$SEL2_5202_out0);
assign v$G10_607_out0 = !(v$SEL1_9027_out0 || v$SEL2_5203_out0);
assign v$G10_608_out0 = !(v$SEL1_9028_out0 || v$SEL2_5204_out0);
assign v$G10_609_out0 = !(v$SEL1_9029_out0 || v$SEL2_5205_out0);
assign v$G10_610_out0 = !(v$SEL1_9030_out0 || v$SEL2_5206_out0);
assign v$G10_611_out0 = !(v$SEL1_9031_out0 || v$SEL2_5207_out0);
assign v$G10_612_out0 = !(v$SEL1_9032_out0 || v$SEL2_5208_out0);
assign v$G10_613_out0 = !(v$SEL1_9033_out0 || v$SEL2_5209_out0);
assign v$G10_614_out0 = !(v$SEL1_9034_out0 || v$SEL2_5210_out0);
assign v$G10_615_out0 = !(v$SEL1_9035_out0 || v$SEL2_5211_out0);
assign v$G10_616_out0 = !(v$SEL1_9036_out0 || v$SEL2_5212_out0);
assign v$G10_617_out0 = !(v$SEL1_9037_out0 || v$SEL2_5213_out0);
assign v$G10_618_out0 = !(v$SEL1_9038_out0 || v$SEL2_5214_out0);
assign v$G10_619_out0 = !(v$SEL1_9039_out0 || v$SEL2_5215_out0);
assign v$G10_620_out0 = !(v$SEL1_9040_out0 || v$SEL2_5216_out0);
assign v$G10_621_out0 = !(v$SEL1_9041_out0 || v$SEL2_5217_out0);
assign v$G10_622_out0 = !(v$SEL1_9042_out0 || v$SEL2_5218_out0);
assign v$G10_623_out0 = !(v$SEL1_9043_out0 || v$SEL2_5219_out0);
assign v$G10_624_out0 = !(v$SEL1_9044_out0 || v$SEL2_5220_out0);
assign v$G10_625_out0 = !(v$SEL1_9045_out0 || v$SEL2_5221_out0);
assign v$G10_626_out0 = !(v$SEL1_9046_out0 || v$SEL2_5222_out0);
assign v$G10_627_out0 = !(v$SEL1_9047_out0 || v$SEL2_5223_out0);
assign v$G10_628_out0 = !(v$SEL1_9048_out0 || v$SEL2_5224_out0);
assign v$G10_635_out0 = !(v$SEL1_9055_out0 || v$SEL2_5231_out0);
assign v$G10_636_out0 = !(v$SEL1_9056_out0 || v$SEL2_5232_out0);
assign v$G10_637_out0 = !(v$SEL1_9057_out0 || v$SEL2_5233_out0);
assign v$G10_638_out0 = !(v$SEL1_9058_out0 || v$SEL2_5234_out0);
assign v$G10_639_out0 = !(v$SEL1_9059_out0 || v$SEL2_5235_out0);
assign v$G10_640_out0 = !(v$SEL1_9060_out0 || v$SEL2_5236_out0);
assign v$G10_641_out0 = !(v$SEL1_9061_out0 || v$SEL2_5237_out0);
assign v$G10_642_out0 = !(v$SEL1_9062_out0 || v$SEL2_5238_out0);
assign v$G10_643_out0 = !(v$SEL1_9063_out0 || v$SEL2_5239_out0);
assign v$G10_644_out0 = !(v$SEL1_9064_out0 || v$SEL2_5240_out0);
assign v$G10_645_out0 = !(v$SEL1_9065_out0 || v$SEL2_5241_out0);
assign v$G10_646_out0 = !(v$SEL1_9066_out0 || v$SEL2_5242_out0);
assign v$G10_647_out0 = !(v$SEL1_9067_out0 || v$SEL2_5243_out0);
assign v$G10_648_out0 = !(v$SEL1_9068_out0 || v$SEL2_5244_out0);
assign v$G10_649_out0 = !(v$SEL1_9069_out0 || v$SEL2_5245_out0);
assign v$G10_650_out0 = !(v$SEL1_9070_out0 || v$SEL2_5246_out0);
assign v$G10_651_out0 = !(v$SEL1_9071_out0 || v$SEL2_5247_out0);
assign v$G10_652_out0 = !(v$SEL1_9072_out0 || v$SEL2_5248_out0);
assign v$G10_653_out0 = !(v$SEL1_9073_out0 || v$SEL2_5249_out0);
assign v$G10_654_out0 = !(v$SEL1_9074_out0 || v$SEL2_5250_out0);
assign v$G10_655_out0 = !(v$SEL1_9075_out0 || v$SEL2_5251_out0);
assign v$G10_656_out0 = !(v$SEL1_9076_out0 || v$SEL2_5252_out0);
assign v$G10_657_out0 = !(v$SEL1_9077_out0 || v$SEL2_5253_out0);
assign v$G10_658_out0 = !(v$SEL1_9078_out0 || v$SEL2_5254_out0);
assign v$G6_2256_out0 = ! v$SEL2_5201_out0;
assign v$G6_2257_out0 = ! v$SEL2_5202_out0;
assign v$G6_2258_out0 = ! v$SEL2_5203_out0;
assign v$G6_2259_out0 = ! v$SEL2_5204_out0;
assign v$G6_2260_out0 = ! v$SEL2_5205_out0;
assign v$G6_2261_out0 = ! v$SEL2_5206_out0;
assign v$G6_2262_out0 = ! v$SEL2_5207_out0;
assign v$G6_2263_out0 = ! v$SEL2_5208_out0;
assign v$G6_2264_out0 = ! v$SEL2_5209_out0;
assign v$G6_2265_out0 = ! v$SEL2_5210_out0;
assign v$G6_2266_out0 = ! v$SEL2_5211_out0;
assign v$G6_2267_out0 = ! v$SEL2_5212_out0;
assign v$G6_2268_out0 = ! v$SEL2_5213_out0;
assign v$G6_2269_out0 = ! v$SEL2_5214_out0;
assign v$G6_2270_out0 = ! v$SEL2_5215_out0;
assign v$G6_2271_out0 = ! v$SEL2_5216_out0;
assign v$G6_2272_out0 = ! v$SEL2_5217_out0;
assign v$G6_2273_out0 = ! v$SEL2_5218_out0;
assign v$G6_2274_out0 = ! v$SEL2_5219_out0;
assign v$G6_2275_out0 = ! v$SEL2_5220_out0;
assign v$G6_2276_out0 = ! v$SEL2_5221_out0;
assign v$G6_2277_out0 = ! v$SEL2_5222_out0;
assign v$G6_2278_out0 = ! v$SEL2_5223_out0;
assign v$G6_2279_out0 = ! v$SEL2_5224_out0;
assign v$G6_2286_out0 = ! v$SEL2_5231_out0;
assign v$G6_2287_out0 = ! v$SEL2_5232_out0;
assign v$G6_2288_out0 = ! v$SEL2_5233_out0;
assign v$G6_2289_out0 = ! v$SEL2_5234_out0;
assign v$G6_2290_out0 = ! v$SEL2_5235_out0;
assign v$G6_2291_out0 = ! v$SEL2_5236_out0;
assign v$G6_2292_out0 = ! v$SEL2_5237_out0;
assign v$G6_2293_out0 = ! v$SEL2_5238_out0;
assign v$G6_2294_out0 = ! v$SEL2_5239_out0;
assign v$G6_2295_out0 = ! v$SEL2_5240_out0;
assign v$G6_2296_out0 = ! v$SEL2_5241_out0;
assign v$G6_2297_out0 = ! v$SEL2_5242_out0;
assign v$G6_2298_out0 = ! v$SEL2_5243_out0;
assign v$G6_2299_out0 = ! v$SEL2_5244_out0;
assign v$G6_2300_out0 = ! v$SEL2_5245_out0;
assign v$G6_2301_out0 = ! v$SEL2_5246_out0;
assign v$G6_2302_out0 = ! v$SEL2_5247_out0;
assign v$G6_2303_out0 = ! v$SEL2_5248_out0;
assign v$G6_2304_out0 = ! v$SEL2_5249_out0;
assign v$G6_2305_out0 = ! v$SEL2_5250_out0;
assign v$G6_2306_out0 = ! v$SEL2_5251_out0;
assign v$G6_2307_out0 = ! v$SEL2_5252_out0;
assign v$G6_2308_out0 = ! v$SEL2_5253_out0;
assign v$G6_2309_out0 = ! v$SEL2_5254_out0;
assign v$MUX21_3294_out0 = v$EQ21_2017_out0 ? v$SEL21_7286_out0 : v$MUX22_11542_out0;
assign v$MUX21_3295_out0 = v$EQ21_2018_out0 ? v$SEL21_7287_out0 : v$MUX22_11543_out0;
assign v$MUX21_3296_out0 = v$EQ21_2019_out0 ? v$SEL21_7288_out0 : v$MUX22_11544_out0;
assign v$MUX21_3297_out0 = v$EQ21_2020_out0 ? v$SEL21_7289_out0 : v$MUX22_11545_out0;
assign v$G5_3846_out0 = ! v$SEL4_4081_out0;
assign v$G5_3847_out0 = ! v$SEL4_4082_out0;
assign v$G5_3848_out0 = ! v$SEL4_4083_out0;
assign v$G5_3849_out0 = ! v$SEL4_4084_out0;
assign v$G5_3850_out0 = ! v$SEL4_4085_out0;
assign v$G5_3851_out0 = ! v$SEL4_4086_out0;
assign v$G5_3852_out0 = ! v$SEL4_4087_out0;
assign v$G5_3853_out0 = ! v$SEL4_4088_out0;
assign v$G5_3854_out0 = ! v$SEL4_4089_out0;
assign v$G5_3855_out0 = ! v$SEL4_4090_out0;
assign v$G5_3856_out0 = ! v$SEL4_4091_out0;
assign v$G5_3857_out0 = ! v$SEL4_4092_out0;
assign v$G5_3858_out0 = ! v$SEL4_4093_out0;
assign v$G5_3859_out0 = ! v$SEL4_4094_out0;
assign v$G5_3860_out0 = ! v$SEL4_4095_out0;
assign v$G5_3861_out0 = ! v$SEL4_4096_out0;
assign v$G5_3862_out0 = ! v$SEL4_4097_out0;
assign v$G5_3863_out0 = ! v$SEL4_4098_out0;
assign v$G5_3864_out0 = ! v$SEL4_4099_out0;
assign v$G5_3865_out0 = ! v$SEL4_4100_out0;
assign v$G5_3866_out0 = ! v$SEL4_4101_out0;
assign v$G5_3867_out0 = ! v$SEL4_4102_out0;
assign v$G5_3868_out0 = ! v$SEL4_4103_out0;
assign v$G5_3869_out0 = ! v$SEL4_4104_out0;
assign v$G5_3876_out0 = ! v$SEL4_4111_out0;
assign v$G5_3877_out0 = ! v$SEL4_4112_out0;
assign v$G5_3878_out0 = ! v$SEL4_4113_out0;
assign v$G5_3879_out0 = ! v$SEL4_4114_out0;
assign v$G5_3880_out0 = ! v$SEL4_4115_out0;
assign v$G5_3881_out0 = ! v$SEL4_4116_out0;
assign v$G5_3882_out0 = ! v$SEL4_4117_out0;
assign v$G5_3883_out0 = ! v$SEL4_4118_out0;
assign v$G5_3884_out0 = ! v$SEL4_4119_out0;
assign v$G5_3885_out0 = ! v$SEL4_4120_out0;
assign v$G5_3886_out0 = ! v$SEL4_4121_out0;
assign v$G5_3887_out0 = ! v$SEL4_4122_out0;
assign v$G5_3888_out0 = ! v$SEL4_4123_out0;
assign v$G5_3889_out0 = ! v$SEL4_4124_out0;
assign v$G5_3890_out0 = ! v$SEL4_4125_out0;
assign v$G5_3891_out0 = ! v$SEL4_4126_out0;
assign v$G5_3892_out0 = ! v$SEL4_4127_out0;
assign v$G5_3893_out0 = ! v$SEL4_4128_out0;
assign v$G5_3894_out0 = ! v$SEL4_4129_out0;
assign v$G5_3895_out0 = ! v$SEL4_4130_out0;
assign v$G5_3896_out0 = ! v$SEL4_4131_out0;
assign v$G5_3897_out0 = ! v$SEL4_4132_out0;
assign v$G5_3898_out0 = ! v$SEL4_4133_out0;
assign v$G5_3899_out0 = ! v$SEL4_4134_out0;
assign v$G11_6081_out0 = !(v$SEL3_1217_out0 || v$SEL4_4081_out0);
assign v$G11_6082_out0 = !(v$SEL3_1218_out0 || v$SEL4_4082_out0);
assign v$G11_6083_out0 = !(v$SEL3_1219_out0 || v$SEL4_4083_out0);
assign v$G11_6084_out0 = !(v$SEL3_1220_out0 || v$SEL4_4084_out0);
assign v$G11_6085_out0 = !(v$SEL3_1221_out0 || v$SEL4_4085_out0);
assign v$G11_6086_out0 = !(v$SEL3_1222_out0 || v$SEL4_4086_out0);
assign v$G11_6087_out0 = !(v$SEL3_1223_out0 || v$SEL4_4087_out0);
assign v$G11_6088_out0 = !(v$SEL3_1224_out0 || v$SEL4_4088_out0);
assign v$G11_6089_out0 = !(v$SEL3_1225_out0 || v$SEL4_4089_out0);
assign v$G11_6090_out0 = !(v$SEL3_1226_out0 || v$SEL4_4090_out0);
assign v$G11_6091_out0 = !(v$SEL3_1227_out0 || v$SEL4_4091_out0);
assign v$G11_6092_out0 = !(v$SEL3_1228_out0 || v$SEL4_4092_out0);
assign v$G11_6093_out0 = !(v$SEL3_1229_out0 || v$SEL4_4093_out0);
assign v$G11_6094_out0 = !(v$SEL3_1230_out0 || v$SEL4_4094_out0);
assign v$G11_6095_out0 = !(v$SEL3_1231_out0 || v$SEL4_4095_out0);
assign v$G11_6096_out0 = !(v$SEL3_1232_out0 || v$SEL4_4096_out0);
assign v$G11_6097_out0 = !(v$SEL3_1233_out0 || v$SEL4_4097_out0);
assign v$G11_6098_out0 = !(v$SEL3_1234_out0 || v$SEL4_4098_out0);
assign v$G11_6099_out0 = !(v$SEL3_1235_out0 || v$SEL4_4099_out0);
assign v$G11_6100_out0 = !(v$SEL3_1236_out0 || v$SEL4_4100_out0);
assign v$G11_6101_out0 = !(v$SEL3_1237_out0 || v$SEL4_4101_out0);
assign v$G11_6102_out0 = !(v$SEL3_1238_out0 || v$SEL4_4102_out0);
assign v$G11_6103_out0 = !(v$SEL3_1239_out0 || v$SEL4_4103_out0);
assign v$G11_6104_out0 = !(v$SEL3_1240_out0 || v$SEL4_4104_out0);
assign v$G11_6111_out0 = !(v$SEL3_1247_out0 || v$SEL4_4111_out0);
assign v$G11_6112_out0 = !(v$SEL3_1248_out0 || v$SEL4_4112_out0);
assign v$G11_6113_out0 = !(v$SEL3_1249_out0 || v$SEL4_4113_out0);
assign v$G11_6114_out0 = !(v$SEL3_1250_out0 || v$SEL4_4114_out0);
assign v$G11_6115_out0 = !(v$SEL3_1251_out0 || v$SEL4_4115_out0);
assign v$G11_6116_out0 = !(v$SEL3_1252_out0 || v$SEL4_4116_out0);
assign v$G11_6117_out0 = !(v$SEL3_1253_out0 || v$SEL4_4117_out0);
assign v$G11_6118_out0 = !(v$SEL3_1254_out0 || v$SEL4_4118_out0);
assign v$G11_6119_out0 = !(v$SEL3_1255_out0 || v$SEL4_4119_out0);
assign v$G11_6120_out0 = !(v$SEL3_1256_out0 || v$SEL4_4120_out0);
assign v$G11_6121_out0 = !(v$SEL3_1257_out0 || v$SEL4_4121_out0);
assign v$G11_6122_out0 = !(v$SEL3_1258_out0 || v$SEL4_4122_out0);
assign v$G11_6123_out0 = !(v$SEL3_1259_out0 || v$SEL4_4123_out0);
assign v$G11_6124_out0 = !(v$SEL3_1260_out0 || v$SEL4_4124_out0);
assign v$G11_6125_out0 = !(v$SEL3_1261_out0 || v$SEL4_4125_out0);
assign v$G11_6126_out0 = !(v$SEL3_1262_out0 || v$SEL4_4126_out0);
assign v$G11_6127_out0 = !(v$SEL3_1263_out0 || v$SEL4_4127_out0);
assign v$G11_6128_out0 = !(v$SEL3_1264_out0 || v$SEL4_4128_out0);
assign v$G11_6129_out0 = !(v$SEL3_1265_out0 || v$SEL4_4129_out0);
assign v$G11_6130_out0 = !(v$SEL3_1266_out0 || v$SEL4_4130_out0);
assign v$G11_6131_out0 = !(v$SEL3_1267_out0 || v$SEL4_4131_out0);
assign v$G11_6132_out0 = !(v$SEL3_1268_out0 || v$SEL4_4132_out0);
assign v$G11_6133_out0 = !(v$SEL3_1269_out0 || v$SEL4_4133_out0);
assign v$G11_6134_out0 = !(v$SEL3_1270_out0 || v$SEL4_4134_out0);
assign v$G8_7762_out0 = ! v$SEL3_1217_out0;
assign v$G8_7763_out0 = ! v$SEL3_1218_out0;
assign v$G8_7764_out0 = ! v$SEL3_1219_out0;
assign v$G8_7765_out0 = ! v$SEL3_1220_out0;
assign v$G8_7766_out0 = ! v$SEL3_1221_out0;
assign v$G8_7767_out0 = ! v$SEL3_1222_out0;
assign v$G8_7768_out0 = ! v$SEL3_1223_out0;
assign v$G8_7769_out0 = ! v$SEL3_1224_out0;
assign v$G8_7770_out0 = ! v$SEL3_1225_out0;
assign v$G8_7771_out0 = ! v$SEL3_1226_out0;
assign v$G8_7772_out0 = ! v$SEL3_1227_out0;
assign v$G8_7773_out0 = ! v$SEL3_1228_out0;
assign v$G8_7774_out0 = ! v$SEL3_1229_out0;
assign v$G8_7775_out0 = ! v$SEL3_1230_out0;
assign v$G8_7776_out0 = ! v$SEL3_1231_out0;
assign v$G8_7777_out0 = ! v$SEL3_1232_out0;
assign v$G8_7778_out0 = ! v$SEL3_1233_out0;
assign v$G8_7779_out0 = ! v$SEL3_1234_out0;
assign v$G8_7780_out0 = ! v$SEL3_1235_out0;
assign v$G8_7781_out0 = ! v$SEL3_1236_out0;
assign v$G8_7782_out0 = ! v$SEL3_1237_out0;
assign v$G8_7783_out0 = ! v$SEL3_1238_out0;
assign v$G8_7784_out0 = ! v$SEL3_1239_out0;
assign v$G8_7785_out0 = ! v$SEL3_1240_out0;
assign v$G8_7792_out0 = ! v$SEL3_1247_out0;
assign v$G8_7793_out0 = ! v$SEL3_1248_out0;
assign v$G8_7794_out0 = ! v$SEL3_1249_out0;
assign v$G8_7795_out0 = ! v$SEL3_1250_out0;
assign v$G8_7796_out0 = ! v$SEL3_1251_out0;
assign v$G8_7797_out0 = ! v$SEL3_1252_out0;
assign v$G8_7798_out0 = ! v$SEL3_1253_out0;
assign v$G8_7799_out0 = ! v$SEL3_1254_out0;
assign v$G8_7800_out0 = ! v$SEL3_1255_out0;
assign v$G8_7801_out0 = ! v$SEL3_1256_out0;
assign v$G8_7802_out0 = ! v$SEL3_1257_out0;
assign v$G8_7803_out0 = ! v$SEL3_1258_out0;
assign v$G8_7804_out0 = ! v$SEL3_1259_out0;
assign v$G8_7805_out0 = ! v$SEL3_1260_out0;
assign v$G8_7806_out0 = ! v$SEL3_1261_out0;
assign v$G8_7807_out0 = ! v$SEL3_1262_out0;
assign v$G8_7808_out0 = ! v$SEL3_1263_out0;
assign v$G8_7809_out0 = ! v$SEL3_1264_out0;
assign v$G8_7810_out0 = ! v$SEL3_1265_out0;
assign v$G8_7811_out0 = ! v$SEL3_1266_out0;
assign v$G8_7812_out0 = ! v$SEL3_1267_out0;
assign v$G8_7813_out0 = ! v$SEL3_1268_out0;
assign v$G8_7814_out0 = ! v$SEL3_1269_out0;
assign v$G8_7815_out0 = ! v$SEL3_1270_out0;
assign v$MUX20_7410_out0 = v$EQ20_6666_out0 ? v$SEL20_5666_out0 : v$MUX21_3294_out0;
assign v$MUX20_7411_out0 = v$EQ20_6667_out0 ? v$SEL20_5667_out0 : v$MUX21_3295_out0;
assign v$MUX20_7412_out0 = v$EQ20_6668_out0 ? v$SEL20_5668_out0 : v$MUX21_3296_out0;
assign v$MUX20_7413_out0 = v$EQ20_6669_out0 ? v$SEL20_5669_out0 : v$MUX21_3297_out0;
assign v$G3_8305_out0 = v$G10_605_out0 && v$G11_6081_out0;
assign v$G3_8306_out0 = v$G10_606_out0 && v$G11_6082_out0;
assign v$G3_8307_out0 = v$G10_607_out0 && v$G11_6083_out0;
assign v$G3_8308_out0 = v$G10_608_out0 && v$G11_6084_out0;
assign v$G3_8309_out0 = v$G10_609_out0 && v$G11_6085_out0;
assign v$G3_8310_out0 = v$G10_610_out0 && v$G11_6086_out0;
assign v$G3_8311_out0 = v$G10_611_out0 && v$G11_6087_out0;
assign v$G3_8312_out0 = v$G10_612_out0 && v$G11_6088_out0;
assign v$G3_8313_out0 = v$G10_613_out0 && v$G11_6089_out0;
assign v$G3_8314_out0 = v$G10_614_out0 && v$G11_6090_out0;
assign v$G3_8315_out0 = v$G10_615_out0 && v$G11_6091_out0;
assign v$G3_8316_out0 = v$G10_616_out0 && v$G11_6092_out0;
assign v$G3_8317_out0 = v$G10_617_out0 && v$G11_6093_out0;
assign v$G3_8318_out0 = v$G10_618_out0 && v$G11_6094_out0;
assign v$G3_8319_out0 = v$G10_619_out0 && v$G11_6095_out0;
assign v$G3_8320_out0 = v$G10_620_out0 && v$G11_6096_out0;
assign v$G3_8321_out0 = v$G10_621_out0 && v$G11_6097_out0;
assign v$G3_8322_out0 = v$G10_622_out0 && v$G11_6098_out0;
assign v$G3_8323_out0 = v$G10_623_out0 && v$G11_6099_out0;
assign v$G3_8324_out0 = v$G10_624_out0 && v$G11_6100_out0;
assign v$G3_8325_out0 = v$G10_625_out0 && v$G11_6101_out0;
assign v$G3_8326_out0 = v$G10_626_out0 && v$G11_6102_out0;
assign v$G3_8327_out0 = v$G10_627_out0 && v$G11_6103_out0;
assign v$G3_8328_out0 = v$G10_628_out0 && v$G11_6104_out0;
assign v$G3_8335_out0 = v$G10_635_out0 && v$G11_6111_out0;
assign v$G3_8336_out0 = v$G10_636_out0 && v$G11_6112_out0;
assign v$G3_8337_out0 = v$G10_637_out0 && v$G11_6113_out0;
assign v$G3_8338_out0 = v$G10_638_out0 && v$G11_6114_out0;
assign v$G3_8339_out0 = v$G10_639_out0 && v$G11_6115_out0;
assign v$G3_8340_out0 = v$G10_640_out0 && v$G11_6116_out0;
assign v$G3_8341_out0 = v$G10_641_out0 && v$G11_6117_out0;
assign v$G3_8342_out0 = v$G10_642_out0 && v$G11_6118_out0;
assign v$G3_8343_out0 = v$G10_643_out0 && v$G11_6119_out0;
assign v$G3_8344_out0 = v$G10_644_out0 && v$G11_6120_out0;
assign v$G3_8345_out0 = v$G10_645_out0 && v$G11_6121_out0;
assign v$G3_8346_out0 = v$G10_646_out0 && v$G11_6122_out0;
assign v$G3_8347_out0 = v$G10_647_out0 && v$G11_6123_out0;
assign v$G3_8348_out0 = v$G10_648_out0 && v$G11_6124_out0;
assign v$G3_8349_out0 = v$G10_649_out0 && v$G11_6125_out0;
assign v$G3_8350_out0 = v$G10_650_out0 && v$G11_6126_out0;
assign v$G3_8351_out0 = v$G10_651_out0 && v$G11_6127_out0;
assign v$G3_8352_out0 = v$G10_652_out0 && v$G11_6128_out0;
assign v$G3_8353_out0 = v$G10_653_out0 && v$G11_6129_out0;
assign v$G3_8354_out0 = v$G10_654_out0 && v$G11_6130_out0;
assign v$G3_8355_out0 = v$G10_655_out0 && v$G11_6131_out0;
assign v$G3_8356_out0 = v$G10_656_out0 && v$G11_6132_out0;
assign v$G3_8357_out0 = v$G10_657_out0 && v$G11_6133_out0;
assign v$G3_8358_out0 = v$G10_658_out0 && v$G11_6134_out0;
assign v$G9_12395_out0 = v$G8_7762_out0 && v$G5_3846_out0;
assign v$G9_12396_out0 = v$G8_7763_out0 && v$G5_3847_out0;
assign v$G9_12397_out0 = v$G8_7764_out0 && v$G5_3848_out0;
assign v$G9_12398_out0 = v$G8_7765_out0 && v$G5_3849_out0;
assign v$G9_12399_out0 = v$G8_7766_out0 && v$G5_3850_out0;
assign v$G9_12400_out0 = v$G8_7767_out0 && v$G5_3851_out0;
assign v$G9_12401_out0 = v$G8_7768_out0 && v$G5_3852_out0;
assign v$G9_12402_out0 = v$G8_7769_out0 && v$G5_3853_out0;
assign v$G9_12403_out0 = v$G8_7770_out0 && v$G5_3854_out0;
assign v$G9_12404_out0 = v$G8_7771_out0 && v$G5_3855_out0;
assign v$G9_12405_out0 = v$G8_7772_out0 && v$G5_3856_out0;
assign v$G9_12406_out0 = v$G8_7773_out0 && v$G5_3857_out0;
assign v$G9_12407_out0 = v$G8_7774_out0 && v$G5_3858_out0;
assign v$G9_12408_out0 = v$G8_7775_out0 && v$G5_3859_out0;
assign v$G9_12409_out0 = v$G8_7776_out0 && v$G5_3860_out0;
assign v$G9_12410_out0 = v$G8_7777_out0 && v$G5_3861_out0;
assign v$G9_12411_out0 = v$G8_7778_out0 && v$G5_3862_out0;
assign v$G9_12412_out0 = v$G8_7779_out0 && v$G5_3863_out0;
assign v$G9_12413_out0 = v$G8_7780_out0 && v$G5_3864_out0;
assign v$G9_12414_out0 = v$G8_7781_out0 && v$G5_3865_out0;
assign v$G9_12415_out0 = v$G8_7782_out0 && v$G5_3866_out0;
assign v$G9_12416_out0 = v$G8_7783_out0 && v$G5_3867_out0;
assign v$G9_12417_out0 = v$G8_7784_out0 && v$G5_3868_out0;
assign v$G9_12418_out0 = v$G8_7785_out0 && v$G5_3869_out0;
assign v$G9_12425_out0 = v$G8_7792_out0 && v$G5_3876_out0;
assign v$G9_12426_out0 = v$G8_7793_out0 && v$G5_3877_out0;
assign v$G9_12427_out0 = v$G8_7794_out0 && v$G5_3878_out0;
assign v$G9_12428_out0 = v$G8_7795_out0 && v$G5_3879_out0;
assign v$G9_12429_out0 = v$G8_7796_out0 && v$G5_3880_out0;
assign v$G9_12430_out0 = v$G8_7797_out0 && v$G5_3881_out0;
assign v$G9_12431_out0 = v$G8_7798_out0 && v$G5_3882_out0;
assign v$G9_12432_out0 = v$G8_7799_out0 && v$G5_3883_out0;
assign v$G9_12433_out0 = v$G8_7800_out0 && v$G5_3884_out0;
assign v$G9_12434_out0 = v$G8_7801_out0 && v$G5_3885_out0;
assign v$G9_12435_out0 = v$G8_7802_out0 && v$G5_3886_out0;
assign v$G9_12436_out0 = v$G8_7803_out0 && v$G5_3887_out0;
assign v$G9_12437_out0 = v$G8_7804_out0 && v$G5_3888_out0;
assign v$G9_12438_out0 = v$G8_7805_out0 && v$G5_3889_out0;
assign v$G9_12439_out0 = v$G8_7806_out0 && v$G5_3890_out0;
assign v$G9_12440_out0 = v$G8_7807_out0 && v$G5_3891_out0;
assign v$G9_12441_out0 = v$G8_7808_out0 && v$G5_3892_out0;
assign v$G9_12442_out0 = v$G8_7809_out0 && v$G5_3893_out0;
assign v$G9_12443_out0 = v$G8_7810_out0 && v$G5_3894_out0;
assign v$G9_12444_out0 = v$G8_7811_out0 && v$G5_3895_out0;
assign v$G9_12445_out0 = v$G8_7812_out0 && v$G5_3896_out0;
assign v$G9_12446_out0 = v$G8_7813_out0 && v$G5_3897_out0;
assign v$G9_12447_out0 = v$G8_7814_out0 && v$G5_3898_out0;
assign v$G9_12448_out0 = v$G8_7815_out0 && v$G5_3899_out0;
assign v$G7_12865_out0 = v$G6_2256_out0 || v$SEL3_1217_out0;
assign v$G7_12866_out0 = v$G6_2257_out0 || v$SEL3_1218_out0;
assign v$G7_12867_out0 = v$G6_2258_out0 || v$SEL3_1219_out0;
assign v$G7_12868_out0 = v$G6_2259_out0 || v$SEL3_1220_out0;
assign v$G7_12869_out0 = v$G6_2260_out0 || v$SEL3_1221_out0;
assign v$G7_12870_out0 = v$G6_2261_out0 || v$SEL3_1222_out0;
assign v$G7_12871_out0 = v$G6_2262_out0 || v$SEL3_1223_out0;
assign v$G7_12872_out0 = v$G6_2263_out0 || v$SEL3_1224_out0;
assign v$G7_12873_out0 = v$G6_2264_out0 || v$SEL3_1225_out0;
assign v$G7_12874_out0 = v$G6_2265_out0 || v$SEL3_1226_out0;
assign v$G7_12875_out0 = v$G6_2266_out0 || v$SEL3_1227_out0;
assign v$G7_12876_out0 = v$G6_2267_out0 || v$SEL3_1228_out0;
assign v$G7_12877_out0 = v$G6_2268_out0 || v$SEL3_1229_out0;
assign v$G7_12878_out0 = v$G6_2269_out0 || v$SEL3_1230_out0;
assign v$G7_12879_out0 = v$G6_2270_out0 || v$SEL3_1231_out0;
assign v$G7_12880_out0 = v$G6_2271_out0 || v$SEL3_1232_out0;
assign v$G7_12881_out0 = v$G6_2272_out0 || v$SEL3_1233_out0;
assign v$G7_12882_out0 = v$G6_2273_out0 || v$SEL3_1234_out0;
assign v$G7_12883_out0 = v$G6_2274_out0 || v$SEL3_1235_out0;
assign v$G7_12884_out0 = v$G6_2275_out0 || v$SEL3_1236_out0;
assign v$G7_12885_out0 = v$G6_2276_out0 || v$SEL3_1237_out0;
assign v$G7_12886_out0 = v$G6_2277_out0 || v$SEL3_1238_out0;
assign v$G7_12887_out0 = v$G6_2278_out0 || v$SEL3_1239_out0;
assign v$G7_12888_out0 = v$G6_2279_out0 || v$SEL3_1240_out0;
assign v$G7_12895_out0 = v$G6_2286_out0 || v$SEL3_1247_out0;
assign v$G7_12896_out0 = v$G6_2287_out0 || v$SEL3_1248_out0;
assign v$G7_12897_out0 = v$G6_2288_out0 || v$SEL3_1249_out0;
assign v$G7_12898_out0 = v$G6_2289_out0 || v$SEL3_1250_out0;
assign v$G7_12899_out0 = v$G6_2290_out0 || v$SEL3_1251_out0;
assign v$G7_12900_out0 = v$G6_2291_out0 || v$SEL3_1252_out0;
assign v$G7_12901_out0 = v$G6_2292_out0 || v$SEL3_1253_out0;
assign v$G7_12902_out0 = v$G6_2293_out0 || v$SEL3_1254_out0;
assign v$G7_12903_out0 = v$G6_2294_out0 || v$SEL3_1255_out0;
assign v$G7_12904_out0 = v$G6_2295_out0 || v$SEL3_1256_out0;
assign v$G7_12905_out0 = v$G6_2296_out0 || v$SEL3_1257_out0;
assign v$G7_12906_out0 = v$G6_2297_out0 || v$SEL3_1258_out0;
assign v$G7_12907_out0 = v$G6_2298_out0 || v$SEL3_1259_out0;
assign v$G7_12908_out0 = v$G6_2299_out0 || v$SEL3_1260_out0;
assign v$G7_12909_out0 = v$G6_2300_out0 || v$SEL3_1261_out0;
assign v$G7_12910_out0 = v$G6_2301_out0 || v$SEL3_1262_out0;
assign v$G7_12911_out0 = v$G6_2302_out0 || v$SEL3_1263_out0;
assign v$G7_12912_out0 = v$G6_2303_out0 || v$SEL3_1264_out0;
assign v$G7_12913_out0 = v$G6_2304_out0 || v$SEL3_1265_out0;
assign v$G7_12914_out0 = v$G6_2305_out0 || v$SEL3_1266_out0;
assign v$G7_12915_out0 = v$G6_2306_out0 || v$SEL3_1267_out0;
assign v$G7_12916_out0 = v$G6_2307_out0 || v$SEL3_1268_out0;
assign v$G7_12917_out0 = v$G6_2308_out0 || v$SEL3_1269_out0;
assign v$G7_12918_out0 = v$G6_2309_out0 || v$SEL3_1270_out0;
assign v$MUX19_4393_out0 = v$EQ19_3689_out0 ? v$SEL19_8464_out0 : v$MUX20_7410_out0;
assign v$MUX19_4394_out0 = v$EQ19_3690_out0 ? v$SEL19_8465_out0 : v$MUX20_7411_out0;
assign v$MUX19_4395_out0 = v$EQ19_3691_out0 ? v$SEL19_8466_out0 : v$MUX20_7412_out0;
assign v$MUX19_4396_out0 = v$EQ19_3692_out0 ? v$SEL19_8467_out0 : v$MUX20_7413_out0;
assign v$Z_8188_out0 = v$G3_8305_out0;
assign v$Z_8189_out0 = v$G3_8306_out0;
assign v$Z_8190_out0 = v$G3_8307_out0;
assign v$Z_8191_out0 = v$G3_8308_out0;
assign v$Z_8192_out0 = v$G3_8309_out0;
assign v$Z_8193_out0 = v$G3_8310_out0;
assign v$Z_8194_out0 = v$G3_8311_out0;
assign v$Z_8195_out0 = v$G3_8312_out0;
assign v$Z_8196_out0 = v$G3_8313_out0;
assign v$Z_8197_out0 = v$G3_8314_out0;
assign v$Z_8198_out0 = v$G3_8315_out0;
assign v$Z_8199_out0 = v$G3_8316_out0;
assign v$Z_8200_out0 = v$G3_8317_out0;
assign v$Z_8201_out0 = v$G3_8318_out0;
assign v$Z_8202_out0 = v$G3_8319_out0;
assign v$Z_8203_out0 = v$G3_8320_out0;
assign v$Z_8204_out0 = v$G3_8321_out0;
assign v$Z_8205_out0 = v$G3_8322_out0;
assign v$Z_8206_out0 = v$G3_8323_out0;
assign v$Z_8207_out0 = v$G3_8324_out0;
assign v$Z_8208_out0 = v$G3_8325_out0;
assign v$Z_8209_out0 = v$G3_8326_out0;
assign v$Z_8210_out0 = v$G3_8327_out0;
assign v$Z_8211_out0 = v$G3_8328_out0;
assign v$Z_8218_out0 = v$G3_8335_out0;
assign v$Z_8219_out0 = v$G3_8336_out0;
assign v$Z_8220_out0 = v$G3_8337_out0;
assign v$Z_8221_out0 = v$G3_8338_out0;
assign v$Z_8222_out0 = v$G3_8339_out0;
assign v$Z_8223_out0 = v$G3_8340_out0;
assign v$Z_8224_out0 = v$G3_8341_out0;
assign v$Z_8225_out0 = v$G3_8342_out0;
assign v$Z_8226_out0 = v$G3_8343_out0;
assign v$Z_8227_out0 = v$G3_8344_out0;
assign v$Z_8228_out0 = v$G3_8345_out0;
assign v$Z_8229_out0 = v$G3_8346_out0;
assign v$Z_8230_out0 = v$G3_8347_out0;
assign v$Z_8231_out0 = v$G3_8348_out0;
assign v$Z_8232_out0 = v$G3_8349_out0;
assign v$Z_8233_out0 = v$G3_8350_out0;
assign v$Z_8234_out0 = v$G3_8351_out0;
assign v$Z_8235_out0 = v$G3_8352_out0;
assign v$Z_8236_out0 = v$G3_8353_out0;
assign v$Z_8237_out0 = v$G3_8354_out0;
assign v$Z_8238_out0 = v$G3_8355_out0;
assign v$Z_8239_out0 = v$G3_8356_out0;
assign v$Z_8240_out0 = v$G3_8357_out0;
assign v$Z_8241_out0 = v$G3_8358_out0;
assign v$G4_12318_out0 = v$G7_12865_out0 && v$G5_3846_out0;
assign v$G4_12319_out0 = v$G7_12866_out0 && v$G5_3847_out0;
assign v$G4_12320_out0 = v$G7_12867_out0 && v$G5_3848_out0;
assign v$G4_12321_out0 = v$G7_12868_out0 && v$G5_3849_out0;
assign v$G4_12322_out0 = v$G7_12869_out0 && v$G5_3850_out0;
assign v$G4_12323_out0 = v$G7_12870_out0 && v$G5_3851_out0;
assign v$G4_12324_out0 = v$G7_12871_out0 && v$G5_3852_out0;
assign v$G4_12325_out0 = v$G7_12872_out0 && v$G5_3853_out0;
assign v$G4_12326_out0 = v$G7_12873_out0 && v$G5_3854_out0;
assign v$G4_12327_out0 = v$G7_12874_out0 && v$G5_3855_out0;
assign v$G4_12328_out0 = v$G7_12875_out0 && v$G5_3856_out0;
assign v$G4_12329_out0 = v$G7_12876_out0 && v$G5_3857_out0;
assign v$G4_12330_out0 = v$G7_12877_out0 && v$G5_3858_out0;
assign v$G4_12331_out0 = v$G7_12878_out0 && v$G5_3859_out0;
assign v$G4_12332_out0 = v$G7_12879_out0 && v$G5_3860_out0;
assign v$G4_12333_out0 = v$G7_12880_out0 && v$G5_3861_out0;
assign v$G4_12334_out0 = v$G7_12881_out0 && v$G5_3862_out0;
assign v$G4_12335_out0 = v$G7_12882_out0 && v$G5_3863_out0;
assign v$G4_12336_out0 = v$G7_12883_out0 && v$G5_3864_out0;
assign v$G4_12337_out0 = v$G7_12884_out0 && v$G5_3865_out0;
assign v$G4_12338_out0 = v$G7_12885_out0 && v$G5_3866_out0;
assign v$G4_12339_out0 = v$G7_12886_out0 && v$G5_3867_out0;
assign v$G4_12340_out0 = v$G7_12887_out0 && v$G5_3868_out0;
assign v$G4_12341_out0 = v$G7_12888_out0 && v$G5_3869_out0;
assign v$G4_12348_out0 = v$G7_12895_out0 && v$G5_3876_out0;
assign v$G4_12349_out0 = v$G7_12896_out0 && v$G5_3877_out0;
assign v$G4_12350_out0 = v$G7_12897_out0 && v$G5_3878_out0;
assign v$G4_12351_out0 = v$G7_12898_out0 && v$G5_3879_out0;
assign v$G4_12352_out0 = v$G7_12899_out0 && v$G5_3880_out0;
assign v$G4_12353_out0 = v$G7_12900_out0 && v$G5_3881_out0;
assign v$G4_12354_out0 = v$G7_12901_out0 && v$G5_3882_out0;
assign v$G4_12355_out0 = v$G7_12902_out0 && v$G5_3883_out0;
assign v$G4_12356_out0 = v$G7_12903_out0 && v$G5_3884_out0;
assign v$G4_12357_out0 = v$G7_12904_out0 && v$G5_3885_out0;
assign v$G4_12358_out0 = v$G7_12905_out0 && v$G5_3886_out0;
assign v$G4_12359_out0 = v$G7_12906_out0 && v$G5_3887_out0;
assign v$G4_12360_out0 = v$G7_12907_out0 && v$G5_3888_out0;
assign v$G4_12361_out0 = v$G7_12908_out0 && v$G5_3889_out0;
assign v$G4_12362_out0 = v$G7_12909_out0 && v$G5_3890_out0;
assign v$G4_12363_out0 = v$G7_12910_out0 && v$G5_3891_out0;
assign v$G4_12364_out0 = v$G7_12911_out0 && v$G5_3892_out0;
assign v$G4_12365_out0 = v$G7_12912_out0 && v$G5_3893_out0;
assign v$G4_12366_out0 = v$G7_12913_out0 && v$G5_3894_out0;
assign v$G4_12367_out0 = v$G7_12914_out0 && v$G5_3895_out0;
assign v$G4_12368_out0 = v$G7_12915_out0 && v$G5_3896_out0;
assign v$G4_12369_out0 = v$G7_12916_out0 && v$G5_3897_out0;
assign v$G4_12370_out0 = v$G7_12917_out0 && v$G5_3898_out0;
assign v$G4_12371_out0 = v$G7_12918_out0 && v$G5_3899_out0;
assign v$MUX18_3258_out0 = v$EQ18_8460_out0 ? v$SEL18_7420_out0 : v$MUX19_4393_out0;
assign v$MUX18_3259_out0 = v$EQ18_8461_out0 ? v$SEL18_7421_out0 : v$MUX19_4394_out0;
assign v$MUX18_3260_out0 = v$EQ18_8462_out0 ? v$SEL18_7422_out0 : v$MUX19_4395_out0;
assign v$MUX18_3261_out0 = v$EQ18_8463_out0 ? v$SEL18_7423_out0 : v$MUX19_4396_out0;
assign v$_4267_out0 = { v$G4_12318_out0,v$G9_12395_out0 };
assign v$_4268_out0 = { v$G4_12319_out0,v$G9_12396_out0 };
assign v$_4269_out0 = { v$G4_12320_out0,v$G9_12397_out0 };
assign v$_4270_out0 = { v$G4_12321_out0,v$G9_12398_out0 };
assign v$_4271_out0 = { v$G4_12322_out0,v$G9_12399_out0 };
assign v$_4272_out0 = { v$G4_12323_out0,v$G9_12400_out0 };
assign v$_4273_out0 = { v$G4_12324_out0,v$G9_12401_out0 };
assign v$_4274_out0 = { v$G4_12325_out0,v$G9_12402_out0 };
assign v$_4275_out0 = { v$G4_12326_out0,v$G9_12403_out0 };
assign v$_4276_out0 = { v$G4_12327_out0,v$G9_12404_out0 };
assign v$_4277_out0 = { v$G4_12328_out0,v$G9_12405_out0 };
assign v$_4278_out0 = { v$G4_12329_out0,v$G9_12406_out0 };
assign v$_4279_out0 = { v$G4_12330_out0,v$G9_12407_out0 };
assign v$_4280_out0 = { v$G4_12331_out0,v$G9_12408_out0 };
assign v$_4281_out0 = { v$G4_12332_out0,v$G9_12409_out0 };
assign v$_4282_out0 = { v$G4_12333_out0,v$G9_12410_out0 };
assign v$_4283_out0 = { v$G4_12334_out0,v$G9_12411_out0 };
assign v$_4284_out0 = { v$G4_12335_out0,v$G9_12412_out0 };
assign v$_4285_out0 = { v$G4_12336_out0,v$G9_12413_out0 };
assign v$_4286_out0 = { v$G4_12337_out0,v$G9_12414_out0 };
assign v$_4287_out0 = { v$G4_12338_out0,v$G9_12415_out0 };
assign v$_4288_out0 = { v$G4_12339_out0,v$G9_12416_out0 };
assign v$_4289_out0 = { v$G4_12340_out0,v$G9_12417_out0 };
assign v$_4290_out0 = { v$G4_12341_out0,v$G9_12418_out0 };
assign v$_4297_out0 = { v$G4_12348_out0,v$G9_12425_out0 };
assign v$_4298_out0 = { v$G4_12349_out0,v$G9_12426_out0 };
assign v$_4299_out0 = { v$G4_12350_out0,v$G9_12427_out0 };
assign v$_4300_out0 = { v$G4_12351_out0,v$G9_12428_out0 };
assign v$_4301_out0 = { v$G4_12352_out0,v$G9_12429_out0 };
assign v$_4302_out0 = { v$G4_12353_out0,v$G9_12430_out0 };
assign v$_4303_out0 = { v$G4_12354_out0,v$G9_12431_out0 };
assign v$_4304_out0 = { v$G4_12355_out0,v$G9_12432_out0 };
assign v$_4305_out0 = { v$G4_12356_out0,v$G9_12433_out0 };
assign v$_4306_out0 = { v$G4_12357_out0,v$G9_12434_out0 };
assign v$_4307_out0 = { v$G4_12358_out0,v$G9_12435_out0 };
assign v$_4308_out0 = { v$G4_12359_out0,v$G9_12436_out0 };
assign v$_4309_out0 = { v$G4_12360_out0,v$G9_12437_out0 };
assign v$_4310_out0 = { v$G4_12361_out0,v$G9_12438_out0 };
assign v$_4311_out0 = { v$G4_12362_out0,v$G9_12439_out0 };
assign v$_4312_out0 = { v$G4_12363_out0,v$G9_12440_out0 };
assign v$_4313_out0 = { v$G4_12364_out0,v$G9_12441_out0 };
assign v$_4314_out0 = { v$G4_12365_out0,v$G9_12442_out0 };
assign v$_4315_out0 = { v$G4_12366_out0,v$G9_12443_out0 };
assign v$_4316_out0 = { v$G4_12367_out0,v$G9_12444_out0 };
assign v$_4317_out0 = { v$G4_12368_out0,v$G9_12445_out0 };
assign v$_4318_out0 = { v$G4_12369_out0,v$G9_12446_out0 };
assign v$_4319_out0 = { v$G4_12370_out0,v$G9_12447_out0 };
assign v$_4320_out0 = { v$G4_12371_out0,v$G9_12448_out0 };
assign v$Z2_4334_out0 = v$Z_8190_out0;
assign v$Z2_4335_out0 = v$Z_8194_out0;
assign v$Z2_4336_out0 = v$Z_8198_out0;
assign v$Z2_4338_out0 = v$Z_8202_out0;
assign v$Z2_4339_out0 = v$Z_8206_out0;
assign v$Z2_4340_out0 = v$Z_8210_out0;
assign v$Z2_4342_out0 = v$Z_8220_out0;
assign v$Z2_4343_out0 = v$Z_8224_out0;
assign v$Z2_4344_out0 = v$Z_8228_out0;
assign v$Z2_4346_out0 = v$Z_8232_out0;
assign v$Z2_4347_out0 = v$Z_8236_out0;
assign v$Z2_4348_out0 = v$Z_8240_out0;
assign v$Z4_5426_out0 = v$Z_8191_out0;
assign v$Z4_5427_out0 = v$Z_8195_out0;
assign v$Z4_5428_out0 = v$Z_8199_out0;
assign v$Z4_5429_out0 = v$Z_8203_out0;
assign v$Z4_5430_out0 = v$Z_8207_out0;
assign v$Z4_5431_out0 = v$Z_8211_out0;
assign v$Z4_5432_out0 = v$Z_8221_out0;
assign v$Z4_5433_out0 = v$Z_8225_out0;
assign v$Z4_5434_out0 = v$Z_8229_out0;
assign v$Z4_5435_out0 = v$Z_8233_out0;
assign v$Z4_5436_out0 = v$Z_8237_out0;
assign v$Z4_5437_out0 = v$Z_8241_out0;
assign v$Z1_12049_out0 = v$Z_8189_out0;
assign v$Z1_12050_out0 = v$Z_8193_out0;
assign v$Z1_12051_out0 = v$Z_8197_out0;
assign v$Z1_12053_out0 = v$Z_8201_out0;
assign v$Z1_12054_out0 = v$Z_8205_out0;
assign v$Z1_12055_out0 = v$Z_8209_out0;
assign v$Z1_12057_out0 = v$Z_8219_out0;
assign v$Z1_12058_out0 = v$Z_8223_out0;
assign v$Z1_12059_out0 = v$Z_8227_out0;
assign v$Z1_12061_out0 = v$Z_8231_out0;
assign v$Z1_12062_out0 = v$Z_8235_out0;
assign v$Z1_12063_out0 = v$Z_8239_out0;
assign v$Z3_12568_out0 = v$Z_8188_out0;
assign v$Z3_12569_out0 = v$Z_8192_out0;
assign v$Z3_12570_out0 = v$Z_8196_out0;
assign v$Z3_12572_out0 = v$Z_8200_out0;
assign v$Z3_12573_out0 = v$Z_8204_out0;
assign v$Z3_12574_out0 = v$Z_8208_out0;
assign v$Z3_12576_out0 = v$Z_8218_out0;
assign v$Z3_12577_out0 = v$Z_8222_out0;
assign v$Z3_12578_out0 = v$Z_8226_out0;
assign v$Z3_12580_out0 = v$Z_8230_out0;
assign v$Z3_12581_out0 = v$Z_8234_out0;
assign v$Z3_12582_out0 = v$Z_8238_out0;
assign v$G4_4055_out0 = ! v$Z4_5426_out0;
assign v$G4_4056_out0 = ! v$Z4_5427_out0;
assign v$G4_4057_out0 = ! v$Z4_5428_out0;
assign v$G4_4058_out0 = ! v$Z4_5429_out0;
assign v$G4_4059_out0 = ! v$Z4_5430_out0;
assign v$G4_4060_out0 = ! v$Z4_5431_out0;
assign v$G4_4061_out0 = ! v$Z4_5432_out0;
assign v$G4_4062_out0 = ! v$Z4_5433_out0;
assign v$G4_4063_out0 = ! v$Z4_5434_out0;
assign v$G4_4064_out0 = ! v$Z4_5435_out0;
assign v$G4_4065_out0 = ! v$Z4_5436_out0;
assign v$G4_4066_out0 = ! v$Z4_5437_out0;
assign v$G6_4184_out0 = ! v$Z2_4334_out0;
assign v$G6_4185_out0 = ! v$Z2_4335_out0;
assign v$G6_4186_out0 = ! v$Z2_4336_out0;
assign v$G6_4188_out0 = ! v$Z2_4338_out0;
assign v$G6_4189_out0 = ! v$Z2_4339_out0;
assign v$G6_4190_out0 = ! v$Z2_4340_out0;
assign v$G6_4192_out0 = ! v$Z2_4342_out0;
assign v$G6_4193_out0 = ! v$Z2_4343_out0;
assign v$G6_4194_out0 = ! v$Z2_4344_out0;
assign v$G6_4196_out0 = ! v$Z2_4346_out0;
assign v$G6_4197_out0 = ! v$Z2_4347_out0;
assign v$G6_4198_out0 = ! v$Z2_4348_out0;
assign v$Y_4474_out0 = v$_4267_out0;
assign v$Y_4475_out0 = v$_4268_out0;
assign v$Y_4476_out0 = v$_4269_out0;
assign v$Y_4477_out0 = v$_4270_out0;
assign v$Y_4478_out0 = v$_4271_out0;
assign v$Y_4479_out0 = v$_4272_out0;
assign v$Y_4480_out0 = v$_4273_out0;
assign v$Y_4481_out0 = v$_4274_out0;
assign v$Y_4482_out0 = v$_4275_out0;
assign v$Y_4483_out0 = v$_4276_out0;
assign v$Y_4484_out0 = v$_4277_out0;
assign v$Y_4485_out0 = v$_4278_out0;
assign v$Y_4486_out0 = v$_4279_out0;
assign v$Y_4487_out0 = v$_4280_out0;
assign v$Y_4488_out0 = v$_4281_out0;
assign v$Y_4489_out0 = v$_4282_out0;
assign v$Y_4490_out0 = v$_4283_out0;
assign v$Y_4491_out0 = v$_4284_out0;
assign v$Y_4492_out0 = v$_4285_out0;
assign v$Y_4493_out0 = v$_4286_out0;
assign v$Y_4494_out0 = v$_4287_out0;
assign v$Y_4495_out0 = v$_4288_out0;
assign v$Y_4496_out0 = v$_4289_out0;
assign v$Y_4497_out0 = v$_4290_out0;
assign v$Y_4504_out0 = v$_4297_out0;
assign v$Y_4505_out0 = v$_4298_out0;
assign v$Y_4506_out0 = v$_4299_out0;
assign v$Y_4507_out0 = v$_4300_out0;
assign v$Y_4508_out0 = v$_4301_out0;
assign v$Y_4509_out0 = v$_4302_out0;
assign v$Y_4510_out0 = v$_4303_out0;
assign v$Y_4511_out0 = v$_4304_out0;
assign v$Y_4512_out0 = v$_4305_out0;
assign v$Y_4513_out0 = v$_4306_out0;
assign v$Y_4514_out0 = v$_4307_out0;
assign v$Y_4515_out0 = v$_4308_out0;
assign v$Y_4516_out0 = v$_4309_out0;
assign v$Y_4517_out0 = v$_4310_out0;
assign v$Y_4518_out0 = v$_4311_out0;
assign v$Y_4519_out0 = v$_4312_out0;
assign v$Y_4520_out0 = v$_4313_out0;
assign v$Y_4521_out0 = v$_4314_out0;
assign v$Y_4522_out0 = v$_4315_out0;
assign v$Y_4523_out0 = v$_4316_out0;
assign v$Y_4524_out0 = v$_4317_out0;
assign v$Y_4525_out0 = v$_4318_out0;
assign v$Y_4526_out0 = v$_4319_out0;
assign v$Y_4527_out0 = v$_4320_out0;
assign v$G9_10504_out0 = v$Z1_12049_out0 && v$Z2_4334_out0;
assign v$G9_10505_out0 = v$Z1_12050_out0 && v$Z2_4335_out0;
assign v$G9_10506_out0 = v$Z1_12051_out0 && v$Z2_4336_out0;
assign v$G9_10508_out0 = v$Z1_12053_out0 && v$Z2_4338_out0;
assign v$G9_10509_out0 = v$Z1_12054_out0 && v$Z2_4339_out0;
assign v$G9_10510_out0 = v$Z1_12055_out0 && v$Z2_4340_out0;
assign v$G9_10512_out0 = v$Z1_12057_out0 && v$Z2_4342_out0;
assign v$G9_10513_out0 = v$Z1_12058_out0 && v$Z2_4343_out0;
assign v$G9_10514_out0 = v$Z1_12059_out0 && v$Z2_4344_out0;
assign v$G9_10516_out0 = v$Z1_12061_out0 && v$Z2_4346_out0;
assign v$G9_10517_out0 = v$Z1_12062_out0 && v$Z2_4347_out0;
assign v$G9_10518_out0 = v$Z1_12063_out0 && v$Z2_4348_out0;
assign v$MUX17_11616_out0 = v$EQ17_3906_out0 ? v$SEL17_11249_out0 : v$MUX18_3258_out0;
assign v$MUX17_11617_out0 = v$EQ17_3907_out0 ? v$SEL17_11250_out0 : v$MUX18_3259_out0;
assign v$MUX17_11618_out0 = v$EQ17_3908_out0 ? v$SEL17_11251_out0 : v$MUX18_3260_out0;
assign v$MUX17_11619_out0 = v$EQ17_3909_out0 ? v$SEL17_11252_out0 : v$MUX18_3261_out0;
assign v$G5_12296_out0 = ! v$Z3_12568_out0;
assign v$G5_12297_out0 = ! v$Z3_12569_out0;
assign v$G5_12298_out0 = ! v$Z3_12570_out0;
assign v$G5_12299_out0 = ! v$Z3_12572_out0;
assign v$G5_12300_out0 = ! v$Z3_12573_out0;
assign v$G5_12301_out0 = ! v$Z3_12574_out0;
assign v$G5_12302_out0 = ! v$Z3_12576_out0;
assign v$G5_12303_out0 = ! v$Z3_12577_out0;
assign v$G5_12304_out0 = ! v$Z3_12578_out0;
assign v$G5_12305_out0 = ! v$Z3_12580_out0;
assign v$G5_12306_out0 = ! v$Z3_12581_out0;
assign v$G5_12307_out0 = ! v$Z3_12582_out0;
assign v$_2700_out0 = { v$Y_4477_out0,v$C3_2001_out0 };
assign v$_2701_out0 = { v$Y_4481_out0,v$C3_2002_out0 };
assign v$_2702_out0 = { v$Y_4485_out0,v$C3_2003_out0 };
assign v$_2703_out0 = { v$Y_4489_out0,v$C3_2004_out0 };
assign v$_2704_out0 = { v$Y_4493_out0,v$C3_2005_out0 };
assign v$_2705_out0 = { v$Y_4497_out0,v$C3_2006_out0 };
assign v$_2706_out0 = { v$Y_4507_out0,v$C3_2007_out0 };
assign v$_2707_out0 = { v$Y_4511_out0,v$C3_2008_out0 };
assign v$_2708_out0 = { v$Y_4515_out0,v$C3_2009_out0 };
assign v$_2709_out0 = { v$Y_4519_out0,v$C3_2010_out0 };
assign v$_2710_out0 = { v$Y_4523_out0,v$C3_2011_out0 };
assign v$_2711_out0 = { v$Y_4527_out0,v$C3_2012_out0 };
assign v$_3462_out0 = { v$Y_4476_out0,v$C5_11958_out0 };
assign v$_3463_out0 = { v$Y_4480_out0,v$C5_11959_out0 };
assign v$_3464_out0 = { v$Y_4484_out0,v$C5_11960_out0 };
assign v$_3466_out0 = { v$Y_4488_out0,v$C5_11962_out0 };
assign v$_3467_out0 = { v$Y_4492_out0,v$C5_11963_out0 };
assign v$_3468_out0 = { v$Y_4496_out0,v$C5_11964_out0 };
assign v$_3470_out0 = { v$Y_4506_out0,v$C5_11966_out0 };
assign v$_3471_out0 = { v$Y_4510_out0,v$C5_11967_out0 };
assign v$_3472_out0 = { v$Y_4514_out0,v$C5_11968_out0 };
assign v$_3474_out0 = { v$Y_4518_out0,v$C5_11970_out0 };
assign v$_3475_out0 = { v$Y_4522_out0,v$C5_11971_out0 };
assign v$_3476_out0 = { v$Y_4526_out0,v$C5_11972_out0 };
assign v$_6022_out0 = { v$Y_4475_out0,v$C6_4537_out0 };
assign v$_6023_out0 = { v$Y_4479_out0,v$C6_4538_out0 };
assign v$_6024_out0 = { v$Y_4483_out0,v$C6_4539_out0 };
assign v$_6026_out0 = { v$Y_4487_out0,v$C6_4541_out0 };
assign v$_6027_out0 = { v$Y_4491_out0,v$C6_4542_out0 };
assign v$_6028_out0 = { v$Y_4495_out0,v$C6_4543_out0 };
assign v$_6030_out0 = { v$Y_4505_out0,v$C6_4545_out0 };
assign v$_6031_out0 = { v$Y_4509_out0,v$C6_4546_out0 };
assign v$_6032_out0 = { v$Y_4513_out0,v$C6_4547_out0 };
assign v$_6034_out0 = { v$Y_4517_out0,v$C6_4549_out0 };
assign v$_6035_out0 = { v$Y_4521_out0,v$C6_4550_out0 };
assign v$_6036_out0 = { v$Y_4525_out0,v$C6_4551_out0 };
assign v$_6148_out0 = { v$Y_4474_out0,v$C4_11589_out0 };
assign v$_6149_out0 = { v$Y_4478_out0,v$C4_11590_out0 };
assign v$_6150_out0 = { v$Y_4482_out0,v$C4_11591_out0 };
assign v$_6152_out0 = { v$Y_4486_out0,v$C4_11593_out0 };
assign v$_6153_out0 = { v$Y_4490_out0,v$C4_11594_out0 };
assign v$_6154_out0 = { v$Y_4494_out0,v$C4_11595_out0 };
assign v$_6156_out0 = { v$Y_4504_out0,v$C4_11597_out0 };
assign v$_6157_out0 = { v$Y_4508_out0,v$C4_11598_out0 };
assign v$_6158_out0 = { v$Y_4512_out0,v$C4_11599_out0 };
assign v$_6160_out0 = { v$Y_4516_out0,v$C4_11601_out0 };
assign v$_6161_out0 = { v$Y_4520_out0,v$C4_11602_out0 };
assign v$_6162_out0 = { v$Y_4524_out0,v$C4_11603_out0 };
assign v$G7_6594_out0 = v$G9_10504_out0 && v$Z3_12568_out0;
assign v$G7_6595_out0 = v$G9_10505_out0 && v$Z3_12569_out0;
assign v$G7_6596_out0 = v$G9_10506_out0 && v$Z3_12570_out0;
assign v$G7_6598_out0 = v$G9_10508_out0 && v$Z3_12572_out0;
assign v$G7_6599_out0 = v$G9_10509_out0 && v$Z3_12573_out0;
assign v$G7_6600_out0 = v$G9_10510_out0 && v$Z3_12574_out0;
assign v$G7_6602_out0 = v$G9_10512_out0 && v$Z3_12576_out0;
assign v$G7_6603_out0 = v$G9_10513_out0 && v$Z3_12577_out0;
assign v$G7_6604_out0 = v$G9_10514_out0 && v$Z3_12578_out0;
assign v$G7_6606_out0 = v$G9_10516_out0 && v$Z3_12580_out0;
assign v$G7_6607_out0 = v$G9_10517_out0 && v$Z3_12581_out0;
assign v$G7_6608_out0 = v$G9_10518_out0 && v$Z3_12582_out0;
assign v$MUX16_11809_out0 = v$EQ16_5760_out0 ? v$SEL16_11943_out0 : v$MUX17_11616_out0;
assign v$MUX16_11810_out0 = v$EQ16_5761_out0 ? v$SEL16_11944_out0 : v$MUX17_11617_out0;
assign v$MUX16_11811_out0 = v$EQ16_5762_out0 ? v$SEL16_11945_out0 : v$MUX17_11618_out0;
assign v$MUX16_11812_out0 = v$EQ16_5763_out0 ? v$SEL16_11946_out0 : v$MUX17_11619_out0;
assign v$MUX5_2765_out0 = v$G6_4184_out0 ? v$_3462_out0 : v$_6022_out0;
assign v$MUX5_2766_out0 = v$G6_4185_out0 ? v$_3463_out0 : v$_6023_out0;
assign v$MUX5_2767_out0 = v$G6_4186_out0 ? v$_3464_out0 : v$_6024_out0;
assign v$MUX5_2769_out0 = v$G6_4188_out0 ? v$_3466_out0 : v$_6026_out0;
assign v$MUX5_2770_out0 = v$G6_4189_out0 ? v$_3467_out0 : v$_6027_out0;
assign v$MUX5_2771_out0 = v$G6_4190_out0 ? v$_3468_out0 : v$_6028_out0;
assign v$MUX5_2773_out0 = v$G6_4192_out0 ? v$_3470_out0 : v$_6030_out0;
assign v$MUX5_2774_out0 = v$G6_4193_out0 ? v$_3471_out0 : v$_6031_out0;
assign v$MUX5_2775_out0 = v$G6_4194_out0 ? v$_3472_out0 : v$_6032_out0;
assign v$MUX5_2777_out0 = v$G6_4196_out0 ? v$_3474_out0 : v$_6034_out0;
assign v$MUX5_2778_out0 = v$G6_4197_out0 ? v$_3475_out0 : v$_6035_out0;
assign v$MUX5_2779_out0 = v$G6_4198_out0 ? v$_3476_out0 : v$_6036_out0;
assign v$LOWER$PART_4327_out0 = v$MUX16_11809_out0;
assign v$LOWER$PART_4328_out0 = v$MUX16_11810_out0;
assign v$LOWER$PART_4329_out0 = v$MUX16_11811_out0;
assign v$LOWER$PART_4330_out0 = v$MUX16_11812_out0;
assign v$G1_11306_out0 = v$G7_6594_out0 && v$Z4_5426_out0;
assign v$G1_11307_out0 = v$G7_6595_out0 && v$Z4_5427_out0;
assign v$G1_11308_out0 = v$G7_6596_out0 && v$Z4_5428_out0;
assign v$G1_11309_out0 = v$G7_6598_out0 && v$Z4_5429_out0;
assign v$G1_11310_out0 = v$G7_6599_out0 && v$Z4_5430_out0;
assign v$G1_11311_out0 = v$G7_6600_out0 && v$Z4_5431_out0;
assign v$G1_11312_out0 = v$G7_6602_out0 && v$Z4_5432_out0;
assign v$G1_11313_out0 = v$G7_6603_out0 && v$Z4_5433_out0;
assign v$G1_11314_out0 = v$G7_6604_out0 && v$Z4_5434_out0;
assign v$G1_11315_out0 = v$G7_6606_out0 && v$Z4_5435_out0;
assign v$G1_11316_out0 = v$G7_6607_out0 && v$Z4_5436_out0;
assign v$G1_11317_out0 = v$G7_6608_out0 && v$Z4_5437_out0;
assign v$MUX15_547_out0 = v$EQ15_11158_out0 ? v$SEL15_3278_out0 : v$LOWER$PART_4327_out0;
assign v$MUX15_548_out0 = v$EQ15_11159_out0 ? v$SEL15_3279_out0 : v$LOWER$PART_4328_out0;
assign v$MUX15_549_out0 = v$EQ15_11160_out0 ? v$SEL15_3280_out0 : v$LOWER$PART_4329_out0;
assign v$MUX15_550_out0 = v$EQ15_11161_out0 ? v$SEL15_3281_out0 : v$LOWER$PART_4330_out0;
assign v$Z_1461_out0 = v$G1_11306_out0;
assign v$Z_1462_out0 = v$G1_11307_out0;
assign v$Z_1463_out0 = v$G1_11308_out0;
assign v$Z_1465_out0 = v$G1_11309_out0;
assign v$Z_1466_out0 = v$G1_11310_out0;
assign v$Z_1467_out0 = v$G1_11311_out0;
assign v$Z_1469_out0 = v$G1_11312_out0;
assign v$Z_1470_out0 = v$G1_11313_out0;
assign v$Z_1471_out0 = v$G1_11314_out0;
assign v$Z_1473_out0 = v$G1_11315_out0;
assign v$Z_1474_out0 = v$G1_11316_out0;
assign v$Z_1475_out0 = v$G1_11317_out0;
assign v$MUX4_1642_out0 = v$G5_12296_out0 ? v$_6148_out0 : v$MUX5_2765_out0;
assign v$MUX4_1643_out0 = v$G5_12297_out0 ? v$_6149_out0 : v$MUX5_2766_out0;
assign v$MUX4_1644_out0 = v$G5_12298_out0 ? v$_6150_out0 : v$MUX5_2767_out0;
assign v$MUX4_1646_out0 = v$G5_12299_out0 ? v$_6152_out0 : v$MUX5_2769_out0;
assign v$MUX4_1647_out0 = v$G5_12300_out0 ? v$_6153_out0 : v$MUX5_2770_out0;
assign v$MUX4_1648_out0 = v$G5_12301_out0 ? v$_6154_out0 : v$MUX5_2771_out0;
assign v$MUX4_1650_out0 = v$G5_12302_out0 ? v$_6156_out0 : v$MUX5_2773_out0;
assign v$MUX4_1651_out0 = v$G5_12303_out0 ? v$_6157_out0 : v$MUX5_2774_out0;
assign v$MUX4_1652_out0 = v$G5_12304_out0 ? v$_6158_out0 : v$MUX5_2775_out0;
assign v$MUX4_1654_out0 = v$G5_12305_out0 ? v$_6160_out0 : v$MUX5_2777_out0;
assign v$MUX4_1655_out0 = v$G5_12306_out0 ? v$_6161_out0 : v$MUX5_2778_out0;
assign v$MUX4_1656_out0 = v$G5_12307_out0 ? v$_6162_out0 : v$MUX5_2779_out0;
assign v$MUX14_3312_out0 = v$EQ14_3647_out0 ? v$SEL14_11462_out0 : v$MUX15_547_out0;
assign v$MUX14_3313_out0 = v$EQ14_3648_out0 ? v$SEL14_11463_out0 : v$MUX15_548_out0;
assign v$MUX14_3314_out0 = v$EQ14_3649_out0 ? v$SEL14_11464_out0 : v$MUX15_549_out0;
assign v$MUX14_3315_out0 = v$EQ14_3650_out0 ? v$SEL14_11465_out0 : v$MUX15_550_out0;
assign v$Z2_4333_out0 = v$Z_1462_out0;
assign v$Z2_4337_out0 = v$Z_1466_out0;
assign v$Z2_4341_out0 = v$Z_1470_out0;
assign v$Z2_4345_out0 = v$Z_1474_out0;
assign v$Z1_12048_out0 = v$Z_1461_out0;
assign v$Z1_12052_out0 = v$Z_1465_out0;
assign v$Z1_12056_out0 = v$Z_1469_out0;
assign v$Z1_12060_out0 = v$Z_1473_out0;
assign v$MUX3_12264_out0 = v$G4_4055_out0 ? v$_2700_out0 : v$MUX4_1642_out0;
assign v$MUX3_12265_out0 = v$G4_4056_out0 ? v$_2701_out0 : v$MUX4_1643_out0;
assign v$MUX3_12266_out0 = v$G4_4057_out0 ? v$_2702_out0 : v$MUX4_1644_out0;
assign v$MUX3_12267_out0 = v$G4_4058_out0 ? v$_2703_out0 : v$MUX4_1646_out0;
assign v$MUX3_12268_out0 = v$G4_4059_out0 ? v$_2704_out0 : v$MUX4_1647_out0;
assign v$MUX3_12269_out0 = v$G4_4060_out0 ? v$_2705_out0 : v$MUX4_1648_out0;
assign v$MUX3_12270_out0 = v$G4_4061_out0 ? v$_2706_out0 : v$MUX4_1650_out0;
assign v$MUX3_12271_out0 = v$G4_4062_out0 ? v$_2707_out0 : v$MUX4_1651_out0;
assign v$MUX3_12272_out0 = v$G4_4063_out0 ? v$_2708_out0 : v$MUX4_1652_out0;
assign v$MUX3_12273_out0 = v$G4_4064_out0 ? v$_2709_out0 : v$MUX4_1654_out0;
assign v$MUX3_12274_out0 = v$G4_4065_out0 ? v$_2710_out0 : v$MUX4_1655_out0;
assign v$MUX3_12275_out0 = v$G4_4066_out0 ? v$_2711_out0 : v$MUX4_1656_out0;
assign v$Z3_12567_out0 = v$Z_1463_out0;
assign v$Z3_12571_out0 = v$Z_1467_out0;
assign v$Z3_12575_out0 = v$Z_1471_out0;
assign v$Z3_12579_out0 = v$Z_1475_out0;
assign v$G6_4183_out0 = ! v$Z2_4333_out0;
assign v$G6_4187_out0 = ! v$Z2_4337_out0;
assign v$G6_4191_out0 = ! v$Z2_4341_out0;
assign v$G6_4195_out0 = ! v$Z2_4345_out0;
assign v$OUT_6200_out0 = v$MUX3_12264_out0;
assign v$OUT_6201_out0 = v$MUX3_12265_out0;
assign v$OUT_6202_out0 = v$MUX3_12266_out0;
assign v$OUT_6204_out0 = v$MUX3_12267_out0;
assign v$OUT_6205_out0 = v$MUX3_12268_out0;
assign v$OUT_6206_out0 = v$MUX3_12269_out0;
assign v$OUT_6208_out0 = v$MUX3_12270_out0;
assign v$OUT_6209_out0 = v$MUX3_12271_out0;
assign v$OUT_6210_out0 = v$MUX3_12272_out0;
assign v$OUT_6212_out0 = v$MUX3_12273_out0;
assign v$OUT_6213_out0 = v$MUX3_12274_out0;
assign v$OUT_6214_out0 = v$MUX3_12275_out0;
assign v$MUX13_9228_out0 = v$EQ13_6491_out0 ? v$SEL13_4694_out0 : v$MUX14_3312_out0;
assign v$MUX13_9229_out0 = v$EQ13_6492_out0 ? v$SEL13_4695_out0 : v$MUX14_3313_out0;
assign v$MUX13_9230_out0 = v$EQ13_6493_out0 ? v$SEL13_4696_out0 : v$MUX14_3314_out0;
assign v$MUX13_9231_out0 = v$EQ13_6494_out0 ? v$SEL13_4697_out0 : v$MUX14_3315_out0;
assign v$G9_10503_out0 = v$Z1_12048_out0 && v$Z2_4333_out0;
assign v$G9_10507_out0 = v$Z1_12052_out0 && v$Z2_4337_out0;
assign v$G9_10511_out0 = v$Z1_12056_out0 && v$Z2_4341_out0;
assign v$G9_10515_out0 = v$Z1_12060_out0 && v$Z2_4345_out0;
assign v$G10_11273_out0 = ! v$Z3_12567_out0;
assign v$G10_11274_out0 = ! v$Z3_12571_out0;
assign v$G10_11275_out0 = ! v$Z3_12575_out0;
assign v$G10_11276_out0 = ! v$Z3_12579_out0;
assign v$_3461_out0 = { v$OUT_6201_out0,v$C5_11957_out0 };
assign v$_3465_out0 = { v$OUT_6205_out0,v$C5_11961_out0 };
assign v$_3469_out0 = { v$OUT_6209_out0,v$C5_11965_out0 };
assign v$_3473_out0 = { v$OUT_6213_out0,v$C5_11969_out0 };
assign v$_6021_out0 = { v$OUT_6200_out0,v$C6_4536_out0 };
assign v$_6025_out0 = { v$OUT_6204_out0,v$C6_4540_out0 };
assign v$_6029_out0 = { v$OUT_6208_out0,v$C6_4544_out0 };
assign v$_6033_out0 = { v$OUT_6212_out0,v$C6_4548_out0 };
assign v$_6147_out0 = { v$OUT_6202_out0,v$C4_11588_out0 };
assign v$_6151_out0 = { v$OUT_6206_out0,v$C4_11592_out0 };
assign v$_6155_out0 = { v$OUT_6210_out0,v$C4_11596_out0 };
assign v$_6159_out0 = { v$OUT_6214_out0,v$C4_11600_out0 };
assign v$G7_6593_out0 = v$G9_10503_out0 && v$Z3_12567_out0;
assign v$G7_6597_out0 = v$G9_10507_out0 && v$Z3_12571_out0;
assign v$G7_6601_out0 = v$G9_10511_out0 && v$Z3_12575_out0;
assign v$G7_6605_out0 = v$G9_10515_out0 && v$Z3_12579_out0;
assign v$MUX12_12609_out0 = v$EQ12_9356_out0 ? v$SEL12_9362_out0 : v$MUX13_9228_out0;
assign v$MUX12_12610_out0 = v$EQ12_9357_out0 ? v$SEL12_9363_out0 : v$MUX13_9229_out0;
assign v$MUX12_12611_out0 = v$EQ12_9358_out0 ? v$SEL12_9364_out0 : v$MUX13_9230_out0;
assign v$MUX12_12612_out0 = v$EQ12_9359_out0 ? v$SEL12_9365_out0 : v$MUX13_9231_out0;
assign v$Z_1460_out0 = v$G7_6593_out0;
assign v$Z_1464_out0 = v$G7_6597_out0;
assign v$Z_1468_out0 = v$G7_6601_out0;
assign v$Z_1472_out0 = v$G7_6605_out0;
assign v$MUX5_2764_out0 = v$G6_4183_out0 ? v$_3461_out0 : v$_6021_out0;
assign v$MUX5_2768_out0 = v$G6_4187_out0 ? v$_3465_out0 : v$_6025_out0;
assign v$MUX5_2772_out0 = v$G6_4191_out0 ? v$_3469_out0 : v$_6029_out0;
assign v$MUX5_2776_out0 = v$G6_4195_out0 ? v$_3473_out0 : v$_6033_out0;
assign v$MUX11_12709_out0 = v$EQ11_4157_out0 ? v$SEL11_4834_out0 : v$MUX12_12609_out0;
assign v$MUX11_12710_out0 = v$EQ11_4158_out0 ? v$SEL11_4835_out0 : v$MUX12_12610_out0;
assign v$MUX11_12711_out0 = v$EQ11_4159_out0 ? v$SEL11_4836_out0 : v$MUX12_12611_out0;
assign v$MUX11_12712_out0 = v$EQ11_4160_out0 ? v$SEL11_4837_out0 : v$MUX12_12612_out0;
assign v$MUX4_1641_out0 = v$G10_11273_out0 ? v$_6147_out0 : v$MUX5_2764_out0;
assign v$MUX4_1645_out0 = v$G10_11274_out0 ? v$_6151_out0 : v$MUX5_2768_out0;
assign v$MUX4_1649_out0 = v$G10_11275_out0 ? v$_6155_out0 : v$MUX5_2772_out0;
assign v$MUX4_1653_out0 = v$G10_11276_out0 ? v$_6159_out0 : v$MUX5_2776_out0;
assign v$MUX8_1711_out0 = v$EQ9_9300_out0 ? v$SEL9_6829_out0 : v$MUX11_12709_out0;
assign v$MUX8_1712_out0 = v$EQ9_9301_out0 ? v$SEL9_6830_out0 : v$MUX11_12710_out0;
assign v$MUX8_1713_out0 = v$EQ9_9302_out0 ? v$SEL9_6831_out0 : v$MUX11_12711_out0;
assign v$MUX8_1714_out0 = v$EQ9_9303_out0 ? v$SEL9_6832_out0 : v$MUX11_12712_out0;
assign v$Z_11031_out0 = v$Z_1460_out0;
assign v$Z_11032_out0 = v$Z_1464_out0;
assign v$Z_11033_out0 = v$Z_1468_out0;
assign v$Z_11034_out0 = v$Z_1472_out0;
assign v$OUT_6199_out0 = v$MUX4_1641_out0;
assign v$OUT_6203_out0 = v$MUX4_1645_out0;
assign v$OUT_6207_out0 = v$MUX4_1649_out0;
assign v$OUT_6211_out0 = v$MUX4_1653_out0;
assign v$MUX10_10936_out0 = v$EQ10_3914_out0 ? v$SEL8_12507_out0 : v$MUX8_1711_out0;
assign v$MUX10_10937_out0 = v$EQ10_3915_out0 ? v$SEL8_12508_out0 : v$MUX8_1712_out0;
assign v$MUX10_10938_out0 = v$EQ10_3916_out0 ? v$SEL8_12509_out0 : v$MUX8_1713_out0;
assign v$MUX10_10939_out0 = v$EQ10_3917_out0 ? v$SEL8_12510_out0 : v$MUX8_1714_out0;
assign v$MUX9_5726_out0 = v$EQ8_9797_out0 ? v$SEL10_6487_out0 : v$MUX10_10936_out0;
assign v$MUX9_5727_out0 = v$EQ8_9798_out0 ? v$SEL10_6488_out0 : v$MUX10_10937_out0;
assign v$MUX9_5728_out0 = v$EQ8_9799_out0 ? v$SEL10_6489_out0 : v$MUX10_10938_out0;
assign v$MUX9_5729_out0 = v$EQ8_9800_out0 ? v$SEL10_6490_out0 : v$MUX10_10939_out0;
assign v$AMOUNT$OF$SHIFT_6455_out0 = v$OUT_6199_out0;
assign v$AMOUNT$OF$SHIFT_6456_out0 = v$OUT_6203_out0;
assign v$AMOUNT$OF$SHIFT_6457_out0 = v$OUT_6207_out0;
assign v$AMOUNT$OF$SHIFT_6458_out0 = v$OUT_6211_out0;
assign v$MUX7_496_out0 = v$EQ7_2788_out0 ? v$SEL7_9719_out0 : v$MUX9_5726_out0;
assign v$MUX7_497_out0 = v$EQ7_2789_out0 ? v$SEL7_9720_out0 : v$MUX9_5727_out0;
assign v$MUX7_498_out0 = v$EQ7_2790_out0 ? v$SEL7_9721_out0 : v$MUX9_5728_out0;
assign v$MUX7_499_out0 = v$EQ7_2791_out0 ? v$SEL7_9722_out0 : v$MUX9_5729_out0;
assign v$SEL4_1017_out0 = v$AMOUNT$OF$SHIFT_6455_out0[3:3];
assign v$SEL4_1018_out0 = v$AMOUNT$OF$SHIFT_6456_out0[3:3];
assign v$SEL4_1019_out0 = v$AMOUNT$OF$SHIFT_6457_out0[3:3];
assign v$SEL4_1020_out0 = v$AMOUNT$OF$SHIFT_6458_out0[3:3];
assign v$SEL6_6178_out0 = v$AMOUNT$OF$SHIFT_6455_out0[5:5];
assign v$SEL6_6179_out0 = v$AMOUNT$OF$SHIFT_6456_out0[5:5];
assign v$SEL6_6180_out0 = v$AMOUNT$OF$SHIFT_6457_out0[5:5];
assign v$SEL6_6181_out0 = v$AMOUNT$OF$SHIFT_6458_out0[5:5];
assign v$SEL5_7496_out0 = v$AMOUNT$OF$SHIFT_6455_out0[4:4];
assign v$SEL5_7497_out0 = v$AMOUNT$OF$SHIFT_6456_out0[4:4];
assign v$SEL5_7498_out0 = v$AMOUNT$OF$SHIFT_6457_out0[4:4];
assign v$SEL5_7499_out0 = v$AMOUNT$OF$SHIFT_6458_out0[4:4];
assign v$SEL1_8929_out0 = v$AMOUNT$OF$SHIFT_6455_out0[0:0];
assign v$SEL1_8930_out0 = v$AMOUNT$OF$SHIFT_6456_out0[0:0];
assign v$SEL1_8931_out0 = v$AMOUNT$OF$SHIFT_6457_out0[0:0];
assign v$SEL1_8932_out0 = v$AMOUNT$OF$SHIFT_6458_out0[0:0];
assign v$SEL3_9405_out0 = v$AMOUNT$OF$SHIFT_6455_out0[2:2];
assign v$SEL3_9406_out0 = v$AMOUNT$OF$SHIFT_6456_out0[2:2];
assign v$SEL3_9407_out0 = v$AMOUNT$OF$SHIFT_6457_out0[2:2];
assign v$SEL3_9408_out0 = v$AMOUNT$OF$SHIFT_6458_out0[2:2];
assign v$SEL2_13163_out0 = v$AMOUNT$OF$SHIFT_6455_out0[1:1];
assign v$SEL2_13164_out0 = v$AMOUNT$OF$SHIFT_6456_out0[1:1];
assign v$SEL2_13165_out0 = v$AMOUNT$OF$SHIFT_6457_out0[1:1];
assign v$SEL2_13166_out0 = v$AMOUNT$OF$SHIFT_6458_out0[1:1];
assign v$EN_563_out0 = v$SEL4_1017_out0;
assign v$EN_564_out0 = v$SEL4_1018_out0;
assign v$EN_573_out0 = v$SEL4_1019_out0;
assign v$EN_574_out0 = v$SEL4_1020_out0;
assign v$EN_3166_out0 = v$SEL3_9405_out0;
assign v$EN_3167_out0 = v$SEL3_9406_out0;
assign v$EN_3172_out0 = v$SEL3_9407_out0;
assign v$EN_3173_out0 = v$SEL3_9408_out0;
assign v$EN_3586_out0 = v$SEL6_6178_out0;
assign v$EN_3587_out0 = v$SEL5_7496_out0;
assign v$EN_3588_out0 = v$SEL1_8929_out0;
assign v$EN_3589_out0 = v$SEL6_6179_out0;
assign v$EN_3590_out0 = v$SEL5_7497_out0;
assign v$EN_3591_out0 = v$SEL1_8930_out0;
assign v$EN_3596_out0 = v$SEL6_6180_out0;
assign v$EN_3597_out0 = v$SEL5_7498_out0;
assign v$EN_3598_out0 = v$SEL1_8931_out0;
assign v$EN_3599_out0 = v$SEL6_6181_out0;
assign v$EN_3600_out0 = v$SEL5_7499_out0;
assign v$EN_3601_out0 = v$SEL1_8932_out0;
assign v$EN_5390_out0 = v$SEL2_13163_out0;
assign v$EN_5391_out0 = v$SEL2_13164_out0;
assign v$EN_5396_out0 = v$SEL2_13165_out0;
assign v$EN_5397_out0 = v$SEL2_13166_out0;
assign v$MUX6_11420_out0 = v$EQ6_3671_out0 ? v$SEL6_8113_out0 : v$MUX7_496_out0;
assign v$MUX6_11421_out0 = v$EQ6_3672_out0 ? v$SEL6_8114_out0 : v$MUX7_497_out0;
assign v$MUX6_11422_out0 = v$EQ6_3673_out0 ? v$SEL6_8115_out0 : v$MUX7_498_out0;
assign v$MUX6_11423_out0 = v$EQ6_3674_out0 ? v$SEL6_8116_out0 : v$MUX7_499_out0;
assign v$MUX5_4698_out0 = v$EQ5_2013_out0 ? v$SEL5_10744_out0 : v$MUX6_11420_out0;
assign v$MUX5_4699_out0 = v$EQ5_2014_out0 ? v$SEL5_10745_out0 : v$MUX6_11421_out0;
assign v$MUX5_4700_out0 = v$EQ5_2015_out0 ? v$SEL5_10746_out0 : v$MUX6_11422_out0;
assign v$MUX5_4701_out0 = v$EQ5_2016_out0 ? v$SEL5_10747_out0 : v$MUX6_11423_out0;
assign v$MUX2_13220_out0 = v$EN_3588_out0 ? v$MUX1_1292_out0 : v$IN_2569_out0;
assign v$MUX2_13223_out0 = v$EN_3591_out0 ? v$MUX1_1298_out0 : v$IN_2572_out0;
assign v$MUX2_13230_out0 = v$EN_3598_out0 ? v$MUX1_1324_out0 : v$IN_2579_out0;
assign v$MUX2_13233_out0 = v$EN_3601_out0 ? v$MUX1_1330_out0 : v$IN_2582_out0;
assign v$MUX4_5324_out0 = v$EQ4_13241_out0 ? v$SEL4_4919_out0 : v$MUX5_4698_out0;
assign v$MUX4_5325_out0 = v$EQ4_13242_out0 ? v$SEL4_4920_out0 : v$MUX5_4699_out0;
assign v$MUX4_5326_out0 = v$EQ4_13243_out0 ? v$SEL4_4921_out0 : v$MUX5_4700_out0;
assign v$MUX4_5327_out0 = v$EQ4_13244_out0 ? v$SEL4_4922_out0 : v$MUX5_4701_out0;
assign v$OUT_10243_out0 = v$MUX2_13220_out0;
assign v$OUT_10249_out0 = v$MUX2_13223_out0;
assign v$OUT_10275_out0 = v$MUX2_13230_out0;
assign v$OUT_10281_out0 = v$MUX2_13233_out0;
assign v$IN_3528_out0 = v$OUT_10243_out0;
assign v$IN_3534_out0 = v$OUT_10249_out0;
assign v$IN_3560_out0 = v$OUT_10275_out0;
assign v$IN_3566_out0 = v$OUT_10281_out0;
assign v$MUX3_5138_out0 = v$EQ3_991_out0 ? v$SEL3_7544_out0 : v$MUX4_5324_out0;
assign v$MUX3_5139_out0 = v$EQ3_992_out0 ? v$SEL3_7545_out0 : v$MUX4_5325_out0;
assign v$MUX3_5140_out0 = v$EQ3_993_out0 ? v$SEL3_7546_out0 : v$MUX4_5326_out0;
assign v$MUX3_5141_out0 = v$EQ3_994_out0 ? v$SEL3_7547_out0 : v$MUX4_5327_out0;
assign v$IN_7583_out0 = v$IN_3528_out0;
assign v$IN_7584_out0 = v$IN_3534_out0;
assign v$IN_7589_out0 = v$IN_3560_out0;
assign v$IN_7590_out0 = v$IN_3566_out0;
assign v$MUX2_9170_out0 = v$EQ2_9605_out0 ? v$SEL2_8895_out0 : v$MUX3_5138_out0;
assign v$MUX2_9171_out0 = v$EQ2_9606_out0 ? v$SEL2_8896_out0 : v$MUX3_5139_out0;
assign v$MUX2_9172_out0 = v$EQ2_9607_out0 ? v$SEL2_8897_out0 : v$MUX3_5140_out0;
assign v$MUX2_9173_out0 = v$EQ2_9608_out0 ? v$SEL2_8898_out0 : v$MUX3_5141_out0;
assign v$MUX1_1635_out0 = v$EQ1_8984_out0 ? v$SEL1_4817_out0 : v$MUX2_9170_out0;
assign v$MUX1_1636_out0 = v$EQ1_8985_out0 ? v$SEL1_4818_out0 : v$MUX2_9171_out0;
assign v$MUX1_1637_out0 = v$EQ1_8986_out0 ? v$SEL1_4819_out0 : v$MUX2_9172_out0;
assign v$MUX1_1638_out0 = v$EQ1_8987_out0 ? v$SEL1_4820_out0 : v$MUX2_9173_out0;
assign v$SEL1_5941_out0 = v$IN_7583_out0[47:2];
assign v$SEL1_5947_out0 = v$IN_7584_out0[47:2];
assign v$SEL1_5973_out0 = v$IN_7589_out0[47:2];
assign v$SEL1_5979_out0 = v$IN_7590_out0[47:2];
assign v$SEL1_10685_out0 = v$IN_7583_out0[45:0];
assign v$SEL1_10691_out0 = v$IN_7584_out0[45:0];
assign v$SEL1_10717_out0 = v$IN_7589_out0[45:0];
assign v$SEL1_10723_out0 = v$IN_7590_out0[45:0];
assign v$_2927_out0 = { v$C2_103_out0,v$SEL1_10685_out0 };
assign v$_2933_out0 = { v$C2_109_out0,v$SEL1_10691_out0 };
assign v$_2959_out0 = { v$C2_135_out0,v$SEL1_10717_out0 };
assign v$_2965_out0 = { v$C2_141_out0,v$SEL1_10723_out0 };
assign v$MUX25_5870_out0 = v$G2_7692_out0 ? v$C2_10483_out0 : v$MUX1_1635_out0;
assign v$MUX25_5871_out0 = v$G2_7693_out0 ? v$C2_10484_out0 : v$MUX1_1636_out0;
assign v$MUX25_5872_out0 = v$G2_7694_out0 ? v$C2_10485_out0 : v$MUX1_1637_out0;
assign v$MUX25_5873_out0 = v$G2_7695_out0 ? v$C2_10486_out0 : v$MUX1_1638_out0;
assign v$_6234_out0 = { v$SEL1_5941_out0,v$C1_3970_out0 };
assign v$_6240_out0 = { v$SEL1_5947_out0,v$C1_3976_out0 };
assign v$_6266_out0 = { v$SEL1_5973_out0,v$C1_4002_out0 };
assign v$_6272_out0 = { v$SEL1_5979_out0,v$C1_4008_out0 };
assign v$MUX1_1290_out0 = v$LEFT$SHIT_1802_out0 ? v$_2927_out0 : v$_6234_out0;
assign v$MUX1_1296_out0 = v$LEFT$SHIT_1808_out0 ? v$_2933_out0 : v$_6240_out0;
assign v$MUX1_1322_out0 = v$LEFT$SHIT_1834_out0 ? v$_2959_out0 : v$_6266_out0;
assign v$MUX1_1328_out0 = v$LEFT$SHIT_1840_out0 ? v$_2965_out0 : v$_6272_out0;
assign v$OUT_6467_out0 = v$MUX25_5870_out0;
assign v$OUT_6468_out0 = v$MUX25_5871_out0;
assign v$OUT_6469_out0 = v$MUX25_5872_out0;
assign v$OUT_6470_out0 = v$MUX25_5873_out0;
assign v$MUX2_1394_out0 = v$EN_5390_out0 ? v$MUX1_1290_out0 : v$IN_7583_out0;
assign v$MUX2_1395_out0 = v$EN_5391_out0 ? v$MUX1_1296_out0 : v$IN_7584_out0;
assign v$MUX2_1400_out0 = v$EN_5396_out0 ? v$MUX1_1322_out0 : v$IN_7589_out0;
assign v$MUX2_1401_out0 = v$EN_5397_out0 ? v$MUX1_1328_out0 : v$IN_7590_out0;
assign {v$A1_1564_out1,v$A1_1564_out0 } = v$LARGER$EXP_6839_out0 + v$SMALLER$EXP_1707_out0 + v$OUT_6467_out0;
assign {v$A1_1565_out1,v$A1_1565_out0 } = v$LARGER$EXP_6840_out0 + v$SMALLER$EXP_1708_out0 + v$OUT_6468_out0;
assign {v$A1_1566_out1,v$A1_1566_out0 } = v$LARGER$EXP_6841_out0 + v$SMALLER$EXP_1709_out0 + v$OUT_6469_out0;
assign {v$A1_1567_out1,v$A1_1567_out0 } = v$LARGER$EXP_6842_out0 + v$SMALLER$EXP_1710_out0 + v$OUT_6470_out0;
assign {v$A2_6750_out1,v$A2_6750_out0 } = v$A1_1564_out0 + v$C1_3957_out0 + v$C2_11416_out0;
assign {v$A2_6751_out1,v$A2_6751_out0 } = v$A1_1565_out0 + v$C1_3958_out0 + v$C2_11417_out0;
assign {v$A2_6752_out1,v$A2_6752_out0 } = v$A1_1566_out0 + v$C1_3959_out0 + v$C2_11418_out0;
assign {v$A2_6753_out1,v$A2_6753_out0 } = v$A1_1567_out0 + v$C1_3960_out0 + v$C2_11419_out0;
assign v$OUT_10241_out0 = v$MUX2_1394_out0;
assign v$OUT_10247_out0 = v$MUX2_1395_out0;
assign v$OUT_10273_out0 = v$MUX2_1400_out0;
assign v$OUT_10279_out0 = v$MUX2_1401_out0;
assign v$NOT$USED$CARRY_13402_out0 = v$A1_1564_out1;
assign v$NOT$USED$CARRY_13403_out0 = v$A1_1565_out1;
assign v$NOT$USED$CARRY_13404_out0 = v$A1_1566_out1;
assign v$NOT$USED$CARRY_13405_out0 = v$A1_1567_out1;
assign v$IN_3531_out0 = v$OUT_10241_out0;
assign v$IN_3537_out0 = v$OUT_10247_out0;
assign v$IN_3563_out0 = v$OUT_10273_out0;
assign v$IN_3569_out0 = v$OUT_10279_out0;
assign v$NOT$USED_11148_out0 = v$A2_6750_out1;
assign v$NOT$USED_11149_out0 = v$A2_6751_out1;
assign v$NOT$USED_11150_out0 = v$A2_6752_out1;
assign v$NOT$USED_11151_out0 = v$A2_6753_out1;
assign v$IN_10873_out0 = v$IN_3531_out0;
assign v$IN_10874_out0 = v$IN_3537_out0;
assign v$IN_10879_out0 = v$IN_3563_out0;
assign v$IN_10880_out0 = v$IN_3569_out0;
assign v$SEL1_5944_out0 = v$IN_10873_out0[47:4];
assign v$SEL1_5950_out0 = v$IN_10874_out0[47:4];
assign v$SEL1_5976_out0 = v$IN_10879_out0[47:4];
assign v$SEL1_5982_out0 = v$IN_10880_out0[47:4];
assign v$SEL1_10688_out0 = v$IN_10873_out0[43:0];
assign v$SEL1_10694_out0 = v$IN_10874_out0[43:0];
assign v$SEL1_10720_out0 = v$IN_10879_out0[43:0];
assign v$SEL1_10726_out0 = v$IN_10880_out0[43:0];
assign v$_2930_out0 = { v$C2_106_out0,v$SEL1_10688_out0 };
assign v$_2936_out0 = { v$C2_112_out0,v$SEL1_10694_out0 };
assign v$_2962_out0 = { v$C2_138_out0,v$SEL1_10720_out0 };
assign v$_2968_out0 = { v$C2_144_out0,v$SEL1_10726_out0 };
assign v$_6237_out0 = { v$SEL1_5944_out0,v$C1_3973_out0 };
assign v$_6243_out0 = { v$SEL1_5950_out0,v$C1_3979_out0 };
assign v$_6269_out0 = { v$SEL1_5976_out0,v$C1_4005_out0 };
assign v$_6275_out0 = { v$SEL1_5982_out0,v$C1_4011_out0 };
assign v$MUX1_1293_out0 = v$LEFT$SHIT_1805_out0 ? v$_2930_out0 : v$_6237_out0;
assign v$MUX1_1299_out0 = v$LEFT$SHIT_1811_out0 ? v$_2936_out0 : v$_6243_out0;
assign v$MUX1_1325_out0 = v$LEFT$SHIT_1837_out0 ? v$_2962_out0 : v$_6269_out0;
assign v$MUX1_1331_out0 = v$LEFT$SHIT_1843_out0 ? v$_2968_out0 : v$_6275_out0;
assign v$MUX2_10556_out0 = v$EN_3166_out0 ? v$MUX1_1293_out0 : v$IN_10873_out0;
assign v$MUX2_10557_out0 = v$EN_3167_out0 ? v$MUX1_1299_out0 : v$IN_10874_out0;
assign v$MUX2_10562_out0 = v$EN_3172_out0 ? v$MUX1_1325_out0 : v$IN_10879_out0;
assign v$MUX2_10563_out0 = v$EN_3173_out0 ? v$MUX1_1331_out0 : v$IN_10880_out0;
assign v$OUT_10244_out0 = v$MUX2_10556_out0;
assign v$OUT_10250_out0 = v$MUX2_10557_out0;
assign v$OUT_10276_out0 = v$MUX2_10562_out0;
assign v$OUT_10282_out0 = v$MUX2_10563_out0;
assign v$IN_3527_out0 = v$OUT_10244_out0;
assign v$IN_3533_out0 = v$OUT_10250_out0;
assign v$IN_3559_out0 = v$OUT_10276_out0;
assign v$IN_3565_out0 = v$OUT_10282_out0;
assign v$IN_3413_out0 = v$IN_3527_out0;
assign v$IN_3414_out0 = v$IN_3533_out0;
assign v$IN_3423_out0 = v$IN_3559_out0;
assign v$IN_3424_out0 = v$IN_3565_out0;
assign v$SEL1_5940_out0 = v$IN_3413_out0[47:8];
assign v$SEL1_5946_out0 = v$IN_3414_out0[47:8];
assign v$SEL1_5972_out0 = v$IN_3423_out0[47:8];
assign v$SEL1_5978_out0 = v$IN_3424_out0[47:8];
assign v$SEL1_10684_out0 = v$IN_3413_out0[39:0];
assign v$SEL1_10690_out0 = v$IN_3414_out0[39:0];
assign v$SEL1_10716_out0 = v$IN_3423_out0[39:0];
assign v$SEL1_10722_out0 = v$IN_3424_out0[39:0];
assign v$_2926_out0 = { v$C2_102_out0,v$SEL1_10684_out0 };
assign v$_2932_out0 = { v$C2_108_out0,v$SEL1_10690_out0 };
assign v$_2958_out0 = { v$C2_134_out0,v$SEL1_10716_out0 };
assign v$_2964_out0 = { v$C2_140_out0,v$SEL1_10722_out0 };
assign v$_6233_out0 = { v$SEL1_5940_out0,v$C1_3969_out0 };
assign v$_6239_out0 = { v$SEL1_5946_out0,v$C1_3975_out0 };
assign v$_6265_out0 = { v$SEL1_5972_out0,v$C1_4001_out0 };
assign v$_6271_out0 = { v$SEL1_5978_out0,v$C1_4007_out0 };
assign v$MUX1_1289_out0 = v$LEFT$SHIT_1801_out0 ? v$_2926_out0 : v$_6233_out0;
assign v$MUX1_1295_out0 = v$LEFT$SHIT_1807_out0 ? v$_2932_out0 : v$_6239_out0;
assign v$MUX1_1321_out0 = v$LEFT$SHIT_1833_out0 ? v$_2958_out0 : v$_6265_out0;
assign v$MUX1_1327_out0 = v$LEFT$SHIT_1839_out0 ? v$_2964_out0 : v$_6271_out0;
assign v$MUX2_1407_out0 = v$EN_563_out0 ? v$MUX1_1289_out0 : v$IN_3413_out0;
assign v$MUX2_1408_out0 = v$EN_564_out0 ? v$MUX1_1295_out0 : v$IN_3414_out0;
assign v$MUX2_1417_out0 = v$EN_573_out0 ? v$MUX1_1321_out0 : v$IN_3423_out0;
assign v$MUX2_1418_out0 = v$EN_574_out0 ? v$MUX1_1327_out0 : v$IN_3424_out0;
assign v$OUT_10240_out0 = v$MUX2_1407_out0;
assign v$OUT_10246_out0 = v$MUX2_1408_out0;
assign v$OUT_10272_out0 = v$MUX2_1417_out0;
assign v$OUT_10278_out0 = v$MUX2_1418_out0;
assign v$IN_3529_out0 = v$OUT_10240_out0;
assign v$IN_3535_out0 = v$OUT_10246_out0;
assign v$IN_3561_out0 = v$OUT_10272_out0;
assign v$IN_3567_out0 = v$OUT_10278_out0;
assign v$IN_2568_out0 = v$IN_3529_out0;
assign v$IN_2571_out0 = v$IN_3535_out0;
assign v$IN_2578_out0 = v$IN_3561_out0;
assign v$IN_2581_out0 = v$IN_3567_out0;
assign v$SEL1_5942_out0 = v$IN_2568_out0[47:16];
assign v$SEL1_5948_out0 = v$IN_2571_out0[47:16];
assign v$SEL1_5974_out0 = v$IN_2578_out0[47:16];
assign v$SEL1_5980_out0 = v$IN_2581_out0[47:16];
assign v$SEL1_10686_out0 = v$IN_2568_out0[31:0];
assign v$SEL1_10692_out0 = v$IN_2571_out0[31:0];
assign v$SEL1_10718_out0 = v$IN_2578_out0[31:0];
assign v$SEL1_10724_out0 = v$IN_2581_out0[31:0];
assign v$_2928_out0 = { v$C2_104_out0,v$SEL1_10686_out0 };
assign v$_2934_out0 = { v$C2_110_out0,v$SEL1_10692_out0 };
assign v$_2960_out0 = { v$C2_136_out0,v$SEL1_10718_out0 };
assign v$_2966_out0 = { v$C2_142_out0,v$SEL1_10724_out0 };
assign v$_6235_out0 = { v$SEL1_5942_out0,v$C1_3971_out0 };
assign v$_6241_out0 = { v$SEL1_5948_out0,v$C1_3977_out0 };
assign v$_6267_out0 = { v$SEL1_5974_out0,v$C1_4003_out0 };
assign v$_6273_out0 = { v$SEL1_5980_out0,v$C1_4009_out0 };
assign v$MUX1_1291_out0 = v$LEFT$SHIT_1803_out0 ? v$_2928_out0 : v$_6235_out0;
assign v$MUX1_1297_out0 = v$LEFT$SHIT_1809_out0 ? v$_2934_out0 : v$_6241_out0;
assign v$MUX1_1323_out0 = v$LEFT$SHIT_1835_out0 ? v$_2960_out0 : v$_6267_out0;
assign v$MUX1_1329_out0 = v$LEFT$SHIT_1841_out0 ? v$_2966_out0 : v$_6273_out0;
assign v$MUX2_13219_out0 = v$EN_3587_out0 ? v$MUX1_1291_out0 : v$IN_2568_out0;
assign v$MUX2_13222_out0 = v$EN_3590_out0 ? v$MUX1_1297_out0 : v$IN_2571_out0;
assign v$MUX2_13229_out0 = v$EN_3597_out0 ? v$MUX1_1323_out0 : v$IN_2578_out0;
assign v$MUX2_13232_out0 = v$EN_3600_out0 ? v$MUX1_1329_out0 : v$IN_2581_out0;
assign v$OUT_10242_out0 = v$MUX2_13219_out0;
assign v$OUT_10248_out0 = v$MUX2_13222_out0;
assign v$OUT_10274_out0 = v$MUX2_13229_out0;
assign v$OUT_10280_out0 = v$MUX2_13232_out0;
assign v$IN_3526_out0 = v$OUT_10242_out0;
assign v$IN_3532_out0 = v$OUT_10248_out0;
assign v$IN_3558_out0 = v$OUT_10274_out0;
assign v$IN_3564_out0 = v$OUT_10280_out0;
assign v$IN_2567_out0 = v$IN_3526_out0;
assign v$IN_2570_out0 = v$IN_3532_out0;
assign v$IN_2577_out0 = v$IN_3558_out0;
assign v$IN_2580_out0 = v$IN_3564_out0;
assign v$SEL1_5939_out0 = v$IN_2567_out0[47:32];
assign v$SEL1_5945_out0 = v$IN_2570_out0[47:32];
assign v$SEL1_5971_out0 = v$IN_2577_out0[47:32];
assign v$SEL1_5977_out0 = v$IN_2580_out0[47:32];
assign v$SEL1_10683_out0 = v$IN_2567_out0[15:0];
assign v$SEL1_10689_out0 = v$IN_2570_out0[15:0];
assign v$SEL1_10715_out0 = v$IN_2577_out0[15:0];
assign v$SEL1_10721_out0 = v$IN_2580_out0[15:0];
assign v$_2925_out0 = { v$C2_101_out0,v$SEL1_10683_out0 };
assign v$_2931_out0 = { v$C2_107_out0,v$SEL1_10689_out0 };
assign v$_2957_out0 = { v$C2_133_out0,v$SEL1_10715_out0 };
assign v$_2963_out0 = { v$C2_139_out0,v$SEL1_10721_out0 };
assign v$_6232_out0 = { v$SEL1_5939_out0,v$C1_3968_out0 };
assign v$_6238_out0 = { v$SEL1_5945_out0,v$C1_3974_out0 };
assign v$_6264_out0 = { v$SEL1_5971_out0,v$C1_4000_out0 };
assign v$_6270_out0 = { v$SEL1_5977_out0,v$C1_4006_out0 };
assign v$MUX1_1288_out0 = v$LEFT$SHIT_1800_out0 ? v$_2925_out0 : v$_6232_out0;
assign v$MUX1_1294_out0 = v$LEFT$SHIT_1806_out0 ? v$_2931_out0 : v$_6238_out0;
assign v$MUX1_1320_out0 = v$LEFT$SHIT_1832_out0 ? v$_2957_out0 : v$_6264_out0;
assign v$MUX1_1326_out0 = v$LEFT$SHIT_1838_out0 ? v$_2963_out0 : v$_6270_out0;
assign v$MUX2_13218_out0 = v$EN_3586_out0 ? v$MUX1_1288_out0 : v$IN_2567_out0;
assign v$MUX2_13221_out0 = v$EN_3589_out0 ? v$MUX1_1294_out0 : v$IN_2570_out0;
assign v$MUX2_13228_out0 = v$EN_3596_out0 ? v$MUX1_1320_out0 : v$IN_2577_out0;
assign v$MUX2_13231_out0 = v$EN_3599_out0 ? v$MUX1_1326_out0 : v$IN_2580_out0;
assign v$OUT_10239_out0 = v$MUX2_13218_out0;
assign v$OUT_10245_out0 = v$MUX2_13221_out0;
assign v$OUT_10271_out0 = v$MUX2_13228_out0;
assign v$OUT_10277_out0 = v$MUX2_13231_out0;
assign v$OUT_3306_out0 = v$OUT_10239_out0;
assign v$OUT_3307_out0 = v$OUT_10245_out0;
assign v$OUT_3308_out0 = v$OUT_10271_out0;
assign v$OUT_3309_out0 = v$OUT_10277_out0;
assign v$SEL2_5605_out0 = v$OUT_3306_out0[46:37];
assign v$SEL2_5606_out0 = v$OUT_3307_out0[46:24];
assign v$SEL2_5607_out0 = v$OUT_3308_out0[46:37];
assign v$SEL2_5608_out0 = v$OUT_3309_out0[46:24];
assign v$_11064_out0 = { v$SEL2_5605_out0,v$A2_6750_out0 };
assign v$_11065_out0 = { v$SEL2_5606_out0,v$A2_6751_out0 };
assign v$_11066_out0 = { v$SEL2_5607_out0,v$A2_6752_out0 };
assign v$_11067_out0 = { v$SEL2_5608_out0,v$A2_6753_out0 };
assign v$MUX2_9187_out0 = v$Z_11031_out0 ? v$C4_5739_out0 : v$_11064_out0;
assign v$MUX2_9188_out0 = v$Z_11032_out0 ? v$C4_5740_out0 : v$_11065_out0;
assign v$MUX2_9189_out0 = v$Z_11033_out0 ? v$C4_5741_out0 : v$_11066_out0;
assign v$MUX2_9190_out0 = v$Z_11034_out0 ? v$C4_5742_out0 : v$_11067_out0;
assign v$_13103_out0 = { v$MUX2_9187_out0,v$SIGN_591_out0 };
assign v$_13104_out0 = { v$MUX2_9188_out0,v$SIGN_592_out0 };
assign v$_13105_out0 = { v$MUX2_9189_out0,v$SIGN_593_out0 };
assign v$_13106_out0 = { v$MUX2_9190_out0,v$SIGN_594_out0 };
assign v$OUT_8119_out0 = v$_13103_out0;
assign v$OUT_8120_out0 = v$_13104_out0;
assign v$OUT_8121_out0 = v$_13105_out0;
assign v$OUT_8122_out0 = v$_13106_out0;
assign v$MUX11_5920_out0 = v$G5_4215_out0 ? v$C9_13387_out0 : v$OUT_8119_out0;
assign v$MUX11_5921_out0 = v$G5_4216_out0 ? v$C9_13388_out0 : v$OUT_8121_out0;
assign v$MUX3_6217_out0 = v$G3_11192_out0 ? v$C1_10547_out0 : v$OUT_8120_out0;
assign v$MUX3_6218_out0 = v$G3_11193_out0 ? v$C1_10548_out0 : v$OUT_8122_out0;
assign v$SINGLE$PRECISION_5416_out0 = v$MUX3_6217_out0;
assign v$SINGLE$PRECISION_5417_out0 = v$MUX3_6218_out0;
assign v$_12090_out0 = { v$C10_4403_out0,v$MUX11_5920_out0 };
assign v$_12091_out0 = { v$C10_4404_out0,v$MUX11_5921_out0 };
assign v$HALF$PRECISION_6871_out0 = v$_12090_out0;
assign v$HALF$PRECISION_6872_out0 = v$_12091_out0;
assign v$MUX12_11834_out0 = v$IS$32$BITS_527_out0 ? v$SINGLE$PRECISION_5416_out0 : v$HALF$PRECISION_6871_out0;
assign v$MUX12_11835_out0 = v$IS$32$BITS_528_out0 ? v$SINGLE$PRECISION_5417_out0 : v$HALF$PRECISION_6872_out0;
assign v$OUT_2054_out0 = v$MUX12_11834_out0;
assign v$OUT_2055_out0 = v$MUX12_11835_out0;
assign v$MUX4_519_out0 = v$MUL_12088_out0 ? v$OUT_2054_out0 : v$MUX2_11385_out0;
assign v$MUX4_520_out0 = v$MUL_12089_out0 ? v$OUT_2055_out0 : v$MUX2_11386_out0;
assign v$SEL4_6522_out0 = v$MUX4_519_out0[15:0];
assign v$SEL4_6523_out0 = v$MUX4_520_out0[15:0];
assign v$SEL5_9159_out0 = v$MUX4_519_out0[31:16];
assign v$SEL5_9160_out0 = v$MUX4_520_out0[31:16];
assign v$MUX3_13078_out0 = v$G12_7750_out0 ? v$REG3_7578_out0 : v$SEL5_9159_out0;
assign v$MUX3_13079_out0 = v$G12_7751_out0 ? v$REG3_7579_out0 : v$SEL5_9160_out0;
assign v$OUT_551_out0 = v$MUX3_13078_out0;
assign v$OUT_552_out0 = v$MUX3_13079_out0;
assign v$FPU$OUT_12069_out0 = v$OUT_551_out0;
assign v$FPU$OUT_12070_out0 = v$OUT_552_out0;
assign v$MUX6_5016_out0 = v$G21_13310_out0 ? v$FPU$OUT_12069_out0 : v$MUX4_42_out0;
assign v$MUX6_5017_out0 = v$G21_13311_out0 ? v$FPU$OUT_12070_out0 : v$MUX4_43_out0;
assign v$DIN3_9801_out0 = v$MUX6_5016_out0;
assign v$DIN3_9802_out0 = v$MUX6_5017_out0;


endmodule

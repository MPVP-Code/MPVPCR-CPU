

    module v$RAM1_12913(q, a, d, we, clk);
    output reg [15:0] q;
    input [15:0] d;
    input [11:0] a;
    input we, clk;
    reg [15:0] ram [4095:0];
     always @(posedge clk) begin
         if (we)
             ram[a] <= d;
         q <= ram[a];
     end

    integer i;
    initial
    begin
        for (i=0; i < 4096; i=i+1)
        begin
            ram[i] = 0;
        end

        ram[0] = 4080;
ram[1] = 4059;
ram[2] = 16201;
ram[3] = 43691;
ram[4] = 15914;
ram[5] = 0;
ram[6] = 0;
ram[7] = 34953;
ram[8] = 15368;
ram[9] = 0;
ram[10] = 0;
ram[11] = 5120;
ram[12] = 14672;
ram[13] = 0;
ram[14] = 0;
ram[15] = 0;
ram[18] = 15944;
ram[19] = 12629;
ram[20] = 0;
ram[21] = 8260;
ram[22] = 0;
ram[23] = 5120;
ram[4080] = 14920;
ram[4081] = 12629;
ram[4082] = 0;
ram[4083] = 8260;
ram[4084] = 0;
ram[4085] = 0;
    end
    endmodule

    

    module v$AROM1_16158(q, a);
    output[43:0] q;
    input [5:0] a;
    reg [43:0] rom [63:0];

    assign q = rom[a];
    integer i;
    initial
    begin
        for (i=0; i < 64; i=i+1)
        begin
            rom[i] = 0;
        end
    
        rom[0] = 1030792151295;
rom[1] = 64424509695;
rom[2] = 1095216660735;
rom[3] = 4026532095;
rom[4] = 1034818683135;
rom[5] = 68451041535;
rom[6] = 1099243192575;
rom[7] = 251658495;
rom[8] = 1031043809535;
rom[9] = 64676167935;
rom[10] = 0;
    end
    endmodule
     

    module v$AROM1_16159(q, a);
    output[43:0] q;
    input [5:0] a;
    reg [43:0] rom [63:0];

    assign q = rom[a];
    integer i;
    initial
    begin
        for (i=0; i < 64; i=i+1)
        begin
            rom[i] = 0;
        end
    
        rom[0] = 1030792151295;
rom[1] = 64424509695;
rom[2] = 1095216660735;
rom[3] = 4026532095;
rom[4] = 1034818683135;
rom[5] = 68451041535;
rom[6] = 1099243192575;
rom[7] = 251658495;
rom[8] = 1031043809535;
rom[9] = 64676167935;
rom[10] = 0;
    end
    endmodule
     

    module v$ROM1_17450(q, a, clk);
    output reg [15:0] q;
    input clk;
    input [11:0] a;
    reg [15:0] rom [4095:0];
    always @(posedge clk) q <= rom[a];
    integer i;
    initial
    begin
        for (i=0; i < 4096; i=i+1)
        begin
            rom[i] = 0;
        end
    
        rom[0] = 3908;
rom[1] = 49668;
rom[2] = 95;
rom[3] = 1539;
rom[4] = 2631;
rom[5] = 49675;
rom[6] = 6657;
rom[7] = 107;
rom[8] = 28673;
rom[9] = 28672;
rom[10] = 28672;
rom[11] = 28677;
rom[12] = 6657;
rom[13] = 49682;
rom[14] = 107;
rom[15] = 28673;
rom[16] = 28672;
rom[17] = 28672;
rom[18] = 28677;
rom[19] = 6657;
rom[20] = 49689;
rom[21] = 107;
rom[22] = 28673;
rom[23] = 28672;
rom[24] = 28672;
rom[25] = 28677;
rom[26] = 5378;
rom[27] = 1035;
rom[28] = 1539;
rom[29] = 2639;
rom[30] = 6657;
rom[31] = 49683;
rom[32] = 49168;
rom[33] = 107;
rom[34] = 28673;
rom[35] = 28672;
rom[36] = 28672;
rom[37] = 0;
rom[38] = 28677;
rom[39] = 6657;
rom[40] = 49688;
rom[41] = 49168;
rom[42] = 107;
rom[43] = 28673;
rom[44] = 28672;
rom[45] = 28672;
rom[46] = 0;
rom[47] = 0;
rom[48] = 28677;
rom[49] = 6657;
rom[50] = 49692;
rom[51] = 49168;
rom[52] = 107;
rom[53] = 28673;
rom[54] = 28672;
rom[55] = 28672;
rom[56] = 28677;
rom[57] = 6657;
rom[58] = 49680;
rom[59] = 49184;
rom[60] = 107;
rom[61] = 28673;
rom[62] = 28672;
rom[63] = 28672;
rom[64] = 28677;
rom[65] = 6657;
rom[66] = 49683;
rom[67] = 49184;
rom[68] = 107;
rom[69] = 28673;
rom[70] = 28672;
rom[71] = 28672;
rom[72] = 0;
rom[73] = 0;
rom[74] = 0;
rom[75] = 0;
rom[76] = 28677;
rom[77] = 1547;
rom[78] = 6145;
rom[79] = 2055;
rom[80] = 28672;
rom[81] = 837;
rom[82] = 1537;
rom[83] = 5056;
rom[84] = 7040;
rom[85] = 5411;
rom[86] = 4864;
rom[87] = 52748;
rom[88] = 327;
rom[89] = 1027;
rom[90] = 28672;
    end
    endmodule
     

    module v$ROM1_17451(q, a, clk);
    output reg [15:0] q;
    input clk;
    input [11:0] a;
    reg [15:0] rom [4095:0];
    always @(posedge clk) q <= rom[a];
    integer i;
    initial
    begin
        for (i=0; i < 4096; i=i+1)
        begin
            rom[i] = 0;
        end
    
        rom[0] = 28672;
rom[1] = 839;
rom[2] = 4992;
rom[3] = 1863;
rom[4] = 2887;
rom[5] = 7104;
rom[6] = 3587;
rom[7] = 7713;
rom[8] = 6912;
rom[9] = 7104;
rom[10] = 7713;
rom[11] = 6912;
rom[12] = 7104;
rom[13] = 7713;
rom[14] = 6912;
rom[15] = 7040;
rom[16] = 5411;
rom[17] = 4864;
rom[18] = 52741;
rom[19] = 327;
rom[20] = 1027;
rom[21] = 52737;
rom[22] = 839;
rom[23] = 4992;
rom[24] = 1863;
rom[25] = 52743;
rom[26] = 2887;
rom[27] = 7104;
rom[28] = 3587;
rom[29] = 7713;
rom[30] = 6912;
rom[31] = 7104;
rom[32] = 7713;
rom[33] = 6912;
rom[34] = 7104;
rom[35] = 7713;
rom[36] = 6912;
rom[37] = 7104;
rom[38] = 7713;
rom[39] = 6912;
rom[40] = 7104;
rom[41] = 7713;
rom[42] = 6912;
rom[43] = 50693;
rom[44] = 837;
rom[45] = 1537;
rom[46] = 5056;
rom[47] = 7040;
rom[48] = 5155;
rom[49] = 4864;
rom[50] = 52745;
rom[51] = 327;
rom[52] = 1027;
rom[53] = 52737;
rom[54] = 839;
rom[55] = 4992;
rom[56] = 1863;
rom[57] = 52747;
rom[58] = 2887;
rom[59] = 7104;
rom[60] = 3587;
rom[61] = 7713;
rom[62] = 6912;
rom[63] = 7104;
rom[64] = 7713;
rom[65] = 6912;
rom[66] = 7104;
rom[67] = 7713;
rom[68] = 6912;
rom[69] = 7104;
rom[70] = 7713;
rom[71] = 6912;
rom[72] = 7104;
rom[73] = 7713;
rom[74] = 6912;
rom[75] = 7104;
rom[76] = 7713;
rom[77] = 6912;
rom[78] = 7104;
rom[79] = 7713;
rom[80] = 6912;
rom[81] = 50697;
rom[82] = 837;
rom[83] = 1537;
rom[84] = 5056;
rom[85] = 7040;
rom[86] = 5411;
rom[87] = 4864;
rom[88] = 52749;
rom[89] = 327;
rom[90] = 1027;
rom[91] = 28672;
    end
    endmodule
     
module main (
	clk);
input clk;
reg  [11:0] v$INT0_15885_out0 = 12'h0;
reg  [11:0] v$INT0_15886_out0 = 12'h0;
reg  [11:0] v$INT1_18533_out0 = 12'h0;
reg  [11:0] v$INT1_18534_out0 = 12'h0;
reg  [11:0] v$INT2_256_out0 = 12'h0;
reg  [11:0] v$INT2_257_out0 = 12'h0;
reg  [11:0] v$INT3_271_out0 = 12'h0;
reg  [11:0] v$INT3_272_out0 = 12'h0;
reg  [11:0] v$PCINTERRUPT_17807_out0 = 12'h0;
reg  [11:0] v$PCINTERRUPT_17808_out0 = 12'h0;
reg  [11:0] v$PCNORMAL_12768_out0 = 12'h0;
reg  [11:0] v$PCNORMAL_12769_out0 = 12'h0;
reg  [11:0] v$REG12_3330_out0 = 12'h0;
reg  [11:0] v$REG9_16088_out0 = 12'h0;
reg  [15:0] v$REG0_16254_out0 = 16'h0;
reg  [15:0] v$REG0_16255_out0 = 16'h0;
reg  [15:0] v$REG10_16463_out0 = 16'h0;
reg  [15:0] v$REG11_9622_out0 = 16'h0;
reg  [15:0] v$REG1_1163_out0 = 16'h0;
reg  [15:0] v$REG1_1164_out0 = 16'h0;
reg  [15:0] v$REG1_13592_out0 = 16'h0;
reg  [15:0] v$REG1_13593_out0 = 16'h0;
reg  [15:0] v$REG1_14099_out0 = 16'h0;
reg  [15:0] v$REG1_14100_out0 = 16'h0;
reg  [15:0] v$REG1_4894_out0 = 16'h0;
reg  [15:0] v$REG1_4895_out0 = 16'h0;
reg  [15:0] v$REG2_15005_out0 = 16'h0;
reg  [15:0] v$REG2_15006_out0 = 16'h0;
reg  [15:0] v$REG2_15617_out0 = 16'h0;
reg  [15:0] v$REG2_15618_out0 = 16'h0;
reg  [15:0] v$REG2_16345_out0 = 16'h0;
reg  [15:0] v$REG2_16346_out0 = 16'h0;
reg  [15:0] v$REG2_17480_out0 = 16'h0;
reg  [15:0] v$REG2_17481_out0 = 16'h0;
reg  [15:0] v$REG3_11001_out0 = 16'h0;
reg  [15:0] v$REG3_11002_out0 = 16'h0;
reg  [15:0] v$REG3_11767_out0 = 16'h0;
reg  [15:0] v$REG3_11768_out0 = 16'h0;
reg  [15:0] v$REG3_2822_out0 = 16'h0;
reg  [15:0] v$REG3_2823_out0 = 16'h0;
reg  [15:0] v$REG4_6650_out0 = 16'h0;
reg  [15:0] v$REG4_6651_out0 = 16'h0;
reg  [1:0] v$REG1_10904_out0 = 2'h0;
reg  [1:0] v$REG1_10905_out0 = 2'h0;
reg  [1:0] v$REG4_10777_out0 = 2'h0;
reg  [23:0] v$REG1_12089_out0 = 24'h0;
reg  [23:0] v$REG2_16798_out0 = 24'h0;
reg  [31:0] v$REG1_7848_out0 = 32'h0;
reg  [31:0] v$REG2_4047_out0 = 32'h0;
reg  [35:0] v$REG3_6998_out0 = 36'h0;
reg  [3:0] v$REG1_18662_out0 = 4'h0;
reg  [3:0] v$REG1_18663_out0 = 4'h0;
reg  [3:0] v$REG1_8890_out0 = 4'h0;
reg  [3:0] v$REG1_8891_out0 = 4'h0;
reg  [4:0] v$REG1_14090_out0 = 5'h0;
reg  [5:0] v$REG1_14834_out0 = 6'h0;
reg  [5:0] v$REG1_14835_out0 = 6'h0;
reg  [5:0] v$REG2_657_out0 = 6'h0;
reg  [5:0] v$REG2_658_out0 = 6'h0;
reg  [7:0] v$REG1_10302_out0 = 8'h0;
reg  [7:0] v$REG1_10303_out0 = 8'h0;
reg  [7:0] v$REG1_4043_out0 = 8'h0;
reg  [7:0] v$REG1_4044_out0 = 8'h0;
reg v$FF0_4326_out0 = 1'b0;
reg v$FF0_4327_out0 = 1'b0;
reg v$FF0_5007_out0 = 1'b0;
reg v$FF0_5008_out0 = 1'b0;
reg v$FF0_655_out0 = 1'b0;
reg v$FF0_656_out0 = 1'b0;
reg v$FF0_9401_out0 = 1'b0;
reg v$FF0_9402_out0 = 1'b0;
reg v$FF10_14203_out0 = 1'b0;
reg v$FF10_14204_out0 = 1'b0;
reg v$FF10_7890_out0 = 1'b0;
reg v$FF10_7891_out0 = 1'b0;
reg v$FF11_2449_out0 = 1'b0;
reg v$FF11_2450_out0 = 1'b0;
reg v$FF12_16427_out0 = 1'b0;
reg v$FF12_16428_out0 = 1'b0;
reg v$FF13_18541_out0 = 1'b0;
reg v$FF13_18542_out0 = 1'b0;
reg v$FF14_10906_out0 = 1'b0;
reg v$FF14_10907_out0 = 1'b0;
reg v$FF15_12716_out0 = 1'b0;
reg v$FF15_12717_out0 = 1'b0;
reg v$FF1_10306_out0 = 1'b0;
reg v$FF1_10307_out0 = 1'b0;
reg v$FF1_11054_out0 = 1'b0;
reg v$FF1_11055_out0 = 1'b0;
reg v$FF1_1178_out0 = 1'b0;
reg v$FF1_1179_out0 = 1'b0;
reg v$FF1_13095_out0 = 1'b0;
reg v$FF1_13096_out0 = 1'b0;
reg v$FF1_13680_out0 = 1'b0;
reg v$FF1_13681_out0 = 1'b0;
reg v$FF1_1376_out0 = 1'b0;
reg v$FF1_1377_out0 = 1'b0;
reg v$FF1_16074_out0 = 1'b0;
reg v$FF1_16075_out0 = 1'b0;
reg v$FF1_16076_out0 = 1'b0;
reg v$FF1_16077_out0 = 1'b0;
reg v$FF1_16078_out0 = 1'b0;
reg v$FF1_16079_out0 = 1'b0;
reg v$FF1_16080_out0 = 1'b0;
reg v$FF1_16081_out0 = 1'b0;
reg v$FF1_16082_out0 = 1'b0;
reg v$FF1_16083_out0 = 1'b0;
reg v$FF1_16084_out0 = 1'b0;
reg v$FF1_16085_out0 = 1'b0;
reg v$FF1_16187_out0 = 1'b0;
reg v$FF1_16188_out0 = 1'b0;
reg v$FF1_16315_out0 = 1'b0;
reg v$FF1_16316_out0 = 1'b0;
reg v$FF1_191_out0 = 1'b0;
reg v$FF1_192_out0 = 1'b0;
reg v$FF1_2525_out0 = 1'b0;
reg v$FF1_2526_out0 = 1'b0;
reg v$FF1_2_out0 = 1'b0;
reg v$FF1_3_out0 = 1'b0;
reg v$FF1_4339_out0 = 1'b0;
reg v$FF1_5226_out0 = 1'b0;
reg v$FF1_5227_out0 = 1'b0;
reg v$FF1_5228_out0 = 1'b0;
reg v$FF1_5229_out0 = 1'b0;
reg v$FF1_5448_out0 = 1'b0;
reg v$FF1_6026_out0 = 1'b0;
reg v$FF1_6027_out0 = 1'b0;
reg v$FF1_6149_out0 = 1'b0;
reg v$FF1_6150_out0 = 1'b0;
reg v$FF1_8223_out0 = 1'b0;
reg v$FF1_8224_out0 = 1'b0;
reg v$FF1_9422_out0 = 1'b0;
reg v$FF1_9423_out0 = 1'b0;
reg v$FF1_9607_out0 = 1'b0;
reg v$FF1_9608_out0 = 1'b0;
reg v$FF1_9630_out0 = 1'b0;
reg v$FF1_9631_out0 = 1'b0;
reg v$FF2_1180_out0 = 1'b0;
reg v$FF2_1181_out0 = 1'b0;
reg v$FF2_13039_out0 = 1'b0;
reg v$FF2_13040_out0 = 1'b0;
reg v$FF2_13041_out0 = 1'b0;
reg v$FF2_13042_out0 = 1'b0;
reg v$FF2_13043_out0 = 1'b0;
reg v$FF2_13044_out0 = 1'b0;
reg v$FF2_13045_out0 = 1'b0;
reg v$FF2_13046_out0 = 1'b0;
reg v$FF2_13047_out0 = 1'b0;
reg v$FF2_13048_out0 = 1'b0;
reg v$FF2_13049_out0 = 1'b0;
reg v$FF2_13050_out0 = 1'b0;
reg v$FF2_13051_out0 = 1'b0;
reg v$FF2_13052_out0 = 1'b0;
reg v$FF2_13053_out0 = 1'b0;
reg v$FF2_13054_out0 = 1'b0;
reg v$FF2_13055_out0 = 1'b0;
reg v$FF2_13056_out0 = 1'b0;
reg v$FF2_13057_out0 = 1'b0;
reg v$FF2_13058_out0 = 1'b0;
reg v$FF2_13059_out0 = 1'b0;
reg v$FF2_13060_out0 = 1'b0;
reg v$FF2_13458_out0 = 1'b0;
reg v$FF2_14629_out0 = 1'b0;
reg v$FF2_14630_out0 = 1'b0;
reg v$FF2_14782_out0 = 1'b0;
reg v$FF2_14783_out0 = 1'b0;
reg v$FF2_14784_out0 = 1'b0;
reg v$FF2_14785_out0 = 1'b0;
reg v$FF2_14786_out0 = 1'b0;
reg v$FF2_14787_out0 = 1'b0;
reg v$FF2_14788_out0 = 1'b0;
reg v$FF2_14789_out0 = 1'b0;
reg v$FF2_14790_out0 = 1'b0;
reg v$FF2_14791_out0 = 1'b0;
reg v$FF2_14792_out0 = 1'b0;
reg v$FF2_14793_out0 = 1'b0;
reg v$FF2_15481_out0 = 1'b0;
reg v$FF2_15482_out0 = 1'b0;
reg v$FF2_1572_out0 = 1'b0;
reg v$FF2_1573_out0 = 1'b0;
reg v$FF2_16336_out0 = 1'b0;
reg v$FF2_16337_out0 = 1'b0;
reg v$FF2_16652_out0 = 1'b0;
reg v$FF2_16653_out0 = 1'b0;
reg v$FF2_2951_out0 = 1'b0;
reg v$FF2_2952_out0 = 1'b0;
reg v$FF2_4345_out0 = 1'b0;
reg v$FF2_4346_out0 = 1'b0;
reg v$FF2_9418_out0 = 1'b0;
reg v$FF2_9419_out0 = 1'b0;
reg v$FF3_10915_out0 = 1'b0;
reg v$FF3_10916_out0 = 1'b0;
reg v$FF3_1296_out0 = 1'b0;
reg v$FF3_1297_out0 = 1'b0;
reg v$FF3_15030_out0 = 1'b0;
reg v$FF3_15031_out0 = 1'b0;
reg v$FF3_15956_out0 = 1'b0;
reg v$FF3_15957_out0 = 1'b0;
reg v$FF3_18116_out0 = 1'b0;
reg v$FF3_18117_out0 = 1'b0;
reg v$FF3_262_out0 = 1'b0;
reg v$FF3_263_out0 = 1'b0;
reg v$FF3_3378_out0 = 1'b0;
reg v$FF3_7331_out0 = 1'b0;
reg v$FF3_7332_out0 = 1'b0;
reg v$FF3_7563_out0 = 1'b0;
reg v$FF3_7564_out0 = 1'b0;
reg v$FF3_9971_out0 = 1'b0;
reg v$FF3_9972_out0 = 1'b0;
reg v$FF3_9973_out0 = 1'b0;
reg v$FF3_9974_out0 = 1'b0;
reg v$FF3_9975_out0 = 1'b0;
reg v$FF3_9976_out0 = 1'b0;
reg v$FF3_9977_out0 = 1'b0;
reg v$FF3_9978_out0 = 1'b0;
reg v$FF3_9979_out0 = 1'b0;
reg v$FF3_9980_out0 = 1'b0;
reg v$FF3_9981_out0 = 1'b0;
reg v$FF3_9982_out0 = 1'b0;
reg v$FF4_13548_out0 = 1'b0;
reg v$FF4_15974_out0 = 1'b0;
reg v$FF4_15975_out0 = 1'b0;
reg v$FF4_15976_out0 = 1'b0;
reg v$FF4_15977_out0 = 1'b0;
reg v$FF4_15978_out0 = 1'b0;
reg v$FF4_15979_out0 = 1'b0;
reg v$FF4_15980_out0 = 1'b0;
reg v$FF4_15981_out0 = 1'b0;
reg v$FF4_15982_out0 = 1'b0;
reg v$FF4_15983_out0 = 1'b0;
reg v$FF4_15984_out0 = 1'b0;
reg v$FF4_15985_out0 = 1'b0;
reg v$FF4_17846_out0 = 1'b0;
reg v$FF4_17847_out0 = 1'b0;
reg v$FF4_18438_out0 = 1'b0;
reg v$FF4_18439_out0 = 1'b0;
reg v$FF4_2347_out0 = 1'b0;
reg v$FF4_2348_out0 = 1'b0;
reg v$FF4_3781_out0 = 1'b0;
reg v$FF4_3782_out0 = 1'b0;
reg v$FF4_7017_out0 = 1'b0;
reg v$FF4_7018_out0 = 1'b0;
reg v$FF4_8055_out0 = 1'b0;
reg v$FF4_8056_out0 = 1'b0;
reg v$FF4_8252_out0 = 1'b0;
reg v$FF4_8253_out0 = 1'b0;
reg v$FF5_16338_out0 = 1'b0;
reg v$FF5_16339_out0 = 1'b0;
reg v$FF5_16426_out0 = 1'b0;
reg v$FF5_1754_out0 = 1'b0;
reg v$FF5_1755_out0 = 1'b0;
reg v$FF5_1756_out0 = 1'b0;
reg v$FF5_1757_out0 = 1'b0;
reg v$FF5_1758_out0 = 1'b0;
reg v$FF5_1759_out0 = 1'b0;
reg v$FF5_1760_out0 = 1'b0;
reg v$FF5_1761_out0 = 1'b0;
reg v$FF5_1762_out0 = 1'b0;
reg v$FF5_1763_out0 = 1'b0;
reg v$FF5_1764_out0 = 1'b0;
reg v$FF5_1765_out0 = 1'b0;
reg v$FF5_18473_out0 = 1'b0;
reg v$FF5_18474_out0 = 1'b0;
reg v$FF5_4744_out0 = 1'b0;
reg v$FF5_4745_out0 = 1'b0;
reg v$FF6_15324_out0 = 1'b0;
reg v$FF6_15325_out0 = 1'b0;
reg v$FF6_16171_out0 = 1'b0;
reg v$FF6_2621_out0 = 1'b0;
reg v$FF6_2622_out0 = 1'b0;
reg v$FF6_2623_out0 = 1'b0;
reg v$FF6_2624_out0 = 1'b0;
reg v$FF6_2625_out0 = 1'b0;
reg v$FF6_2626_out0 = 1'b0;
reg v$FF6_2627_out0 = 1'b0;
reg v$FF6_2628_out0 = 1'b0;
reg v$FF6_2629_out0 = 1'b0;
reg v$FF6_2630_out0 = 1'b0;
reg v$FF6_2631_out0 = 1'b0;
reg v$FF6_2632_out0 = 1'b0;
reg v$FF6_8963_out0 = 1'b0;
reg v$FF6_8964_out0 = 1'b0;
reg v$FF7_12756_out0 = 1'b0;
reg v$FF7_12757_out0 = 1'b0;
reg v$FF7_14553_out0 = 1'b0;
reg v$FF7_14554_out0 = 1'b0;
reg v$FF7_18120_out0 = 1'b0;
reg v$FF7_18121_out0 = 1'b0;
reg v$FF7_8087_out0 = 1'b0;
reg v$FF7_8088_out0 = 1'b0;
reg v$FF7_8298_out0 = 1'b0;
reg v$FF7_8299_out0 = 1'b0;
reg v$FF7_8300_out0 = 1'b0;
reg v$FF7_8301_out0 = 1'b0;
reg v$FF7_8302_out0 = 1'b0;
reg v$FF7_8303_out0 = 1'b0;
reg v$FF7_8304_out0 = 1'b0;
reg v$FF7_8305_out0 = 1'b0;
reg v$FF7_8306_out0 = 1'b0;
reg v$FF7_8307_out0 = 1'b0;
reg v$FF7_8308_out0 = 1'b0;
reg v$FF7_8309_out0 = 1'b0;
reg v$FF8_10337_out0 = 1'b0;
reg v$FF8_10338_out0 = 1'b0;
reg v$FF8_14460_out0 = 1'b0;
reg v$FF8_14461_out0 = 1'b0;
reg v$FF8_14462_out0 = 1'b0;
reg v$FF8_14463_out0 = 1'b0;
reg v$FF8_14464_out0 = 1'b0;
reg v$FF8_14465_out0 = 1'b0;
reg v$FF8_14466_out0 = 1'b0;
reg v$FF8_14467_out0 = 1'b0;
reg v$FF8_14468_out0 = 1'b0;
reg v$FF8_14469_out0 = 1'b0;
reg v$FF8_14470_out0 = 1'b0;
reg v$FF8_14471_out0 = 1'b0;
reg v$FF8_16727_out0 = 1'b0;
reg v$FF8_16728_out0 = 1'b0;
reg v$FF8_8026_out0 = 1'b0;
reg v$FF8_8027_out0 = 1'b0;
reg v$FF9_10664_out0 = 1'b0;
reg v$FF9_10665_out0 = 1'b0;
reg v$FF9_16021_out0 = 1'b0;
reg v$FF9_16022_out0 = 1'b0;
reg v$LSB$FF_18514_out0 = 1'b0;
reg v$LSB$FF_18515_out0 = 1'b0;
reg v$REG13_296_out0 = 1'b0;
reg v$REG14_5459_out0 = 1'b0;
reg v$REG1_7074_out0 = 1'b0;
reg v$REG1_8824_out0 = 1'b0;
reg v$REG2_11798_out0 = 1'b0;
reg v$REG2_11799_out0 = 1'b0;
reg v$REG2_18373_out0 = 1'b0;
reg v$REG2_5128_out0 = 1'b0;
reg v$REG3_17753_out0 = 1'b0;
reg v$REG3_17754_out0 = 1'b0;
reg v$REG4_10994_out0 = 1'b0;
reg v$REG7_6181_out0 = 1'b0;
reg v$REG8_4106_out0 = 1'b0;
reg v$S$FF_10816_out0 = 1'b0;
reg v$S$FF_10817_out0 = 1'b0;
wire  [10:0] v$C1_15804_out0;
wire  [10:0] v$C1_15805_out0;
wire  [10:0] v$SEL5_16175_out0;
wire  [10:0] v$SEL5_16176_out0;
wire  [11:0] v$A1_14820_out0;
wire  [11:0] v$A1_14821_out0;
wire  [11:0] v$ADDRESS_15194_out0;
wire  [11:0] v$ADDRESS_15195_out0;
wire  [11:0] v$ADDRESS_15901_out0;
wire  [11:0] v$ADDRESS_15902_out0;
wire  [11:0] v$ADDRESS_5811_out0;
wire  [11:0] v$ADDRESS_5812_out0;
wire  [11:0] v$ADD_2955_out0;
wire  [11:0] v$ADD_2956_out0;
wire  [11:0] v$A_2543_out0;
wire  [11:0] v$A_2544_out0;
wire  [11:0] v$A_2545_out0;
wire  [11:0] v$A_2546_out0;
wire  [11:0] v$B_12130_out0;
wire  [11:0] v$B_12131_out0;
wire  [11:0] v$B_12132_out0;
wire  [11:0] v$B_12133_out0;
wire  [11:0] v$C1_15940_out0;
wire  [11:0] v$C1_15941_out0;
wire  [11:0] v$C4_15906_out0;
wire  [11:0] v$C4_15907_out0;
wire  [11:0] v$END_16598_out0;
wire  [11:0] v$END_16599_out0;
wire  [11:0] v$MUX1_1851_out0;
wire  [11:0] v$MUX2_3722_out0;
wire  [11:0] v$MUX2_3723_out0;
wire  [11:0] v$MUX3_9123_out0;
wire  [11:0] v$MUX4_1574_out0;
wire  [11:0] v$MUX4_1575_out0;
wire  [11:0] v$MUX5_16988_out0;
wire  [11:0] v$MUX5_16989_out0;
wire  [11:0] v$MUX6_14420_out0;
wire  [11:0] v$MUX6_14421_out0;
wire  [11:0] v$MUX6_6903_out0;
wire  [11:0] v$MUX7_1135_out0;
wire  [11:0] v$MUX7_1136_out0;
wire  [11:0] v$MUX8_12286_out0;
wire  [11:0] v$MUX8_12287_out0;
wire  [11:0] v$N$VIEWER_1615_out0;
wire  [11:0] v$N$VIEWER_1616_out0;
wire  [11:0] v$NEXTINSTRUCTIONADDRESS_18408_out0;
wire  [11:0] v$NEXTINSTRUCTIONADDRESS_18409_out0;
wire  [11:0] v$N_11753_out0;
wire  [11:0] v$N_11754_out0;
wire  [11:0] v$N_11963_out0;
wire  [11:0] v$N_11964_out0;
wire  [11:0] v$N_14507_out0;
wire  [11:0] v$N_14508_out0;
wire  [11:0] v$N_14843_out0;
wire  [11:0] v$N_14844_out0;
wire  [11:0] v$N_1621_out0;
wire  [11:0] v$N_1622_out0;
wire  [11:0] v$N_17937_out0;
wire  [11:0] v$N_17938_out0;
wire  [11:0] v$N_18295_out0;
wire  [11:0] v$N_18296_out0;
wire  [11:0] v$N_8269_out0;
wire  [11:0] v$N_8270_out0;
wire  [11:0] v$PC$NEXT0_1935_out0;
wire  [11:0] v$PC$NEXT1_3497_out0;
wire  [11:0] v$PCNEXT$VIEWER_15772_out0;
wire  [11:0] v$PCNEXT$VIEWER_15773_out0;
wire  [11:0] v$PCNEXT_6654_out0;
wire  [11:0] v$PCNEXT_6655_out0;
wire  [11:0] v$PC_3147_out0;
wire  [11:0] v$PC_3148_out0;
wire  [11:0] v$RAM$ADDR$VIEWER_15934_out0;
wire  [11:0] v$RAM$ADDR$VIEWER_15935_out0;
wire  [11:0] v$RAM$ADDR0_12525_out0;
wire  [11:0] v$RAM$ADDR1_6454_out0;
wire  [11:0] v$RAM$ADDR_15228_out0;
wire  [11:0] v$RAM$ADDR_15229_out0;
wire  [11:0] v$RAM$ADDR_6413_out0;
wire  [11:0] v$RAM$ADDR_6414_out0;
wire  [11:0] v$RAMADDR0_16982_out0;
wire  [11:0] v$RAMADDR1_12657_out0;
wire  [11:0] v$RAMADDRESS_12721_out0;
wire  [11:0] v$RAMADDRESS_12722_out0;
wire  [11:0] v$RAMADDRESS_6988_out0;
wire  [11:0] v$RAMADDRESS_6989_out0;
wire  [11:0] v$RAMADDRMUX_14376_out0;
wire  [11:0] v$RAMADDRMUX_14377_out0;
wire  [11:0] v$RAMADDRMUX_418_out0;
wire  [11:0] v$RAMADDRMUX_419_out0;
wire  [11:0] v$RAMADDRMUX_4746_out0;
wire  [11:0] v$RAMADDRMUX_4747_out0;
wire  [11:0] v$RAMADDRMUX_4816_out0;
wire  [11:0] v$RAMADDRMUX_4817_out0;
wire  [11:0] v$RAMADDR_13607_out0;
wire  [11:0] v$RAMADDR_18656_out0;
wire  [11:0] v$RAMADDR_8766_out0;
wire  [11:0] v$RAMAddress_2262_out0;
wire  [11:0] v$RAMAddress_2263_out0;
wire  [11:0] v$SEL1_11971_out0;
wire  [11:0] v$SEL1_11972_out0;
wire  [11:0] v$SEL1_3249_out0;
wire  [11:0] v$SEL1_3250_out0;
wire  [11:0] v$SEL2_13746_out0;
wire  [11:0] v$SEL2_13747_out0;
wire  [11:0] v$SEL3_1251_out0;
wire  [11:0] v$SEL3_1252_out0;
wire  [11:0] v$SEL4_1364_out0;
wire  [11:0] v$SEL4_1365_out0;
wire  [11:0] v$SEL8_12749_out0;
wire  [11:0] v$SUM_13667_out0;
wire  [11:0] v$SUM_13668_out0;
wire  [11:0] v$_14024_out0;
wire  [11:0] v$_14025_out0;
wire  [11:0] v$_14601_out0;
wire  [11:0] v$_14605_out0;
wire  [11:0] v$_14635_out0;
wire  [11:0] v$_14639_out0;
wire  [11:0] v$_16367_out0;
wire  [11:0] v$_16368_out0;
wire  [11:0] v$_16749_out0;
wire  [11:0] v$_16753_out0;
wire  [11:0] v$_3985_out0;
wire  [11:0] v$_3985_out1;
wire  [11:0] v$_3986_out0;
wire  [11:0] v$_3986_out1;
wire  [11:0] v$_3987_out0;
wire  [11:0] v$_3987_out1;
wire  [11:0] v$_3988_out0;
wire  [11:0] v$_3988_out1;
wire  [11:0] v$_3989_out0;
wire  [11:0] v$_3989_out1;
wire  [11:0] v$_4802_out0;
wire  [11:0] v$_4806_out0;
wire  [11:0] v$_7539_out0;
wire  [11:0] v$_7539_out1;
wire  [11:0] v$_7540_out0;
wire  [11:0] v$_7540_out1;
wire  [11:0] v$_7541_out0;
wire  [11:0] v$_7541_out1;
wire  [11:0] v$_7542_out0;
wire  [11:0] v$_7542_out1;
wire  [11:0] v$_7543_out0;
wire  [11:0] v$_7543_out1;
wire  [11:0] v$_7720_out0;
wire  [11:0] v$_7721_out0;
wire  [12:0] v$C10_8949_out0;
wire  [12:0] v$C10_8950_out0;
wire  [12:0] v$C4_2451_out0;
wire  [12:0] v$C4_2452_out0;
wire  [12:0] v$C6_1535_out0;
wire  [12:0] v$C6_1536_out0;
wire  [12:0] v$C7_6037_out0;
wire  [12:0] v$C7_6038_out0;
wire  [12:0] v$C8_8206_out0;
wire  [12:0] v$C8_8207_out0;
wire  [13:0] v$_14600_out0;
wire  [13:0] v$_14604_out0;
wire  [13:0] v$_14634_out0;
wire  [13:0] v$_14638_out0;
wire  [13:0] v$_16748_out0;
wire  [13:0] v$_16752_out0;
wire  [13:0] v$_4801_out0;
wire  [13:0] v$_4805_out0;
wire  [14:0] v$C2_18012_out0;
wire  [14:0] v$C2_18013_out0;
wire  [14:0] v$C4_8256_out0;
wire  [14:0] v$C4_8258_out0;
wire  [14:0] v$MUX2_13630_out0;
wire  [14:0] v$MUX2_13632_out0;
wire  [14:0] v$SEL2_6165_out0;
wire  [14:0] v$SEL2_6166_out0;
wire  [14:0] v$_11383_out0;
wire  [14:0] v$_11384_out0;
wire  [14:0] v$_14599_out0;
wire  [14:0] v$_14603_out0;
wire  [14:0] v$_14633_out0;
wire  [14:0] v$_14637_out0;
wire  [14:0] v$_15153_out0;
wire  [14:0] v$_15154_out0;
wire  [14:0] v$_15846_out0;
wire  [14:0] v$_15848_out0;
wire  [14:0] v$_16747_out0;
wire  [14:0] v$_16751_out0;
wire  [14:0] v$_4800_out0;
wire  [14:0] v$_4804_out0;
wire  [15:0] v$A$COMPARATOR$IN_1467_out0;
wire  [15:0] v$A$COMPARATOR$IN_1468_out0;
wire  [15:0] v$A$IN$MULTIPLIER_4076_out0;
wire  [15:0] v$A$IN$MULTIPLIER_4077_out0;
wire  [15:0] v$A$SAVED$PIPELINED_16524_out0;
wire  [15:0] v$A$SAVED_14631_out0;
wire  [15:0] v$A$SAVED_14632_out0;
wire  [15:0] v$A$SAVED_16525_out0;
wire  [15:0] v$A$SAVED_3698_out0;
wire  [15:0] v$A$SAVED_3699_out0;
wire  [15:0] v$A$SAVED_9967_out0;
wire  [15:0] v$A$SAVED_9968_out0;
wire  [15:0] v$A$VIEW_16308_out0;
wire  [15:0] v$A$VIEW_16309_out0;
wire  [15:0] v$A1_13701_out0;
wire  [15:0] v$A1_13702_out0;
wire  [15:0] v$A1_6409_out0;
wire  [15:0] v$A1_6410_out0;
wire  [15:0] v$A1_9430_out0;
wire  [15:0] v$A1_9431_out0;
wire  [15:0] v$ADDEROUT_3504_out0;
wire  [15:0] v$ADDEROUT_3505_out0;
wire  [15:0] v$ALUOUT$LOADSTORE_18633_out0;
wire  [15:0] v$ALUOUT$LOADSTORE_18634_out0;
wire  [15:0] v$ALUOUT_10219_out0;
wire  [15:0] v$ALUOUT_10220_out0;
wire  [15:0] v$ALUOUT_16542_out0;
wire  [15:0] v$ALUOUT_16543_out0;
wire  [15:0] v$ALUOUT_18072_out0;
wire  [15:0] v$ALUOUT_18073_out0;
wire  [15:0] v$ALUOUT_5760_out0;
wire  [15:0] v$ALUOUT_5761_out0;
wire  [15:0] v$ALUOUT_6922_out0;
wire  [15:0] v$ALUOUT_6923_out0;
wire  [15:0] v$ANDOUT_7376_out0;
wire  [15:0] v$ANDOUT_7377_out0;
wire  [15:0] v$A_11042_out0;
wire  [15:0] v$A_11043_out0;
wire  [15:0] v$A_13811_out0;
wire  [15:0] v$A_13813_out0;
wire  [15:0] v$A_13815_out0;
wire  [15:0] v$A_13817_out0;
wire  [15:0] v$A_16090_out0;
wire  [15:0] v$A_16420_out0;
wire  [15:0] v$A_16421_out0;
wire  [15:0] v$A_17045_out0;
wire  [15:0] v$A_17046_out0;
wire  [15:0] v$A_18293_out0;
wire  [15:0] v$A_18294_out0;
wire  [15:0] v$A_2293_out0;
wire  [15:0] v$A_2547_out0;
wire  [15:0] v$A_2548_out0;
wire  [15:0] v$A_3242_out0;
wire  [15:0] v$A_3243_out0;
wire  [15:0] v$A_4196_out0;
wire  [15:0] v$A_4197_out0;
wire  [15:0] v$A_8693_out0;
wire  [15:0] v$A_8694_out0;
wire  [15:0] v$A_9404_out0;
wire  [15:0] v$A_9405_out0;
wire  [15:0] v$B$COMPARATOR$IN_17962_out0;
wire  [15:0] v$B$COMPARATOR$IN_17963_out0;
wire  [15:0] v$B$IN$MULTIPLIER_15471_out0;
wire  [15:0] v$B$IN$MULTIPLIER_15472_out0;
wire  [15:0] v$B$IN_11650_out0;
wire  [15:0] v$B$IN_11651_out0;
wire  [15:0] v$B$MERGE_16587_out0;
wire  [15:0] v$B$MERGE_16588_out0;
wire  [15:0] v$B$SAVED$PIPELINED_17730_out0;
wire  [15:0] v$B$SAVED_17731_out0;
wire  [15:0] v$B$SAVED_3884_out0;
wire  [15:0] v$B$SAVED_3885_out0;
wire  [15:0] v$B$SAVED_4358_out0;
wire  [15:0] v$B$SAVED_4359_out0;
wire  [15:0] v$B$SAVED_4748_out0;
wire  [15:0] v$B$SAVED_4749_out0;
wire  [15:0] v$B_10007_out0;
wire  [15:0] v$B_10008_out0;
wire  [15:0] v$B_11720_out0;
wire  [15:0] v$B_11721_out0;
wire  [15:0] v$B_12138_out0;
wire  [15:0] v$B_14066_out0;
wire  [15:0] v$B_14067_out0;
wire  [15:0] v$B_17051_out0;
wire  [15:0] v$B_17052_out0;
wire  [15:0] v$B_17746_out0;
wire  [15:0] v$B_17747_out0;
wire  [15:0] v$B_17974_out0;
wire  [15:0] v$B_17975_out0;
wire  [15:0] v$B_18099_out0;
wire  [15:0] v$B_18100_out0;
wire  [15:0] v$B_3366_out0;
wire  [15:0] v$B_3367_out0;
wire  [15:0] v$B_4825_out0;
wire  [15:0] v$B_4827_out0;
wire  [15:0] v$B_4829_out0;
wire  [15:0] v$B_4831_out0;
wire  [15:0] v$B_6548_out0;
wire  [15:0] v$C10_6384_out0;
wire  [15:0] v$C10_6385_out0;
wire  [15:0] v$C1_16322_out0;
wire  [15:0] v$C1_16323_out0;
wire  [15:0] v$C1_18208_out0;
wire  [15:0] v$C1_18209_out0;
wire  [15:0] v$C1_5961_out0;
wire  [15:0] v$C1_5966_out0;
wire  [15:0] v$C1_5971_out0;
wire  [15:0] v$C1_5979_out0;
wire  [15:0] v$C1_5981_out0;
wire  [15:0] v$C1_5989_out0;
wire  [15:0] v$C1_5992_out0;
wire  [15:0] v$C1_6000_out0;
wire  [15:0] v$C1_6006_out0;
wire  [15:0] v$C1_6009_out0;
wire  [15:0] v$C1_6014_out0;
wire  [15:0] v$C1_6019_out0;
wire  [15:0] v$C2_10009_out0;
wire  [15:0] v$C2_10010_out0;
wire  [15:0] v$C2_103_out0;
wire  [15:0] v$C2_108_out0;
wire  [15:0] v$C2_113_out0;
wire  [15:0] v$C2_121_out0;
wire  [15:0] v$C2_12207_out0;
wire  [15:0] v$C2_12208_out0;
wire  [15:0] v$C2_123_out0;
wire  [15:0] v$C2_131_out0;
wire  [15:0] v$C2_134_out0;
wire  [15:0] v$C2_142_out0;
wire  [15:0] v$C2_148_out0;
wire  [15:0] v$C2_151_out0;
wire  [15:0] v$C2_156_out0;
wire  [15:0] v$C2_161_out0;
wire  [15:0] v$C3_12205_out0;
wire  [15:0] v$C3_12206_out0;
wire  [15:0] v$C7_1708_out0;
wire  [15:0] v$C7_1709_out0;
wire  [15:0] v$C9_18760_out0;
wire  [15:0] v$C9_18761_out0;
wire  [15:0] v$C9_3300_out0;
wire  [15:0] v$C9_3301_out0;
wire  [15:0] v$COUNTERTHRESHOLD_17949_out0;
wire  [15:0] v$COUNTERTHRESHOLD_17950_out0;
wire  [15:0] v$COUNTERVALUE_2986_out0;
wire  [15:0] v$COUNTERVALUE_2987_out0;
wire  [15:0] v$C_18106_out0;
wire  [15:0] v$C_18107_out0;
wire  [15:0] v$DATA$IN0_10404_out0;
wire  [15:0] v$DATA$IN1_15283_out0;
wire  [15:0] v$DATA$IN_1607_out0;
wire  [15:0] v$DATA$IN_1608_out0;
wire  [15:0] v$DATA$IN_7075_out0;
wire  [15:0] v$DATA$IN_7076_out0;
wire  [15:0] v$DATA$OUT0_12300_out0;
wire  [15:0] v$DATA$OUT1_15602_out0;
wire  [15:0] v$DATA$OUT_1307_out0;
wire  [15:0] v$DATA$OUT_1308_out0;
wire  [15:0] v$DATA$OUT_7608_out0;
wire  [15:0] v$DATA$OUT_7609_out0;
wire  [15:0] v$DATAIN0_11058_out0;
wire  [15:0] v$DATAIN1_9634_out0;
wire  [15:0] v$DATAINCP_10990_out0;
wire  [15:0] v$DATAINCP_10991_out0;
wire  [15:0] v$DATA_14086_out0;
wire  [15:0] v$DATA_14087_out0;
wire  [15:0] v$DATA_4354_out0;
wire  [15:0] v$DATA_4355_out0;
wire  [15:0] v$DIN$FIRST$MUX_7494_out0;
wire  [15:0] v$DIN$FIRST$MUX_7495_out0;
wire  [15:0] v$DIN3$VIEWER_2208_out0;
wire  [15:0] v$DIN3$VIEWER_2209_out0;
wire  [15:0] v$DIN3_14418_out0;
wire  [15:0] v$DIN3_14419_out0;
wire  [15:0] v$DIN_1723_out0;
wire  [15:0] v$DIN_1724_out0;
wire  [15:0] v$DIN_1803_out0;
wire  [15:0] v$DIN_1804_out0;
wire  [15:0] v$DM1_7858_out0;
wire  [15:0] v$DM1_7858_out1;
wire  [15:0] v$DOUT1_3157_out0;
wire  [15:0] v$DOUT1_3158_out0;
wire  [15:0] v$DOUT2_3513_out0;
wire  [15:0] v$DOUT2_3514_out0;
wire  [15:0] v$FPU$A_15881_out0;
wire  [15:0] v$FPU$A_15882_out0;
wire  [15:0] v$FPU$B$EN_7012_out0;
wire  [15:0] v$FPU$B_7013_out0;
wire  [15:0] v$FPU$OUT_17011_out0;
wire  [15:0] v$FPU$OUT_17012_out0;
wire  [15:0] v$FPU$OUT_7736_out0;
wire  [15:0] v$HAZ$DECTECTOR$A_17951_out0;
wire  [15:0] v$HAZ$DECTECTOR$A_17952_out0;
wire  [15:0] v$HAZ$DETECTOR$B_5070_out0;
wire  [15:0] v$HAZ$DETECTOR$B_5071_out0;
wire  [15:0] v$INSTR$READ0_14172_out0;
wire  [15:0] v$INSTR$READ1_11970_out0;
wire  [15:0] v$INSTR$READ_14891_out0;
wire  [15:0] v$INSTR$READ_14892_out0;
wire  [15:0] v$INSTR$READ_7221_out0;
wire  [15:0] v$INSTR$READ_7222_out0;
wire  [15:0] v$IN_13563_out0;
wire  [15:0] v$IN_13565_out0;
wire  [15:0] v$IN_13567_out0;
wire  [15:0] v$IN_13568_out0;
wire  [15:0] v$IN_13569_out0;
wire  [15:0] v$IN_13571_out0;
wire  [15:0] v$IN_13572_out0;
wire  [15:0] v$IN_13573_out0;
wire  [15:0] v$IN_193_out0;
wire  [15:0] v$IN_194_out0;
wire  [15:0] v$IN_4360_out0;
wire  [15:0] v$IN_4361_out0;
wire  [15:0] v$IN_4362_out0;
wire  [15:0] v$IN_4363_out0;
wire  [15:0] v$IN_4364_out0;
wire  [15:0] v$IN_4365_out0;
wire  [15:0] v$IN_4366_out0;
wire  [15:0] v$IN_4367_out0;
wire  [15:0] v$IN_9566_out0;
wire  [15:0] v$IN_9567_out0;
wire  [15:0] v$IN_9568_out0;
wire  [15:0] v$IN_9569_out0;
wire  [15:0] v$IN_9570_out0;
wire  [15:0] v$IN_9571_out0;
wire  [15:0] v$IN_9572_out0;
wire  [15:0] v$IN_9573_out0;
wire  [15:0] v$IR$READ$IN$PREV$CYCLE_6188_out0;
wire  [15:0] v$IR$READ$IN$PREV$CYCLE_6189_out0;
wire  [15:0] v$IR1$VIEWER_7428_out0;
wire  [15:0] v$IR1$VIEWER_7429_out0;
wire  [15:0] v$IR1_13389_out0;
wire  [15:0] v$IR1_13390_out0;
wire  [15:0] v$IR1_15998_out0;
wire  [15:0] v$IR1_15999_out0;
wire  [15:0] v$IR1_16680_out0;
wire  [15:0] v$IR1_16681_out0;
wire  [15:0] v$IR1_18034_out0;
wire  [15:0] v$IR1_18035_out0;
wire  [15:0] v$IR1_22_out0;
wire  [15:0] v$IR1_23_out0;
wire  [15:0] v$IR1_4156_out0;
wire  [15:0] v$IR1_4157_out0;
wire  [15:0] v$IR1_646_out0;
wire  [15:0] v$IR1_647_out0;
wire  [15:0] v$IR1_7613_out0;
wire  [15:0] v$IR1_7614_out0;
wire  [15:0] v$IR2$VIEWER_16300_out0;
wire  [15:0] v$IR2$VIEWER_16301_out0;
wire  [15:0] v$IR2_16559_out0;
wire  [15:0] v$IR2_16560_out0;
wire  [15:0] v$IR2_1750_out0;
wire  [15:0] v$IR2_1751_out0;
wire  [15:0] v$IR2_17953_out0;
wire  [15:0] v$IR2_17954_out0;
wire  [15:0] v$IR2_2217_out0;
wire  [15:0] v$IR2_2218_out0;
wire  [15:0] v$IR2_2933_out0;
wire  [15:0] v$IR2_2934_out0;
wire  [15:0] v$IR2_3286_out0;
wire  [15:0] v$IR2_3287_out0;
wire  [15:0] v$IR2_3948_out0;
wire  [15:0] v$IR2_3949_out0;
wire  [15:0] v$IR2_7773_out0;
wire  [15:0] v$IR2_7774_out0;
wire  [15:0] v$LDST$RAMDOUT_1159_out0;
wire  [15:0] v$LDST$RAMDOUT_1160_out0;
wire  [15:0] v$LDST$RMN_7728_out0;
wire  [15:0] v$LDST$RMN_7729_out0;
wire  [15:0] v$LDSTN_3039_out0;
wire  [15:0] v$LDSTN_3040_out0;
wire  [15:0] v$LDSTRM_7644_out0;
wire  [15:0] v$LDSTRM_7645_out0;
wire  [15:0] v$LOAD$STORE$OUT_17575_out0;
wire  [15:0] v$LOAD$STORE$OUT_17576_out0;
wire  [15:0] v$LOWER$PART_7478_out0;
wire  [15:0] v$LOWER$PART_7479_out0;
wire  [15:0] v$MULTIPLY$DENORMALIZATION$16$BIT_11716_out0;
wire  [15:0] v$MULTIPLY$DENORMALIZATION$16$BIT_11717_out0;
wire  [15:0] v$MUX10_16829_out0;
wire  [15:0] v$MUX10_16830_out0;
wire  [15:0] v$MUX11_8669_out0;
wire  [15:0] v$MUX11_8670_out0;
wire  [15:0] v$MUX13_2549_out0;
wire  [15:0] v$MUX13_2550_out0;
wire  [15:0] v$MUX14_18722_out0;
wire  [15:0] v$MUX15_7008_out0;
wire  [15:0] v$MUX15_7009_out0;
wire  [15:0] v$MUX16_18527_out0;
wire  [15:0] v$MUX16_18528_out0;
wire  [15:0] v$MUX1_11751_out0;
wire  [15:0] v$MUX1_11752_out0;
wire  [15:0] v$MUX1_15262_out0;
wire  [15:0] v$MUX1_15263_out0;
wire  [15:0] v$MUX1_17728_out0;
wire  [15:0] v$MUX1_17729_out0;
wire  [15:0] v$MUX1_1811_out0;
wire  [15:0] v$MUX1_1812_out0;
wire  [15:0] v$MUX1_18328_out0;
wire  [15:0] v$MUX1_18329_out0;
wire  [15:0] v$MUX1_1996_out0;
wire  [15:0] v$MUX1_1997_out0;
wire  [15:0] v$MUX1_2603_out0;
wire  [15:0] v$MUX1_2604_out0;
wire  [15:0] v$MUX1_4041_out0;
wire  [15:0] v$MUX1_4042_out0;
wire  [15:0] v$MUX1_5819_out0;
wire  [15:0] v$MUX1_5820_out0;
wire  [15:0] v$MUX1_6677_out0;
wire  [15:0] v$MUX1_6678_out0;
wire  [15:0] v$MUX1_6679_out0;
wire  [15:0] v$MUX1_6680_out0;
wire  [15:0] v$MUX1_6681_out0;
wire  [15:0] v$MUX1_6682_out0;
wire  [15:0] v$MUX1_6683_out0;
wire  [15:0] v$MUX1_6684_out0;
wire  [15:0] v$MUX2_10668_out0;
wire  [15:0] v$MUX2_10669_out0;
wire  [15:0] v$MUX2_11980_out0;
wire  [15:0] v$MUX2_11981_out0;
wire  [15:0] v$MUX2_12038_out0;
wire  [15:0] v$MUX2_12039_out0;
wire  [15:0] v$MUX2_12040_out0;
wire  [15:0] v$MUX2_12041_out0;
wire  [15:0] v$MUX2_12042_out0;
wire  [15:0] v$MUX2_12043_out0;
wire  [15:0] v$MUX2_12044_out0;
wire  [15:0] v$MUX2_12045_out0;
wire  [15:0] v$MUX2_15190_out0;
wire  [15:0] v$MUX2_15191_out0;
wire  [15:0] v$MUX2_15843_out0;
wire  [15:0] v$MUX3_1584_out0;
wire  [15:0] v$MUX3_1585_out0;
wire  [15:0] v$MUX3_18386_out0;
wire  [15:0] v$MUX3_18387_out0;
wire  [15:0] v$MUX3_1957_out0;
wire  [15:0] v$MUX3_1958_out0;
wire  [15:0] v$MUX3_1959_out0;
wire  [15:0] v$MUX3_1960_out0;
wire  [15:0] v$MUX3_1961_out0;
wire  [15:0] v$MUX3_1962_out0;
wire  [15:0] v$MUX3_1963_out0;
wire  [15:0] v$MUX3_1964_out0;
wire  [15:0] v$MUX3_3880_out0;
wire  [15:0] v$MUX3_3881_out0;
wire  [15:0] v$MUX4_15990_out0;
wire  [15:0] v$MUX4_15991_out0;
wire  [15:0] v$MUX4_15992_out0;
wire  [15:0] v$MUX4_15993_out0;
wire  [15:0] v$MUX4_15994_out0;
wire  [15:0] v$MUX4_15995_out0;
wire  [15:0] v$MUX4_15996_out0;
wire  [15:0] v$MUX4_15997_out0;
wire  [15:0] v$MUX4_1651_out0;
wire  [15:0] v$MUX4_1652_out0;
wire  [15:0] v$MUX4_17721_out0;
wire  [15:0] v$MUX4_17722_out0;
wire  [15:0] v$MUX4_3842_out0;
wire  [15:0] v$MUX4_45_out0;
wire  [15:0] v$MUX4_46_out0;
wire  [15:0] v$MUX4_5935_out0;
wire  [15:0] v$MUX4_5936_out0;
wire  [15:0] v$MUX5_10896_out0;
wire  [15:0] v$MUX5_11943_out0;
wire  [15:0] v$MUX5_11944_out0;
wire  [15:0] v$MUX5_14082_out0;
wire  [15:0] v$MUX5_14083_out0;
wire  [15:0] v$MUX6_5051_out0;
wire  [15:0] v$MUX6_5052_out0;
wire  [15:0] v$MUX6_7439_out0;
wire  [15:0] v$MUX6_7440_out0;
wire  [15:0] v$MUX9_17941_out0;
wire  [15:0] v$MUX9_17942_out0;
wire  [15:0] v$NEXTENDED_14372_out0;
wire  [15:0] v$NEXTENDED_14373_out0;
wire  [15:0] v$NEXTENDED_1909_out0;
wire  [15:0] v$NEXTENDED_1910_out0;
wire  [15:0] v$OP1_15212_out0;
wire  [15:0] v$OP1_15213_out0;
wire  [15:0] v$OP1_5416_out0;
wire  [15:0] v$OP1_5417_out0;
wire  [15:0] v$OP2_10191_out0;
wire  [15:0] v$OP2_10192_out0;
wire  [15:0] v$OP2_13995_out0;
wire  [15:0] v$OP2_13996_out0;
wire  [15:0] v$OP2_15055_out0;
wire  [15:0] v$OP2_15056_out0;
wire  [15:0] v$OP2_7579_out0;
wire  [15:0] v$OP2_7580_out0;
wire  [15:0] v$OUT_12478_out0;
wire  [15:0] v$OUT_12480_out0;
wire  [15:0] v$OUT_1321_out0;
wire  [15:0] v$OUT_1322_out0;
wire  [15:0] v$OUT_14505_out0;
wire  [15:0] v$OUT_14506_out0;
wire  [15:0] v$OUT_3176_out0;
wire  [15:0] v$OUT_3177_out0;
wire  [15:0] v$OUT_3178_out0;
wire  [15:0] v$OUT_3179_out0;
wire  [15:0] v$OUT_3180_out0;
wire  [15:0] v$OUT_3181_out0;
wire  [15:0] v$OUT_3182_out0;
wire  [15:0] v$OUT_3183_out0;
wire  [15:0] v$OUT_5259_out0;
wire  [15:0] v$OUT_5260_out0;
wire  [15:0] v$PIN_2935_out0;
wire  [15:0] v$PIN_2936_out0;
wire  [15:0] v$R0TEST_14040_out0;
wire  [15:0] v$R0TEST_14041_out0;
wire  [15:0] v$R0TEST_8236_out0;
wire  [15:0] v$R0TEST_8237_out0;
wire  [15:0] v$R0_3278_out0;
wire  [15:0] v$R0_3279_out0;
wire  [15:0] v$R1TEST_15146_out0;
wire  [15:0] v$R1TEST_15147_out0;
wire  [15:0] v$R1TEST_8249_out0;
wire  [15:0] v$R1TEST_8250_out0;
wire  [15:0] v$R1_13766_out0;
wire  [15:0] v$R1_13767_out0;
wire  [15:0] v$R2TEST_15718_out0;
wire  [15:0] v$R2TEST_15719_out0;
wire  [15:0] v$R2TEST_15806_out0;
wire  [15:0] v$R2TEST_15807_out0;
wire  [15:0] v$R2_7958_out0;
wire  [15:0] v$R2_7959_out0;
wire  [15:0] v$R3TEST_11804_out0;
wire  [15:0] v$R3TEST_11805_out0;
wire  [15:0] v$R3TEST_7537_out0;
wire  [15:0] v$R3TEST_7538_out0;
wire  [15:0] v$R3_10746_out0;
wire  [15:0] v$R3_10747_out0;
wire  [15:0] v$RAM1_12913_out0;
wire  [15:0] v$RAMDIN_7038_out0;
wire  [15:0] v$RAMDIN_7039_out0;
wire  [15:0] v$RAMDOUT$DATAPATH_642_out0;
wire  [15:0] v$RAMDOUT$DATAPATH_643_out0;
wire  [15:0] v$RAMDOUT0_9099_out0;
wire  [15:0] v$RAMDOUT1_8315_out0;
wire  [15:0] v$RAMDOUT_16779_out0;
wire  [15:0] v$RAMDOUT_16780_out0;
wire  [15:0] v$RAMDOUT_5423_out0;
wire  [15:0] v$RAMDOUT_5424_out0;
wire  [15:0] v$RAMDOUT_68_out0;
wire  [15:0] v$RAMDOUT_69_out0;
wire  [15:0] v$RAMDOUT_7917_out0;
wire  [15:0] v$RAMDOUT_7918_out0;
wire  [15:0] v$RAMDOutOut_3187_out0;
wire  [15:0] v$RAMDOutOut_3188_out0;
wire  [15:0] v$RDOUT_10345_out0;
wire  [15:0] v$RDOUT_10346_out0;
wire  [15:0] v$RD_2226_out0;
wire  [15:0] v$RD_2227_out0;
wire  [15:0] v$REGDIN_16498_out0;
wire  [15:0] v$REGDIN_16499_out0;
wire  [15:0] v$REGDIN_18379_out0;
wire  [15:0] v$REGDIN_18380_out0;
wire  [15:0] v$RMN_6155_out0;
wire  [15:0] v$RMN_6156_out0;
wire  [15:0] v$RMORIGINAL_12978_out0;
wire  [15:0] v$RMORIGINAL_12979_out0;
wire  [15:0] v$RM_10242_out0;
wire  [15:0] v$RM_10243_out0;
wire  [15:0] v$RM_16193_out0;
wire  [15:0] v$RM_16194_out0;
wire  [15:0] v$RM_18197_out0;
wire  [15:0] v$RM_18198_out0;
wire  [15:0] v$RM_18596_out0;
wire  [15:0] v$RM_18597_out0;
wire  [15:0] v$RM_9426_out0;
wire  [15:0] v$RM_9427_out0;
wire  [15:0] v$ROM1_17450_out0;
wire  [15:0] v$ROM1_17451_out0;
wire  [15:0] v$R_18353_out0;
wire  [15:0] v$R_18354_out0;
wire  [15:0] v$R_59_out0;
wire  [15:0] v$R_60_out0;
wire  [15:0] v$SEL11_3703_out0;
wire  [15:0] v$SEL12_1192_out0;
wire  [15:0] v$SEL1_15387_out0;
wire  [15:0] v$SEL1_15392_out0;
wire  [15:0] v$SEL1_15397_out0;
wire  [15:0] v$SEL1_15402_out0;
wire  [15:0] v$SEL1_15407_out0;
wire  [15:0] v$SEL1_15412_out0;
wire  [15:0] v$SEL1_15418_out0;
wire  [15:0] v$SEL1_15422_out0;
wire  [15:0] v$SEL1_15428_out0;
wire  [15:0] v$SEL1_15435_out0;
wire  [15:0] v$SEL1_15440_out0;
wire  [15:0] v$SEL1_15445_out0;
wire  [15:0] v$SEL1_16688_out0;
wire  [15:0] v$SEL1_16692_out0;
wire  [15:0] v$SEL1_8696_out0;
wire  [15:0] v$SEL1_8701_out0;
wire  [15:0] v$SEL1_8706_out0;
wire  [15:0] v$SEL1_8711_out0;
wire  [15:0] v$SEL1_8716_out0;
wire  [15:0] v$SEL1_8721_out0;
wire  [15:0] v$SEL1_8727_out0;
wire  [15:0] v$SEL1_8731_out0;
wire  [15:0] v$SEL1_8737_out0;
wire  [15:0] v$SEL1_8744_out0;
wire  [15:0] v$SEL1_8749_out0;
wire  [15:0] v$SEL1_8754_out0;
wire  [15:0] v$SEL2_13852_out0;
wire  [15:0] v$SEL2_13856_out0;
wire  [15:0] v$SEL2_6393_out0;
wire  [15:0] v$SEL2_6394_out0;
wire  [15:0] v$SEL3_7366_out0;
wire  [15:0] v$SEL3_7370_out0;
wire  [15:0] v$SEL4_9556_out0;
wire  [15:0] v$SEL4_9557_out0;
wire  [15:0] v$SEL5_13590_out0;
wire  [15:0] v$SEL5_13591_out0;
wire  [15:0] v$SHIFT1OUT_7581_out0;
wire  [15:0] v$SHIFT1OUT_7582_out0;
wire  [15:0] v$SHIFT2OUT_15679_out0;
wire  [15:0] v$SHIFT2OUT_15680_out0;
wire  [15:0] v$SHIFT4OUT_5942_out0;
wire  [15:0] v$SHIFT4OUT_5943_out0;
wire  [15:0] v$SHIFT8OUT_8011_out0;
wire  [15:0] v$SHIFT8OUT_8012_out0;
wire  [15:0] v$SUM_10304_out0;
wire  [15:0] v$SUM_10305_out0;
wire  [15:0] v$THRESHOLD_15533_out0;
wire  [15:0] v$THRESHOLD_15534_out0;
wire  [15:0] v$UART$DOUT_17461_out0;
wire  [15:0] v$UART$DOUT_17462_out0;
wire  [15:0] v$XOR1_5078_out0;
wire  [15:0] v$XOR1_5079_out0;
wire  [15:0] v$XOR1_9542_out0;
wire  [15:0] v$XOR1_9543_out0;
wire  [15:0] v$_11646_out0;
wire  [15:0] v$_11647_out0;
wire  [15:0] v$_11757_out0;
wire  [15:0] v$_11758_out0;
wire  [15:0] v$_11808_out0;
wire  [15:0] v$_11809_out0;
wire  [15:0] v$_11810_out0;
wire  [15:0] v$_11811_out0;
wire  [15:0] v$_11812_out0;
wire  [15:0] v$_11813_out0;
wire  [15:0] v$_11814_out0;
wire  [15:0] v$_11815_out0;
wire  [15:0] v$_12228_out0;
wire  [15:0] v$_12229_out0;
wire  [15:0] v$_13304_out0;
wire  [15:0] v$_13305_out0;
wire  [15:0] v$_13306_out0;
wire  [15:0] v$_13307_out0;
wire  [15:0] v$_13308_out0;
wire  [15:0] v$_13309_out0;
wire  [15:0] v$_13310_out0;
wire  [15:0] v$_13311_out0;
wire  [15:0] v$_1477_out0;
wire  [15:0] v$_1478_out0;
wire  [15:0] v$_1479_out0;
wire  [15:0] v$_1480_out0;
wire  [15:0] v$_1481_out0;
wire  [15:0] v$_1482_out0;
wire  [15:0] v$_1483_out0;
wire  [15:0] v$_1484_out0;
wire  [15:0] v$_1494_out0;
wire  [15:0] v$_1495_out0;
wire  [15:0] v$_16367_out1;
wire  [15:0] v$_16368_out1;
wire  [15:0] v$_16369_out0;
wire  [15:0] v$_16370_out0;
wire  [15:0] v$_17478_out0;
wire  [15:0] v$_17479_out0;
wire  [15:0] v$_18233_out0;
wire  [15:0] v$_18234_out0;
wire  [15:0] v$_18235_out0;
wire  [15:0] v$_18236_out0;
wire  [15:0] v$_18237_out0;
wire  [15:0] v$_18416_out0;
wire  [15:0] v$_18418_out0;
wire  [15:0] v$_4867_out0;
wire  [15:0] v$_4868_out0;
wire  [15:0] v$_4869_out0;
wire  [15:0] v$_4870_out0;
wire  [15:0] v$_4871_out0;
wire  [15:0] v$_6913_out0;
wire  [15:0] v$_6914_out0;
wire  [15:0] v$_9445_out0;
wire  [15:0] v$_9446_out0;
wire  [15:0] v$_9447_out0;
wire  [15:0] v$_9448_out0;
wire  [15:0] v$_9449_out0;
wire  [15:0] v$_9450_out0;
wire  [15:0] v$_9451_out0;
wire  [15:0] v$_9452_out0;
wire  [15:0] v$_9931_out1;
wire  [15:0] v$_9932_out1;
wire  [19:0] v$SEL1_15389_out0;
wire  [19:0] v$SEL1_15394_out0;
wire  [19:0] v$SEL1_15399_out0;
wire  [19:0] v$SEL1_15403_out0;
wire  [19:0] v$SEL1_15409_out0;
wire  [19:0] v$SEL1_15413_out0;
wire  [19:0] v$SEL1_15420_out0;
wire  [19:0] v$SEL1_15437_out0;
wire  [19:0] v$SEL1_15442_out0;
wire  [19:0] v$SEL1_15447_out0;
wire  [19:0] v$SEL1_8698_out0;
wire  [19:0] v$SEL1_8703_out0;
wire  [19:0] v$SEL1_8708_out0;
wire  [19:0] v$SEL1_8712_out0;
wire  [19:0] v$SEL1_8718_out0;
wire  [19:0] v$SEL1_8722_out0;
wire  [19:0] v$SEL1_8729_out0;
wire  [19:0] v$SEL1_8746_out0;
wire  [19:0] v$SEL1_8751_out0;
wire  [19:0] v$SEL1_8756_out0;
wire  [1:0] v$2_12738_out0;
wire  [1:0] v$2_12739_out0;
wire  [1:0] v$5_7508_out0;
wire  [1:0] v$5_7509_out0;
wire  [1:0] v$7_14010_out0;
wire  [1:0] v$7_14011_out0;
wire  [1:0] v$8_1193_out0;
wire  [1:0] v$8_1194_out0;
wire  [1:0] v$AD1VIEWER_7010_out0;
wire  [1:0] v$AD1VIEWER_7011_out0;
wire  [1:0] v$AD1_1840_out0;
wire  [1:0] v$AD1_1841_out0;
wire  [1:0] v$AD1_18672_out0;
wire  [1:0] v$AD1_18673_out0;
wire  [1:0] v$AD1_6656_out0;
wire  [1:0] v$AD1_6657_out0;
wire  [1:0] v$AD1_7604_out0;
wire  [1:0] v$AD1_7605_out0;
wire  [1:0] v$AD2$viewer_15750_out0;
wire  [1:0] v$AD2$viewer_15751_out0;
wire  [1:0] v$AD2_15661_out0;
wire  [1:0] v$AD2_15662_out0;
wire  [1:0] v$AD2_3939_out0;
wire  [1:0] v$AD2_3940_out0;
wire  [1:0] v$AD2_6401_out0;
wire  [1:0] v$AD2_6402_out0;
wire  [1:0] v$AD2_9095_out0;
wire  [1:0] v$AD2_9096_out0;
wire  [1:0] v$AD3$VIEWER_8318_out0;
wire  [1:0] v$AD3$VIEWER_8319_out0;
wire  [1:0] v$AD3_13143_out0;
wire  [1:0] v$AD3_13144_out0;
wire  [1:0] v$AD3_15144_out0;
wire  [1:0] v$AD3_15145_out0;
wire  [1:0] v$C1_14253_out0;
wire  [1:0] v$C1_14254_out0;
wire  [1:0] v$C1_3018_out0;
wire  [1:0] v$C1_3019_out0;
wire  [1:0] v$C1_5965_out0;
wire  [1:0] v$C1_5970_out0;
wire  [1:0] v$C1_5975_out0;
wire  [1:0] v$C1_5980_out0;
wire  [1:0] v$C1_5985_out0;
wire  [1:0] v$C1_5990_out0;
wire  [1:0] v$C1_5996_out0;
wire  [1:0] v$C1_5999_out0;
wire  [1:0] v$C1_6005_out0;
wire  [1:0] v$C1_6013_out0;
wire  [1:0] v$C1_6018_out0;
wire  [1:0] v$C1_6023_out0;
wire  [1:0] v$C1_7724_out0;
wire  [1:0] v$C1_7725_out0;
wire  [1:0] v$C1_7972_out0;
wire  [1:0] v$C1_7976_out0;
wire  [1:0] v$C2_107_out0;
wire  [1:0] v$C2_112_out0;
wire  [1:0] v$C2_117_out0;
wire  [1:0] v$C2_122_out0;
wire  [1:0] v$C2_127_out0;
wire  [1:0] v$C2_132_out0;
wire  [1:0] v$C2_13386_out0;
wire  [1:0] v$C2_13387_out0;
wire  [1:0] v$C2_138_out0;
wire  [1:0] v$C2_141_out0;
wire  [1:0] v$C2_147_out0;
wire  [1:0] v$C2_155_out0;
wire  [1:0] v$C2_160_out0;
wire  [1:0] v$C2_165_out0;
wire  [1:0] v$C3_3302_out0;
wire  [1:0] v$C3_3303_out0;
wire  [1:0] v$C3_3304_out0;
wire  [1:0] v$C3_3305_out0;
wire  [1:0] v$C3_3306_out0;
wire  [1:0] v$C3_3307_out0;
wire  [1:0] v$C3_3308_out0;
wire  [1:0] v$C3_3309_out0;
wire  [1:0] v$C4_16302_out0;
wire  [1:0] v$C4_16303_out0;
wire  [1:0] v$C4_16509_out0;
wire  [1:0] v$C4_16510_out0;
wire  [1:0] v$C4_16511_out0;
wire  [1:0] v$C4_16512_out0;
wire  [1:0] v$C4_16513_out0;
wire  [1:0] v$C4_16514_out0;
wire  [1:0] v$C4_16515_out0;
wire  [1:0] v$C4_16516_out0;
wire  [1:0] v$C4_16517_out0;
wire  [1:0] v$C4_16518_out0;
wire  [1:0] v$C5_16909_out0;
wire  [1:0] v$C5_16911_out0;
wire  [1:0] v$C5_16912_out0;
wire  [1:0] v$C5_16913_out0;
wire  [1:0] v$C5_16914_out0;
wire  [1:0] v$C5_16915_out0;
wire  [1:0] v$C5_16916_out0;
wire  [1:0] v$C5_16917_out0;
wire  [1:0] v$C5_16918_out0;
wire  [1:0] v$C5_16919_out0;
wire  [1:0] v$C6_6534_out0;
wire  [1:0] v$C6_6535_out0;
wire  [1:0] v$C6_6536_out0;
wire  [1:0] v$C6_6537_out0;
wire  [1:0] v$C6_6538_out0;
wire  [1:0] v$C6_6539_out0;
wire  [1:0] v$C6_6540_out0;
wire  [1:0] v$C6_6541_out0;
wire  [1:0] v$C6_6542_out0;
wire  [1:0] v$C6_6543_out0;
wire  [1:0] v$C6_6544_out0;
wire  [1:0] v$C6_6545_out0;
wire  [1:0] v$END_388_out0;
wire  [1:0] v$END_389_out0;
wire  [1:0] v$FPU$OP_12762_out0;
wire  [1:0] v$FPU$OP_12763_out0;
wire  [1:0] v$FPU$OP_14068_out0;
wire  [1:0] v$FPU$OP_14069_out0;
wire  [1:0] v$FPU$OP_15736_out0;
wire  [1:0] v$FPU$OP_15737_out0;
wire  [1:0] v$INTERRUPTNUMBER_39_out0;
wire  [1:0] v$INTERRUPTNUMBER_40_out0;
wire  [1:0] v$IR1$D_14847_out0;
wire  [1:0] v$IR1$D_14848_out0;
wire  [1:0] v$IR1$D_4219_out0;
wire  [1:0] v$IR1$D_4220_out0;
wire  [1:0] v$IR1$FPU$OP$CODE_18316_out0;
wire  [1:0] v$IR1$FPU$OP$CODE_18317_out0;
wire  [1:0] v$IR1$FPU$OP_3837_out0;
wire  [1:0] v$IR1$FPU$OP_3838_out0;
wire  [1:0] v$IR1$M_12632_out0;
wire  [1:0] v$IR1$M_12633_out0;
wire  [1:0] v$IR1$M_13247_out0;
wire  [1:0] v$IR1$M_13248_out0;
wire  [1:0] v$IR1$RD$VIEWER_18371_out0;
wire  [1:0] v$IR1$RD$VIEWER_18372_out0;
wire  [1:0] v$IR1$RD_5489_out0;
wire  [1:0] v$IR1$RD_5490_out0;
wire  [1:0] v$IR1$RM$VIEWER_7910_out0;
wire  [1:0] v$IR1$RM$VIEWER_7911_out0;
wire  [1:0] v$IR1$RM_18301_out0;
wire  [1:0] v$IR1$RM_18302_out0;
wire  [1:0] v$IR1$RM_18_out0;
wire  [1:0] v$IR1$RM_19_out0;
wire  [1:0] v$IR2$D_14491_out0;
wire  [1:0] v$IR2$D_14492_out0;
wire  [1:0] v$IR2$D_4898_out0;
wire  [1:0] v$IR2$D_4899_out0;
wire  [1:0] v$IR2$FPU$OP_1687_out0;
wire  [1:0] v$IR2$FPU$OP_1688_out0;
wire  [1:0] v$IR2$FPU$OP_2881_out0;
wire  [1:0] v$IR2$FPU$OP_2882_out0;
wire  [1:0] v$IR2$FPU$OP_7546_out0;
wire  [1:0] v$IR2$FPU$OP_7547_out0;
wire  [1:0] v$IR2$M_12993_out0;
wire  [1:0] v$IR2$M_12994_out0;
wire  [1:0] v$IR2$M_8832_out0;
wire  [1:0] v$IR2$M_8833_out0;
wire  [1:0] v$IR2$RD$VIEWER_9124_out0;
wire  [1:0] v$IR2$RD$VIEWER_9125_out0;
wire  [1:0] v$IR2$RD_13291_out0;
wire  [1:0] v$IR2$RD_13292_out0;
wire  [1:0] v$IR2$RD_16358_out0;
wire  [1:0] v$IR2$RD_16359_out0;
wire  [1:0] v$MUX10_3626_out0;
wire  [1:0] v$MUX10_3627_out0;
wire  [1:0] v$MUX11_4487_out0;
wire  [1:0] v$MUX11_4488_out0;
wire  [1:0] v$MUX16_8689_out0;
wire  [1:0] v$MUX1_8336_out0;
wire  [1:0] v$MUX1_8337_out0;
wire  [1:0] v$MUX2_2884_out0;
wire  [1:0] v$MUX2_2885_out0;
wire  [1:0] v$MUX5_7954_out0;
wire  [1:0] v$MUX5_7955_out0;
wire  [1:0] v$MUX6_1311_out0;
wire  [1:0] v$MUX6_1312_out0;
wire  [1:0] v$MUX9_7648_out0;
wire  [1:0] v$MUX9_7649_out0;
wire  [1:0] v$NINTERRUPT_1595_out0;
wire  [1:0] v$NINTERRUPT_1596_out0;
wire  [1:0] v$NINT_2845_out0;
wire  [1:0] v$NINT_2846_out0;
wire  [1:0] v$OP_1323_out0;
wire  [1:0] v$OP_1324_out0;
wire  [1:0] v$RD$FPU_12947_out0;
wire  [1:0] v$RD$OUT_17889_out0;
wire  [1:0] v$RD_11793_out0;
wire  [1:0] v$S$REG_3443_out0;
wire  [1:0] v$S$REG_3444_out0;
wire  [1:0] v$SEL10_12823_out0;
wire  [1:0] v$SEL10_12824_out0;
wire  [1:0] v$SEL13_4841_out0;
wire  [1:0] v$SEL13_4842_out0;
wire  [1:0] v$SEL1_5240_out0;
wire  [1:0] v$SEL1_5241_out0;
wire  [1:0] v$SEL4_9443_out0;
wire  [1:0] v$SEL4_9444_out0;
wire  [1:0] v$SEL5_644_out0;
wire  [1:0] v$SEL5_645_out0;
wire  [1:0] v$SEL6_3008_out0;
wire  [1:0] v$SEL6_3009_out0;
wire  [1:0] v$SEL8_15116_out0;
wire  [1:0] v$SEL8_15117_out0;
wire  [1:0] v$SEL9_7983_out0;
wire  [1:0] v$SEL9_7984_out0;
wire  [1:0] v$SHIFT_7019_out0;
wire  [1:0] v$SHIFT_7020_out0;
wire  [1:0] v$SHIFT_8028_out0;
wire  [1:0] v$SHIFT_8029_out0;
wire  [1:0] v$SR_16801_out0;
wire  [1:0] v$SR_16802_out0;
wire  [1:0] v$SR_16803_out0;
wire  [1:0] v$SR_16804_out0;
wire  [1:0] v$SR_16805_out0;
wire  [1:0] v$SR_16806_out0;
wire  [1:0] v$SR_16807_out0;
wire  [1:0] v$SR_16808_out0;
wire  [1:0] v$SR_4368_out0;
wire  [1:0] v$SR_4369_out0;
wire  [1:0] v$SR_4370_out0;
wire  [1:0] v$SR_4371_out0;
wire  [1:0] v$SR_4372_out0;
wire  [1:0] v$SR_4373_out0;
wire  [1:0] v$SR_4374_out0;
wire  [1:0] v$SR_4375_out0;
wire  [1:0] v$SR_9927_out0;
wire  [1:0] v$SR_9928_out0;
wire  [1:0] v$XOR1_5009_out0;
wire  [1:0] v$XOR1_5010_out0;
wire  [1:0] v$XOR1_8327_out0;
wire  [1:0] v$XOR1_8328_out0;
wire  [1:0] v$XOR2_18493_out0;
wire  [1:0] v$XOR2_18494_out0;
wire  [1:0] v$XOR3_4037_out0;
wire  [1:0] v$XOR3_4038_out0;
wire  [1:0] v$Y_6483_out0;
wire  [1:0] v$Y_6484_out0;
wire  [1:0] v$Y_6485_out0;
wire  [1:0] v$Y_6486_out0;
wire  [1:0] v$Y_6487_out0;
wire  [1:0] v$Y_6488_out0;
wire  [1:0] v$Y_6489_out0;
wire  [1:0] v$Y_6490_out0;
wire  [1:0] v$Y_6491_out0;
wire  [1:0] v$Y_6492_out0;
wire  [1:0] v$Y_6493_out0;
wire  [1:0] v$Y_6494_out0;
wire  [1:0] v$Y_6495_out0;
wire  [1:0] v$Y_6496_out0;
wire  [1:0] v$Y_6497_out0;
wire  [1:0] v$Y_6498_out0;
wire  [1:0] v$Y_6499_out0;
wire  [1:0] v$Y_6500_out0;
wire  [1:0] v$Y_6501_out0;
wire  [1:0] v$Y_6502_out0;
wire  [1:0] v$Y_6503_out0;
wire  [1:0] v$Y_6504_out0;
wire  [1:0] v$Y_6505_out0;
wire  [1:0] v$Y_6506_out0;
wire  [1:0] v$Y_6507_out0;
wire  [1:0] v$Y_6508_out0;
wire  [1:0] v$Y_6509_out0;
wire  [1:0] v$Y_6510_out0;
wire  [1:0] v$Y_6511_out0;
wire  [1:0] v$Y_6512_out0;
wire  [1:0] v$Y_6513_out0;
wire  [1:0] v$Y_6514_out0;
wire  [1:0] v$Y_6515_out0;
wire  [1:0] v$Y_6516_out0;
wire  [1:0] v$Y_6517_out0;
wire  [1:0] v$Y_6518_out0;
wire  [1:0] v$Y_6519_out0;
wire  [1:0] v$Y_6520_out0;
wire  [1:0] v$Y_6521_out0;
wire  [1:0] v$Y_6522_out0;
wire  [1:0] v$Y_6523_out0;
wire  [1:0] v$Y_6524_out0;
wire  [1:0] v$Y_6525_out0;
wire  [1:0] v$Y_6526_out0;
wire  [1:0] v$Y_6527_out0;
wire  [1:0] v$Y_6528_out0;
wire  [1:0] v$Y_6529_out0;
wire  [1:0] v$Y_6530_out0;
wire  [1:0] v$_10237_out0;
wire  [1:0] v$_10238_out0;
wire  [1:0] v$_10239_out0;
wire  [1:0] v$_10240_out0;
wire  [1:0] v$_10241_out0;
wire  [1:0] v$_10446_out1;
wire  [1:0] v$_10447_out1;
wire  [1:0] v$_10448_out1;
wire  [1:0] v$_10449_out1;
wire  [1:0] v$_10450_out1;
wire  [1:0] v$_10772_out1;
wire  [1:0] v$_10773_out1;
wire  [1:0] v$_10774_out1;
wire  [1:0] v$_10775_out1;
wire  [1:0] v$_10776_out1;
wire  [1:0] v$_10791_out0;
wire  [1:0] v$_10792_out0;
wire  [1:0] v$_10810_out0;
wire  [1:0] v$_10810_out1;
wire  [1:0] v$_10811_out0;
wire  [1:0] v$_10811_out1;
wire  [1:0] v$_10910_out1;
wire  [1:0] v$_10911_out1;
wire  [1:0] v$_10912_out1;
wire  [1:0] v$_10913_out1;
wire  [1:0] v$_10914_out1;
wire  [1:0] v$_10958_out0;
wire  [1:0] v$_10959_out0;
wire  [1:0] v$_10960_out0;
wire  [1:0] v$_10961_out0;
wire  [1:0] v$_10962_out0;
wire  [1:0] v$_10974_out0;
wire  [1:0] v$_10975_out0;
wire  [1:0] v$_11099_out1;
wire  [1:0] v$_11100_out1;
wire  [1:0] v$_11101_out1;
wire  [1:0] v$_11102_out1;
wire  [1:0] v$_11103_out1;
wire  [1:0] v$_11816_out0;
wire  [1:0] v$_11816_out1;
wire  [1:0] v$_11817_out0;
wire  [1:0] v$_11817_out1;
wire  [1:0] v$_1199_out0;
wire  [1:0] v$_1200_out0;
wire  [1:0] v$_1201_out0;
wire  [1:0] v$_1202_out0;
wire  [1:0] v$_1203_out0;
wire  [1:0] v$_1273_out0;
wire  [1:0] v$_1274_out0;
wire  [1:0] v$_12840_out0;
wire  [1:0] v$_12840_out1;
wire  [1:0] v$_12841_out0;
wire  [1:0] v$_12841_out1;
wire  [1:0] v$_12842_out0;
wire  [1:0] v$_12842_out1;
wire  [1:0] v$_12843_out0;
wire  [1:0] v$_12843_out1;
wire  [1:0] v$_12844_out0;
wire  [1:0] v$_12844_out1;
wire  [1:0] v$_12845_out0;
wire  [1:0] v$_12845_out1;
wire  [1:0] v$_12846_out0;
wire  [1:0] v$_12846_out1;
wire  [1:0] v$_12847_out0;
wire  [1:0] v$_12847_out1;
wire  [1:0] v$_12848_out0;
wire  [1:0] v$_12848_out1;
wire  [1:0] v$_12849_out0;
wire  [1:0] v$_12849_out1;
wire  [1:0] v$_12850_out0;
wire  [1:0] v$_12850_out1;
wire  [1:0] v$_12851_out0;
wire  [1:0] v$_12851_out1;
wire  [1:0] v$_1302_out1;
wire  [1:0] v$_1303_out1;
wire  [1:0] v$_1304_out1;
wire  [1:0] v$_1305_out1;
wire  [1:0] v$_13065_out0;
wire  [1:0] v$_13066_out0;
wire  [1:0] v$_1306_out1;
wire  [1:0] v$_13151_out0;
wire  [1:0] v$_13151_out1;
wire  [1:0] v$_13152_out0;
wire  [1:0] v$_13152_out1;
wire  [1:0] v$_13221_out0;
wire  [1:0] v$_13222_out0;
wire  [1:0] v$_13256_out0;
wire  [1:0] v$_13256_out1;
wire  [1:0] v$_13257_out0;
wire  [1:0] v$_13257_out1;
wire  [1:0] v$_13283_out0;
wire  [1:0] v$_13283_out1;
wire  [1:0] v$_13284_out0;
wire  [1:0] v$_13284_out1;
wire  [1:0] v$_13289_out1;
wire  [1:0] v$_13290_out1;
wire  [1:0] v$_13293_out0;
wire  [1:0] v$_13294_out0;
wire  [1:0] v$_13295_out0;
wire  [1:0] v$_13296_out0;
wire  [1:0] v$_13297_out0;
wire  [1:0] v$_13410_out0;
wire  [1:0] v$_13411_out0;
wire  [1:0] v$_13437_out0;
wire  [1:0] v$_13438_out0;
wire  [1:0] v$_13439_out0;
wire  [1:0] v$_13440_out0;
wire  [1:0] v$_13441_out0;
wire  [1:0] v$_1353_out1;
wire  [1:0] v$_1354_out1;
wire  [1:0] v$_1355_out1;
wire  [1:0] v$_1356_out1;
wire  [1:0] v$_1357_out1;
wire  [1:0] v$_14164_out0;
wire  [1:0] v$_14165_out0;
wire  [1:0] v$_14166_out0;
wire  [1:0] v$_14167_out0;
wire  [1:0] v$_14212_out0;
wire  [1:0] v$_14213_out0;
wire  [1:0] v$_14612_out0;
wire  [1:0] v$_14613_out0;
wire  [1:0] v$_1473_out0;
wire  [1:0] v$_1473_out1;
wire  [1:0] v$_1474_out0;
wire  [1:0] v$_1474_out1;
wire  [1:0] v$_14774_out0;
wire  [1:0] v$_14775_out0;
wire  [1:0] v$_14836_out0;
wire  [1:0] v$_14837_out0;
wire  [1:0] v$_14838_out0;
wire  [1:0] v$_14839_out0;
wire  [1:0] v$_14840_out0;
wire  [1:0] v$_14895_out0;
wire  [1:0] v$_14896_out0;
wire  [1:0] v$_14998_out0;
wire  [1:0] v$_14999_out0;
wire  [1:0] v$_15000_out0;
wire  [1:0] v$_15001_out0;
wire  [1:0] v$_15002_out0;
wire  [1:0] v$_15013_out0;
wire  [1:0] v$_15014_out0;
wire  [1:0] v$_15015_out0;
wire  [1:0] v$_15016_out0;
wire  [1:0] v$_15017_out0;
wire  [1:0] v$_15018_out0;
wire  [1:0] v$_15018_out1;
wire  [1:0] v$_15019_out0;
wire  [1:0] v$_15019_out1;
wire  [1:0] v$_15148_out1;
wire  [1:0] v$_15149_out1;
wire  [1:0] v$_15150_out1;
wire  [1:0] v$_15151_out1;
wire  [1:0] v$_15152_out1;
wire  [1:0] v$_15298_out0;
wire  [1:0] v$_15299_out0;
wire  [1:0] v$_15708_out0;
wire  [1:0] v$_15709_out0;
wire  [1:0] v$_15710_out0;
wire  [1:0] v$_15711_out0;
wire  [1:0] v$_15712_out0;
wire  [1:0] v$_1576_out0;
wire  [1:0] v$_1577_out0;
wire  [1:0] v$_1578_out0;
wire  [1:0] v$_1579_out0;
wire  [1:0] v$_1580_out0;
wire  [1:0] v$_15923_out0;
wire  [1:0] v$_15924_out0;
wire  [1:0] v$_15954_out0;
wire  [1:0] v$_15955_out0;
wire  [1:0] v$_16000_out0;
wire  [1:0] v$_16001_out0;
wire  [1:0] v$_1604_out0;
wire  [1:0] v$_1604_out1;
wire  [1:0] v$_1605_out0;
wire  [1:0] v$_1605_out1;
wire  [1:0] v$_16130_out1;
wire  [1:0] v$_16131_out1;
wire  [1:0] v$_16132_out1;
wire  [1:0] v$_16133_out1;
wire  [1:0] v$_16134_out1;
wire  [1:0] v$_16135_out0;
wire  [1:0] v$_16136_out0;
wire  [1:0] v$_16231_out0;
wire  [1:0] v$_16231_out1;
wire  [1:0] v$_16232_out0;
wire  [1:0] v$_16232_out1;
wire  [1:0] v$_16265_out1;
wire  [1:0] v$_16266_out1;
wire  [1:0] v$_16267_out1;
wire  [1:0] v$_16268_out1;
wire  [1:0] v$_16269_out1;
wire  [1:0] v$_16310_out0;
wire  [1:0] v$_16311_out0;
wire  [1:0] v$_16312_out0;
wire  [1:0] v$_16313_out0;
wire  [1:0] v$_16314_out0;
wire  [1:0] v$_16737_out0;
wire  [1:0] v$_16738_out0;
wire  [1:0] v$_16740_out1;
wire  [1:0] v$_16741_out1;
wire  [1:0] v$_16742_out1;
wire  [1:0] v$_16743_out1;
wire  [1:0] v$_16744_out1;
wire  [1:0] v$_16775_out0;
wire  [1:0] v$_16776_out0;
wire  [1:0] v$_1696_out0;
wire  [1:0] v$_1696_out1;
wire  [1:0] v$_1697_out0;
wire  [1:0] v$_1697_out1;
wire  [1:0] v$_17057_out0;
wire  [1:0] v$_17058_out0;
wire  [1:0] v$_17456_out0;
wire  [1:0] v$_17457_out0;
wire  [1:0] v$_17458_out0;
wire  [1:0] v$_17459_out0;
wire  [1:0] v$_17460_out0;
wire  [1:0] v$_1793_out0;
wire  [1:0] v$_1794_out0;
wire  [1:0] v$_1795_out0;
wire  [1:0] v$_17969_out0;
wire  [1:0] v$_1796_out0;
wire  [1:0] v$_17970_out0;
wire  [1:0] v$_1797_out0;
wire  [1:0] v$_18188_out1;
wire  [1:0] v$_18189_out1;
wire  [1:0] v$_18190_out1;
wire  [1:0] v$_18191_out1;
wire  [1:0] v$_18192_out1;
wire  [1:0] v$_18297_out1;
wire  [1:0] v$_18298_out1;
wire  [1:0] v$_1829_out0;
wire  [1:0] v$_1830_out0;
wire  [1:0] v$_18326_out0;
wire  [1:0] v$_18327_out0;
wire  [1:0] v$_18410_out0;
wire  [1:0] v$_18411_out0;
wire  [1:0] v$_18518_out0;
wire  [1:0] v$_18519_out0;
wire  [1:0] v$_1854_out1;
wire  [1:0] v$_1855_out1;
wire  [1:0] v$_18565_out0;
wire  [1:0] v$_18566_out0;
wire  [1:0] v$_1856_out1;
wire  [1:0] v$_1857_out1;
wire  [1:0] v$_1858_out1;
wire  [1:0] v$_18664_out0;
wire  [1:0] v$_18665_out0;
wire  [1:0] v$_18666_out0;
wire  [1:0] v$_18667_out0;
wire  [1:0] v$_18668_out0;
wire  [1:0] v$_212_out0;
wire  [1:0] v$_212_out1;
wire  [1:0] v$_213_out0;
wire  [1:0] v$_213_out1;
wire  [1:0] v$_2264_out0;
wire  [1:0] v$_2265_out0;
wire  [1:0] v$_2289_out0;
wire  [1:0] v$_2289_out1;
wire  [1:0] v$_2290_out0;
wire  [1:0] v$_2290_out1;
wire  [1:0] v$_229_out0;
wire  [1:0] v$_229_out1;
wire  [1:0] v$_230_out0;
wire  [1:0] v$_230_out1;
wire  [1:0] v$_2453_out0;
wire  [1:0] v$_2454_out0;
wire  [1:0] v$_2455_out0;
wire  [1:0] v$_2456_out0;
wire  [1:0] v$_2457_out0;
wire  [1:0] v$_2669_out0;
wire  [1:0] v$_2670_out0;
wire  [1:0] v$_2840_out0;
wire  [1:0] v$_2841_out0;
wire  [1:0] v$_2842_out0;
wire  [1:0] v$_2843_out0;
wire  [1:0] v$_2844_out0;
wire  [1:0] v$_2922_out1;
wire  [1:0] v$_2923_out1;
wire  [1:0] v$_2924_out1;
wire  [1:0] v$_2925_out1;
wire  [1:0] v$_2926_out1;
wire  [1:0] v$_3145_out0;
wire  [1:0] v$_3146_out0;
wire  [1:0] v$_3636_out0;
wire  [1:0] v$_3637_out0;
wire  [1:0] v$_3638_out0;
wire  [1:0] v$_3639_out0;
wire  [1:0] v$_3640_out0;
wire  [1:0] v$_3701_out0;
wire  [1:0] v$_3701_out1;
wire  [1:0] v$_3702_out0;
wire  [1:0] v$_3702_out1;
wire  [1:0] v$_3785_out0;
wire  [1:0] v$_3786_out0;
wire  [1:0] v$_5082_out0;
wire  [1:0] v$_5083_out0;
wire  [1:0] v$_5142_out0;
wire  [1:0] v$_5142_out1;
wire  [1:0] v$_5143_out0;
wire  [1:0] v$_5143_out1;
wire  [1:0] v$_54_out0;
wire  [1:0] v$_54_out1;
wire  [1:0] v$_55_out0;
wire  [1:0] v$_55_out1;
wire  [1:0] v$_5896_out0;
wire  [1:0] v$_5897_out0;
wire  [1:0] v$_5898_out0;
wire  [1:0] v$_5899_out0;
wire  [1:0] v$_5900_out0;
wire  [1:0] v$_6075_out1;
wire  [1:0] v$_6076_out1;
wire  [1:0] v$_6182_out0;
wire  [1:0] v$_6183_out0;
wire  [1:0] v$_6266_out0;
wire  [1:0] v$_6267_out0;
wire  [1:0] v$_6268_out0;
wire  [1:0] v$_6269_out0;
wire  [1:0] v$_6270_out0;
wire  [1:0] v$_6271_out0;
wire  [1:0] v$_6272_out0;
wire  [1:0] v$_6273_out0;
wire  [1:0] v$_6274_out0;
wire  [1:0] v$_6275_out0;
wire  [1:0] v$_6276_out0;
wire  [1:0] v$_6277_out0;
wire  [1:0] v$_6278_out0;
wire  [1:0] v$_6279_out0;
wire  [1:0] v$_6280_out0;
wire  [1:0] v$_6281_out0;
wire  [1:0] v$_6282_out0;
wire  [1:0] v$_6283_out0;
wire  [1:0] v$_6284_out0;
wire  [1:0] v$_6285_out0;
wire  [1:0] v$_6286_out0;
wire  [1:0] v$_6287_out0;
wire  [1:0] v$_6288_out0;
wire  [1:0] v$_6289_out0;
wire  [1:0] v$_6290_out0;
wire  [1:0] v$_6291_out0;
wire  [1:0] v$_6292_out0;
wire  [1:0] v$_6293_out0;
wire  [1:0] v$_6294_out0;
wire  [1:0] v$_6295_out0;
wire  [1:0] v$_6296_out0;
wire  [1:0] v$_6297_out0;
wire  [1:0] v$_6298_out0;
wire  [1:0] v$_6299_out0;
wire  [1:0] v$_6300_out0;
wire  [1:0] v$_6301_out0;
wire  [1:0] v$_6302_out0;
wire  [1:0] v$_6303_out0;
wire  [1:0] v$_6304_out0;
wire  [1:0] v$_6305_out0;
wire  [1:0] v$_6306_out0;
wire  [1:0] v$_6307_out0;
wire  [1:0] v$_6308_out0;
wire  [1:0] v$_6309_out0;
wire  [1:0] v$_6310_out0;
wire  [1:0] v$_6311_out0;
wire  [1:0] v$_6312_out0;
wire  [1:0] v$_6313_out0;
wire  [1:0] v$_650_out0;
wire  [1:0] v$_651_out0;
wire  [1:0] v$_652_out0;
wire  [1:0] v$_653_out0;
wire  [1:0] v$_654_out0;
wire  [1:0] v$_7067_out1;
wire  [1:0] v$_7068_out1;
wire  [1:0] v$_7069_out1;
wire  [1:0] v$_7070_out1;
wire  [1:0] v$_7071_out1;
wire  [1:0] v$_7374_out0;
wire  [1:0] v$_7374_out1;
wire  [1:0] v$_7375_out0;
wire  [1:0] v$_7375_out1;
wire  [1:0] v$_7467_out0;
wire  [1:0] v$_7467_out1;
wire  [1:0] v$_7468_out0;
wire  [1:0] v$_7468_out1;
wire  [1:0] v$_7552_out0;
wire  [1:0] v$_7553_out0;
wire  [1:0] v$_7554_out0;
wire  [1:0] v$_7555_out0;
wire  [1:0] v$_7556_out0;
wire  [1:0] v$_7734_out0;
wire  [1:0] v$_7735_out0;
wire  [1:0] v$_7768_out1;
wire  [1:0] v$_7769_out1;
wire  [1:0] v$_7770_out1;
wire  [1:0] v$_7771_out1;
wire  [1:0] v$_7772_out1;
wire  [1:0] v$_7868_out0;
wire  [1:0] v$_7869_out0;
wire  [1:0] v$_7870_out0;
wire  [1:0] v$_7871_out0;
wire  [1:0] v$_7872_out0;
wire  [1:0] v$_8208_out0;
wire  [1:0] v$_8208_out1;
wire  [1:0] v$_8209_out0;
wire  [1:0] v$_8209_out1;
wire  [1:0] v$_82_out0;
wire  [1:0] v$_8329_out0;
wire  [1:0] v$_8330_out0;
wire  [1:0] v$_8331_out0;
wire  [1:0] v$_8332_out0;
wire  [1:0] v$_8333_out0;
wire  [1:0] v$_83_out0;
wire  [1:0] v$_8452_out0;
wire  [1:0] v$_8452_out1;
wire  [1:0] v$_8453_out0;
wire  [1:0] v$_8453_out1;
wire  [1:0] v$_8454_out0;
wire  [1:0] v$_8454_out1;
wire  [1:0] v$_8455_out0;
wire  [1:0] v$_8455_out1;
wire  [1:0] v$_8456_out0;
wire  [1:0] v$_8456_out1;
wire  [1:0] v$_8457_out0;
wire  [1:0] v$_8457_out1;
wire  [1:0] v$_8458_out0;
wire  [1:0] v$_8458_out1;
wire  [1:0] v$_8459_out0;
wire  [1:0] v$_8459_out1;
wire  [1:0] v$_8460_out0;
wire  [1:0] v$_8460_out1;
wire  [1:0] v$_8461_out0;
wire  [1:0] v$_8461_out1;
wire  [1:0] v$_8462_out0;
wire  [1:0] v$_8462_out1;
wire  [1:0] v$_8463_out0;
wire  [1:0] v$_8463_out1;
wire  [1:0] v$_84_out0;
wire  [1:0] v$_85_out0;
wire  [1:0] v$_86_out0;
wire  [1:0] v$_8906_out0;
wire  [1:0] v$_8907_out0;
wire  [1:0] v$_8908_out0;
wire  [1:0] v$_8909_out0;
wire  [1:0] v$_8910_out0;
wire  [1:0] v$_9062_out1;
wire  [1:0] v$_9063_out1;
wire  [1:0] v$_9064_out1;
wire  [1:0] v$_9065_out1;
wire  [1:0] v$_9066_out1;
wire  [1:0] v$_909_out0;
wire  [1:0] v$_910_out0;
wire  [1:0] v$_9420_out0;
wire  [1:0] v$_9420_out1;
wire  [1:0] v$_9421_out0;
wire  [1:0] v$_9421_out1;
wire  [1:0] v$_9436_out0;
wire  [1:0] v$_9437_out0;
wire  [1:0] v$_9457_out0;
wire  [1:0] v$_9458_out0;
wire  [1:0] v$_9911_out0;
wire  [1:0] v$_9912_out0;
wire  [1:0] v$_9917_out0;
wire  [1:0] v$_9918_out0;
wire  [21:0] v$SEL1_15390_out0;
wire  [21:0] v$SEL1_15395_out0;
wire  [21:0] v$SEL1_15400_out0;
wire  [21:0] v$SEL1_15405_out0;
wire  [21:0] v$SEL1_15410_out0;
wire  [21:0] v$SEL1_15415_out0;
wire  [21:0] v$SEL1_15421_out0;
wire  [21:0] v$SEL1_15438_out0;
wire  [21:0] v$SEL1_15443_out0;
wire  [21:0] v$SEL1_15448_out0;
wire  [21:0] v$SEL1_8699_out0;
wire  [21:0] v$SEL1_8704_out0;
wire  [21:0] v$SEL1_8709_out0;
wire  [21:0] v$SEL1_8714_out0;
wire  [21:0] v$SEL1_8719_out0;
wire  [21:0] v$SEL1_8724_out0;
wire  [21:0] v$SEL1_8730_out0;
wire  [21:0] v$SEL1_8747_out0;
wire  [21:0] v$SEL1_8752_out0;
wire  [21:0] v$SEL1_8757_out0;
wire  [22:0] v$A$MANTISA$MUL_2654_out0;
wire  [22:0] v$A$MANTISA$MUL_2655_out0;
wire  [22:0] v$A$MANTISA_11825_out0;
wire  [22:0] v$A$MANTISA_11826_out0;
wire  [22:0] v$A$MANTISA_14549_out0;
wire  [22:0] v$A$MANTISA_14550_out0;
wire  [22:0] v$A$MANTISA_17915_out0;
wire  [22:0] v$A$MANTISA_17916_out0;
wire  [22:0] v$B$MANTISA$MUL_8165_out0;
wire  [22:0] v$B$MANTISA$MUL_8166_out0;
wire  [22:0] v$B$MANTISA_3002_out0;
wire  [22:0] v$B$MANTISA_3003_out0;
wire  [22:0] v$B$MANTISA_4070_out0;
wire  [22:0] v$B$MANTISA_4071_out0;
wire  [22:0] v$B$MANTISA_4908_out0;
wire  [22:0] v$B$MANTISA_4909_out0;
wire  [22:0] v$C5_15619_out0;
wire  [22:0] v$C5_15620_out0;
wire  [22:0] v$MANTISA$ADDITION_13173_out0;
wire  [22:0] v$MANTISA$ADDITION_13174_out0;
wire  [22:0] v$MANTISA$RESULT$BEFORE$MERGE_18716_out0;
wire  [22:0] v$MANTISA$RESULT$BEFORE$MERGE_18717_out0;
wire  [22:0] v$MANTISA$RESULT$FPU$ADDER_11900_out0;
wire  [22:0] v$MANTISA$RESULT$FPU$ADDER_11901_out0;
wire  [22:0] v$MANTISA$RESULT_6546_out0;
wire  [22:0] v$MANTISA$RESULT_6547_out0;
wire  [22:0] v$MUX1_1933_out0;
wire  [22:0] v$MUX1_1934_out0;
wire  [22:0] v$MUX2_1609_out0;
wire  [22:0] v$MUX2_1610_out0;
wire  [22:0] v$MUX2_2973_out0;
wire  [22:0] v$MUX2_2974_out0;
wire  [22:0] v$MUX6_12770_out0;
wire  [22:0] v$MUX6_12771_out0;
wire  [22:0] v$MUX7_12742_out0;
wire  [22:0] v$MUX7_12743_out0;
wire  [22:0] v$MUX8_7077_out0;
wire  [22:0] v$MUX8_7078_out0;
wire  [22:0] v$OUT1_10407_out0;
wire  [22:0] v$OUT1_10408_out0;
wire  [22:0] v$SEL1_14363_out0;
wire  [22:0] v$SEL1_14364_out0;
wire  [22:0] v$SEL1_15388_out0;
wire  [22:0] v$SEL1_15393_out0;
wire  [22:0] v$SEL1_15398_out0;
wire  [22:0] v$SEL1_15401_out0;
wire  [22:0] v$SEL1_15408_out0;
wire  [22:0] v$SEL1_15411_out0;
wire  [22:0] v$SEL1_15416_out0;
wire  [22:0] v$SEL1_15419_out0;
wire  [22:0] v$SEL1_15436_out0;
wire  [22:0] v$SEL1_15441_out0;
wire  [22:0] v$SEL1_15446_out0;
wire  [22:0] v$SEL1_15748_out0;
wire  [22:0] v$SEL1_15749_out0;
wire  [22:0] v$SEL1_6028_out0;
wire  [22:0] v$SEL1_8697_out0;
wire  [22:0] v$SEL1_8702_out0;
wire  [22:0] v$SEL1_8707_out0;
wire  [22:0] v$SEL1_8710_out0;
wire  [22:0] v$SEL1_8717_out0;
wire  [22:0] v$SEL1_8720_out0;
wire  [22:0] v$SEL1_8725_out0;
wire  [22:0] v$SEL1_8728_out0;
wire  [22:0] v$SEL1_8745_out0;
wire  [22:0] v$SEL1_8750_out0;
wire  [22:0] v$SEL1_8755_out0;
wire  [22:0] v$SEL2_11011_out0;
wire  [22:0] v$SEL2_11012_out0;
wire  [22:0] v$SEL2_6033_out0;
wire  [22:0] v$SEL2_6034_out0;
wire  [22:0] v$SEL2_8100_out0;
wire  [22:0] v$SEL3_11894_out0;
wire  [22:0] v$SEL3_11895_out0;
wire  [22:0] v$SEL3_14249_out0;
wire  [22:0] v$SEL3_14250_out0;
wire  [22:0] v$SEL4_12976_out0;
wire  [22:0] v$SEL4_12977_out0;
wire  [22:0] v$SEL4_2279_out0;
wire  [22:0] v$SEL4_2280_out0;
wire  [22:0] v$SEL4_7557_out0;
wire  [22:0] v$SEL5_10328_out0;
wire  [22:0] v$SEL6_4441_out0;
wire  [22:0] v$SEL6_4442_out0;
wire  [22:0] v$SEL8_17494_out0;
wire  [22:0] v$SEL8_17495_out0;
wire  [22:0] v$SEL8_17651_out0;
wire  [22:0] v$SEL8_17652_out0;
wire  [22:0] v$SEL8_17653_out0;
wire  [22:0] v$SEL8_17654_out0;
wire  [22:0] v$SEL8_17655_out0;
wire  [22:0] v$SEL8_17656_out0;
wire  [22:0] v$SEL8_17657_out0;
wire  [22:0] v$SEL8_17658_out0;
wire  [22:0] v$SEL8_17659_out0;
wire  [22:0] v$SEL8_17660_out0;
wire  [22:0] v$SEL8_17661_out0;
wire  [22:0] v$SEL8_17662_out0;
wire  [22:0] v$SEL8_7275_out0;
wire  [22:0] v$SEL8_7276_out0;
wire  [22:0] v$_16242_out0;
wire  [22:0] v$_16243_out0;
wire  [22:0] v$_1685_out0;
wire  [22:0] v$_1686_out0;
wire  [22:0] v$_18088_out0;
wire  [22:0] v$_18089_out0;
wire  [22:0] v$_2231_out0;
wire  [22:0] v$_2232_out0;
wire  [23:0] v$A$MANTISA$COMPARATOR_7501_out0;
wire  [23:0] v$A$MANTISA$COMPARATOR_7502_out0;
wire  [23:0] v$A$MANTISA_3756_out0;
wire  [23:0] v$A$MANTISA_3757_out0;
wire  [23:0] v$A$MANTISSA_13185_out0;
wire  [23:0] v$A$MANTISSA_13186_out0;
wire  [23:0] v$A$VIEW_11027_out0;
wire  [23:0] v$A1_13595_out0;
wire  [23:0] v$A1_13596_out0;
wire  [23:0] v$A1_13597_out0;
wire  [23:0] v$A1_13598_out0;
wire  [23:0] v$A1_13599_out0;
wire  [23:0] v$A1_15214_out0;
wire  [23:0] v$A1_15215_out0;
wire  [23:0] v$A1_15216_out0;
wire  [23:0] v$A1_15217_out0;
wire  [23:0] v$A1_15218_out0;
wire  [23:0] v$A1_15219_out0;
wire  [23:0] v$A1_15220_out0;
wire  [23:0] v$A1_15221_out0;
wire  [23:0] v$A1_15222_out0;
wire  [23:0] v$A1_15223_out0;
wire  [23:0] v$A1_15224_out0;
wire  [23:0] v$A1_15225_out0;
wire  [23:0] v$ADDER$A_3696_out0;
wire  [23:0] v$ADDER$A_3697_out0;
wire  [23:0] v$ADDER$B_6442_out0;
wire  [23:0] v$ADDER$B_6443_out0;
wire  [23:0] v$A_14255_out0;
wire  [23:0] v$A_14801_out0;
wire  [23:0] v$A_3463_out0;
wire  [23:0] v$A_5418_out0;
wire  [23:0] v$B$MANTISA$COMPARATOR_15865_out0;
wire  [23:0] v$B$MANTISA$COMPARATOR_15866_out0;
wire  [23:0] v$B$MANTISA_15588_out0;
wire  [23:0] v$B$MANTISA_15589_out0;
wire  [23:0] v$B$MANTISSA_2673_out0;
wire  [23:0] v$B$MANTISSA_2674_out0;
wire  [23:0] v$B$SHIFTED_13792_out0;
wire  [23:0] v$B$VIEW_5730_out0;
wire  [23:0] v$B2_8415_out0;
wire  [23:0] v$B2_8416_out0;
wire  [23:0] v$B2_8417_out0;
wire  [23:0] v$B2_8418_out0;
wire  [23:0] v$B2_8419_out0;
wire  [23:0] v$B_13561_out0;
wire  [23:0] v$B_1965_out0;
wire  [23:0] v$B_81_out0;
wire  [23:0] v$B_8359_out0;
wire  [23:0] v$C1_16233_out0;
wire  [23:0] v$C1_16234_out0;
wire  [23:0] v$C1_4454_out0;
wire  [23:0] v$C1_4455_out0;
wire  [23:0] v$C1_4456_out0;
wire  [23:0] v$C1_4457_out0;
wire  [23:0] v$C1_4458_out0;
wire  [23:0] v$C1_4459_out0;
wire  [23:0] v$C1_4460_out0;
wire  [23:0] v$C1_4461_out0;
wire  [23:0] v$C2_7814_out0;
wire  [23:0] v$C3_18437_out0;
wire  [23:0] v$C4_17973_out0;
wire  [23:0] v$C5_3961_out0;
wire  [23:0] v$C5_3962_out0;
wire  [23:0] v$C5_3963_out0;
wire  [23:0] v$C5_3964_out0;
wire  [23:0] v$C5_3965_out0;
wire  [23:0] v$C5_3966_out0;
wire  [23:0] v$C5_3967_out0;
wire  [23:0] v$C5_3968_out0;
wire  [23:0] v$C5_3969_out0;
wire  [23:0] v$C5_3970_out0;
wire  [23:0] v$C5_3971_out0;
wire  [23:0] v$C5_3972_out0;
wire  [23:0] v$C7_14643_out0;
wire  [23:0] v$C7_14644_out0;
wire  [23:0] v$C8_13621_out0;
wire  [23:0] v$C8_13622_out0;
wire  [23:0] v$C9_15264_out0;
wire  [23:0] v$C9_15265_out0;
wire  [23:0] v$END1_9929_out0;
wire  [23:0] v$END1_9930_out0;
wire  [23:0] v$END_1870_out0;
wire  [23:0] v$END_1871_out0;
wire  [23:0] v$FINAL$RESULT_2572_out0;
wire  [23:0] v$IGNORE_12634_out0;
wire  [23:0] v$IN_11071_out0;
wire  [23:0] v$IN_11072_out0;
wire  [23:0] v$IN_11642_out0;
wire  [23:0] v$IN_11643_out0;
wire  [23:0] v$IN_11781_out0;
wire  [23:0] v$IN_11782_out0;
wire  [23:0] v$IN_11783_out0;
wire  [23:0] v$IN_11784_out0;
wire  [23:0] v$IN_11785_out0;
wire  [23:0] v$IN_11786_out0;
wire  [23:0] v$IN_11787_out0;
wire  [23:0] v$IN_11790_out0;
wire  [23:0] v$IN_11791_out0;
wire  [23:0] v$IN_11792_out0;
wire  [23:0] v$IN_13165_out0;
wire  [23:0] v$IN_13166_out0;
wire  [23:0] v$IN_13167_out0;
wire  [23:0] v$IN_13168_out0;
wire  [23:0] v$IN_13169_out0;
wire  [23:0] v$IN_13170_out0;
wire  [23:0] v$IN_13171_out0;
wire  [23:0] v$IN_13172_out0;
wire  [23:0] v$IN_13562_out0;
wire  [23:0] v$IN_13564_out0;
wire  [23:0] v$IN_15603_out0;
wire  [23:0] v$IN_15604_out0;
wire  [23:0] v$IN_15605_out0;
wire  [23:0] v$IN_15606_out0;
wire  [23:0] v$IN_15607_out0;
wire  [23:0] v$IN_15608_out0;
wire  [23:0] v$IN_15609_out0;
wire  [23:0] v$IN_15612_out0;
wire  [23:0] v$IN_15613_out0;
wire  [23:0] v$IN_15614_out0;
wire  [23:0] v$IN_17987_out0;
wire  [23:0] v$IN_17988_out0;
wire  [23:0] v$IN_18262_out0;
wire  [23:0] v$IN_18263_out0;
wire  [23:0] v$IN_3856_out0;
wire  [23:0] v$IN_3857_out0;
wire  [23:0] v$IN_3858_out0;
wire  [23:0] v$IN_3859_out0;
wire  [23:0] v$IN_3860_out0;
wire  [23:0] v$IN_3861_out0;
wire  [23:0] v$IN_3862_out0;
wire  [23:0] v$IN_3863_out0;
wire  [23:0] v$IN_3864_out0;
wire  [23:0] v$IN_3865_out0;
wire  [23:0] v$IN_3872_out0;
wire  [23:0] v$IN_3873_out0;
wire  [23:0] v$IN_3874_out0;
wire  [23:0] v$IN_4190_out0;
wire  [23:0] v$IN_4191_out0;
wire  [23:0] v$IN_5018_out0;
wire  [23:0] v$IN_5019_out0;
wire  [23:0] v$IN_5020_out0;
wire  [23:0] v$IN_5021_out0;
wire  [23:0] v$IN_5022_out0;
wire  [23:0] v$IN_5023_out0;
wire  [23:0] v$IN_5024_out0;
wire  [23:0] v$IN_5025_out0;
wire  [23:0] v$IN_5026_out0;
wire  [23:0] v$IN_5027_out0;
wire  [23:0] v$IN_5028_out0;
wire  [23:0] v$IN_5029_out0;
wire  [23:0] v$IN_5032_out0;
wire  [23:0] v$IN_5033_out0;
wire  [23:0] v$IN_5034_out0;
wire  [23:0] v$IN_5035_out0;
wire  [23:0] v$IN_5036_out0;
wire  [23:0] v$IN_5037_out0;
wire  [23:0] v$IN_5147_out0;
wire  [23:0] v$IN_5148_out0;
wire  [23:0] v$IN_5149_out0;
wire  [23:0] v$IN_5150_out0;
wire  [23:0] v$IN_5151_out0;
wire  [23:0] v$IN_5152_out0;
wire  [23:0] v$IN_5153_out0;
wire  [23:0] v$IN_5154_out0;
wire  [23:0] v$IN_5155_out0;
wire  [23:0] v$IN_5156_out0;
wire  [23:0] v$IN_5157_out0;
wire  [23:0] v$IN_5158_out0;
wire  [23:0] v$IN_5159_out0;
wire  [23:0] v$IN_5160_out0;
wire  [23:0] v$IN_5161_out0;
wire  [23:0] v$IN_5162_out0;
wire  [23:0] v$IN_5163_out0;
wire  [23:0] v$IN_5164_out0;
wire  [23:0] v$IN_5165_out0;
wire  [23:0] v$IN_5166_out0;
wire  [23:0] v$IN_5167_out0;
wire  [23:0] v$IN_5168_out0;
wire  [23:0] v$IN_5169_out0;
wire  [23:0] v$IN_5170_out0;
wire  [23:0] v$IN_5171_out0;
wire  [23:0] v$IN_5172_out0;
wire  [23:0] v$IN_5173_out0;
wire  [23:0] v$IN_5174_out0;
wire  [23:0] v$IN_5175_out0;
wire  [23:0] v$IN_5176_out0;
wire  [23:0] v$IN_5177_out0;
wire  [23:0] v$IN_5178_out0;
wire  [23:0] v$IN_5179_out0;
wire  [23:0] v$IN_5180_out0;
wire  [23:0] v$IN_5181_out0;
wire  [23:0] v$IN_5182_out0;
wire  [23:0] v$IN_5195_out0;
wire  [23:0] v$IN_5196_out0;
wire  [23:0] v$IN_5197_out0;
wire  [23:0] v$IN_5198_out0;
wire  [23:0] v$IN_5199_out0;
wire  [23:0] v$IN_5200_out0;
wire  [23:0] v$IN_5201_out0;
wire  [23:0] v$IN_5202_out0;
wire  [23:0] v$IN_5203_out0;
wire  [23:0] v$IN_5204_out0;
wire  [23:0] v$IN_5205_out0;
wire  [23:0] v$IN_5206_out0;
wire  [23:0] v$IN_5207_out0;
wire  [23:0] v$IN_5208_out0;
wire  [23:0] v$IN_5209_out0;
wire  [23:0] v$IN_8294_out0;
wire  [23:0] v$IN_8295_out0;
wire  [23:0] v$LZD$INPUT_8837_out0;
wire  [23:0] v$LZD$INPUT_8838_out0;
wire  [23:0] v$MULTIPLIER$OUT_14973_out0;
wire  [23:0] v$MULTIPLIER$OUT_9343_out0;
wire  [23:0] v$MULTIPLIER_3669_out0;
wire  [23:0] v$MULTIPLIER_3671_out0;
wire  [23:0] v$MULTIPLIER_3672_out0;
wire  [23:0] v$MULTIPLIER_3673_out0;
wire  [23:0] v$MULTIPLIER_3674_out0;
wire  [23:0] v$MULTIPLIER_3675_out0;
wire  [23:0] v$MULTIPLIER_3676_out0;
wire  [23:0] v$MULTIPLIER_3677_out0;
wire  [23:0] v$MULTIPLIER_3678_out0;
wire  [23:0] v$MULTIPLIER_3679_out0;
wire  [23:0] v$MULTIPLIER_3680_out0;
wire  [23:0] v$MULTIPLIER_6355_out0;
wire  [23:0] v$MUX1_11630_out0;
wire  [23:0] v$MUX1_11631_out0;
wire  [23:0] v$MUX1_11632_out0;
wire  [23:0] v$MUX1_11633_out0;
wire  [23:0] v$MUX1_11634_out0;
wire  [23:0] v$MUX1_11635_out0;
wire  [23:0] v$MUX1_11636_out0;
wire  [23:0] v$MUX1_11637_out0;
wire  [23:0] v$MUX1_14183_out0;
wire  [23:0] v$MUX1_14184_out0;
wire  [23:0] v$MUX1_2349_out0;
wire  [23:0] v$MUX1_2350_out0;
wire  [23:0] v$MUX1_2351_out0;
wire  [23:0] v$MUX1_2352_out0;
wire  [23:0] v$MUX1_2353_out0;
wire  [23:0] v$MUX1_2354_out0;
wire  [23:0] v$MUX1_2355_out0;
wire  [23:0] v$MUX1_2356_out0;
wire  [23:0] v$MUX1_2357_out0;
wire  [23:0] v$MUX1_2358_out0;
wire  [23:0] v$MUX1_2359_out0;
wire  [23:0] v$MUX1_2360_out0;
wire  [23:0] v$MUX1_2361_out0;
wire  [23:0] v$MUX1_2362_out0;
wire  [23:0] v$MUX1_2363_out0;
wire  [23:0] v$MUX1_2364_out0;
wire  [23:0] v$MUX1_2365_out0;
wire  [23:0] v$MUX1_2366_out0;
wire  [23:0] v$MUX1_2367_out0;
wire  [23:0] v$MUX1_2368_out0;
wire  [23:0] v$MUX1_2369_out0;
wire  [23:0] v$MUX1_2370_out0;
wire  [23:0] v$MUX1_2371_out0;
wire  [23:0] v$MUX1_2372_out0;
wire  [23:0] v$MUX1_2373_out0;
wire  [23:0] v$MUX1_2374_out0;
wire  [23:0] v$MUX1_2375_out0;
wire  [23:0] v$MUX1_2376_out0;
wire  [23:0] v$MUX1_2377_out0;
wire  [23:0] v$MUX1_2378_out0;
wire  [23:0] v$MUX1_2379_out0;
wire  [23:0] v$MUX1_2380_out0;
wire  [23:0] v$MUX1_2381_out0;
wire  [23:0] v$MUX1_2382_out0;
wire  [23:0] v$MUX1_2383_out0;
wire  [23:0] v$MUX1_2384_out0;
wire  [23:0] v$MUX1_2397_out0;
wire  [23:0] v$MUX1_2398_out0;
wire  [23:0] v$MUX1_2399_out0;
wire  [23:0] v$MUX1_2400_out0;
wire  [23:0] v$MUX1_2401_out0;
wire  [23:0] v$MUX1_2402_out0;
wire  [23:0] v$MUX1_2403_out0;
wire  [23:0] v$MUX1_2404_out0;
wire  [23:0] v$MUX1_2405_out0;
wire  [23:0] v$MUX1_2406_out0;
wire  [23:0] v$MUX1_2407_out0;
wire  [23:0] v$MUX1_2408_out0;
wire  [23:0] v$MUX1_2409_out0;
wire  [23:0] v$MUX1_2410_out0;
wire  [23:0] v$MUX1_2411_out0;
wire  [23:0] v$MUX1_2888_out0;
wire  [23:0] v$MUX1_8338_out0;
wire  [23:0] v$MUX1_8339_out0;
wire  [23:0] v$MUX1_8340_out0;
wire  [23:0] v$MUX1_8341_out0;
wire  [23:0] v$MUX1_8342_out0;
wire  [23:0] v$MUX1_8343_out0;
wire  [23:0] v$MUX1_8344_out0;
wire  [23:0] v$MUX1_8345_out0;
wire  [23:0] v$MUX1_8346_out0;
wire  [23:0] v$MUX1_8347_out0;
wire  [23:0] v$MUX1_8348_out0;
wire  [23:0] v$MUX1_8349_out0;
wire  [23:0] v$MUX2_12458_out0;
wire  [23:0] v$MUX2_14827_out0;
wire  [23:0] v$MUX2_14828_out0;
wire  [23:0] v$MUX2_14829_out0;
wire  [23:0] v$MUX2_15234_out0;
wire  [23:0] v$MUX2_15235_out0;
wire  [23:0] v$MUX2_15236_out0;
wire  [23:0] v$MUX2_15237_out0;
wire  [23:0] v$MUX2_15238_out0;
wire  [23:0] v$MUX2_15239_out0;
wire  [23:0] v$MUX2_15240_out0;
wire  [23:0] v$MUX2_15243_out0;
wire  [23:0] v$MUX2_15244_out0;
wire  [23:0] v$MUX2_15245_out0;
wire  [23:0] v$MUX2_18043_out0;
wire  [23:0] v$MUX2_18573_out0;
wire  [23:0] v$MUX2_18574_out0;
wire  [23:0] v$MUX2_18575_out0;
wire  [23:0] v$MUX2_18576_out0;
wire  [23:0] v$MUX2_18577_out0;
wire  [23:0] v$MUX2_18578_out0;
wire  [23:0] v$MUX2_18579_out0;
wire  [23:0] v$MUX2_18586_out0;
wire  [23:0] v$MUX2_18587_out0;
wire  [23:0] v$MUX2_18588_out0;
wire  [23:0] v$MUX2_2475_out0;
wire  [23:0] v$MUX2_2476_out0;
wire  [23:0] v$MUX2_2477_out0;
wire  [23:0] v$MUX2_2478_out0;
wire  [23:0] v$MUX2_2479_out0;
wire  [23:0] v$MUX2_2480_out0;
wire  [23:0] v$MUX2_2481_out0;
wire  [23:0] v$MUX2_2484_out0;
wire  [23:0] v$MUX2_2485_out0;
wire  [23:0] v$MUX2_2486_out0;
wire  [23:0] v$MUX2_2492_out0;
wire  [23:0] v$MUX2_2493_out0;
wire  [23:0] v$MUX2_2494_out0;
wire  [23:0] v$MUX2_2495_out0;
wire  [23:0] v$MUX2_2496_out0;
wire  [23:0] v$MUX2_2497_out0;
wire  [23:0] v$MUX2_2498_out0;
wire  [23:0] v$MUX2_2499_out0;
wire  [23:0] v$MUX2_2500_out0;
wire  [23:0] v$MUX2_2501_out0;
wire  [23:0] v$MUX2_2502_out0;
wire  [23:0] v$MUX2_2503_out0;
wire  [23:0] v$MUX2_2506_out0;
wire  [23:0] v$MUX2_2507_out0;
wire  [23:0] v$MUX2_2508_out0;
wire  [23:0] v$MUX2_2509_out0;
wire  [23:0] v$MUX2_2510_out0;
wire  [23:0] v$MUX2_2511_out0;
wire  [23:0] v$MUX3_12800_out0;
wire  [23:0] v$MUX3_12801_out0;
wire  [23:0] v$MUX3_17902_out0;
wire  [23:0] v$MUX3_3107_out0;
wire  [23:0] v$MUX3_3108_out0;
wire  [23:0] v$MUX3_3771_out0;
wire  [23:0] v$MUX3_3772_out0;
wire  [23:0] v$MUX3_7636_out0;
wire  [23:0] v$MUX4_5890_out0;
wire  [23:0] v$MUX4_5891_out0;
wire  [23:0] v$MUX4_8103_out0;
wire  [23:0] v$MUX5_10310_out0;
wire  [23:0] v$MUX5_1611_out0;
wire  [23:0] v$MUX5_1612_out0;
wire  [23:0] v$MUX5_6222_out0;
wire  [23:0] v$MUX5_6223_out0;
wire  [23:0] v$MUX7_3280_out0;
wire  [23:0] v$MUX7_3281_out0;
wire  [23:0] v$MUX8_5397_out0;
wire  [23:0] v$MUX8_5398_out0;
wire  [23:0] v$MUX9_2458_out0;
wire  [23:0] v$MUX9_2459_out0;
wire  [23:0] v$OP1$MANTISA$ADDER_3643_out0;
wire  [23:0] v$OP1$MANTISA$ADDER_3644_out0;
wire  [23:0] v$OP1$MANTISA$MULTIPLY_11887_out0;
wire  [23:0] v$OP1$MANTISA$MULTIPLY_11888_out0;
wire  [23:0] v$OP1$MANTISA_11806_out0;
wire  [23:0] v$OP1$MANTISA_11807_out0;
wire  [23:0] v$OP1$MANTISA_3789_out0;
wire  [23:0] v$OP1$MANTISA_3790_out0;
wire  [23:0] v$OP1$MANTISA_9121_out0;
wire  [23:0] v$OP1$MANTISA_9122_out0;
wire  [23:0] v$OP1_14185_out0;
wire  [23:0] v$OP1_14186_out0;
wire  [23:0] v$OP1_14187_out0;
wire  [23:0] v$OP1_14188_out0;
wire  [23:0] v$OP1_14189_out0;
wire  [23:0] v$OP1_14190_out0;
wire  [23:0] v$OP1_14191_out0;
wire  [23:0] v$OP1_14192_out0;
wire  [23:0] v$OP1_14193_out0;
wire  [23:0] v$OP1_14194_out0;
wire  [23:0] v$OP1_14195_out0;
wire  [23:0] v$OP1_14196_out0;
wire  [23:0] v$OP1_3379_out0;
wire  [23:0] v$OP1_3380_out0;
wire  [23:0] v$OP1_3381_out0;
wire  [23:0] v$OP1_3382_out0;
wire  [23:0] v$OP1_3383_out0;
wire  [23:0] v$OP1_3384_out0;
wire  [23:0] v$OP1_3385_out0;
wire  [23:0] v$OP1_3386_out0;
wire  [23:0] v$OP1_3387_out0;
wire  [23:0] v$OP1_3388_out0;
wire  [23:0] v$OP1_3389_out0;
wire  [23:0] v$OP1_3390_out0;
wire  [23:0] v$OP1_4100_out0;
wire  [23:0] v$OP1_4101_out0;
wire  [23:0] v$OP2$MANTISA$ADDER_7490_out0;
wire  [23:0] v$OP2$MANTISA$ADDER_7491_out0;
wire  [23:0] v$OP2$MANTISA$MULTIPLY_2462_out0;
wire  [23:0] v$OP2$MANTISA$MULTIPLY_2463_out0;
wire  [23:0] v$OP2$MANTISA_2656_out0;
wire  [23:0] v$OP2$MANTISA_2657_out0;
wire  [23:0] v$OP2$MANTISA_3510_out0;
wire  [23:0] v$OP2$MANTISA_3511_out0;
wire  [23:0] v$OP2$MANTISA_9544_out0;
wire  [23:0] v$OP2$MANTISA_9545_out0;
wire  [23:0] v$OP2_10374_out0;
wire  [23:0] v$OP2_10375_out0;
wire  [23:0] v$OP2_10376_out0;
wire  [23:0] v$OP2_10377_out0;
wire  [23:0] v$OP2_10378_out0;
wire  [23:0] v$OP2_10379_out0;
wire  [23:0] v$OP2_10380_out0;
wire  [23:0] v$OP2_10381_out0;
wire  [23:0] v$OP2_10382_out0;
wire  [23:0] v$OP2_10383_out0;
wire  [23:0] v$OP2_10384_out0;
wire  [23:0] v$OP2_10385_out0;
wire  [23:0] v$OP2_12455_out0;
wire  [23:0] v$OP2_3670_out0;
wire  [23:0] v$OP2_4162_out0;
wire  [23:0] v$OP2_4163_out0;
wire  [23:0] v$OP2_4862_out0;
wire  [23:0] v$OP2_6354_out0;
wire  [23:0] v$OP2_6356_out0;
wire  [23:0] v$OP2_6357_out0;
wire  [23:0] v$OP2_6358_out0;
wire  [23:0] v$OP2_6359_out0;
wire  [23:0] v$OP2_6360_out0;
wire  [23:0] v$OP2_6361_out0;
wire  [23:0] v$OP2_6362_out0;
wire  [23:0] v$OP2_6363_out0;
wire  [23:0] v$OP2_6364_out0;
wire  [23:0] v$OP2_6365_out0;
wire  [23:0] v$OUT_10011_out0;
wire  [23:0] v$OUT_10012_out0;
wire  [23:0] v$OUT_10013_out0;
wire  [23:0] v$OUT_10014_out0;
wire  [23:0] v$OUT_10015_out0;
wire  [23:0] v$OUT_10016_out0;
wire  [23:0] v$OUT_10017_out0;
wire  [23:0] v$OUT_10018_out0;
wire  [23:0] v$OUT_14901_out0;
wire  [23:0] v$OUT_14902_out0;
wire  [23:0] v$OUT_14903_out0;
wire  [23:0] v$OUT_14904_out0;
wire  [23:0] v$OUT_14905_out0;
wire  [23:0] v$OUT_14906_out0;
wire  [23:0] v$OUT_14907_out0;
wire  [23:0] v$OUT_14908_out0;
wire  [23:0] v$OUT_14909_out0;
wire  [23:0] v$OUT_14910_out0;
wire  [23:0] v$OUT_14911_out0;
wire  [23:0] v$OUT_14912_out0;
wire  [23:0] v$OUT_14913_out0;
wire  [23:0] v$OUT_14914_out0;
wire  [23:0] v$OUT_14915_out0;
wire  [23:0] v$OUT_14916_out0;
wire  [23:0] v$OUT_14917_out0;
wire  [23:0] v$OUT_14918_out0;
wire  [23:0] v$OUT_14919_out0;
wire  [23:0] v$OUT_14920_out0;
wire  [23:0] v$OUT_14921_out0;
wire  [23:0] v$OUT_14922_out0;
wire  [23:0] v$OUT_14923_out0;
wire  [23:0] v$OUT_14924_out0;
wire  [23:0] v$OUT_14925_out0;
wire  [23:0] v$OUT_14926_out0;
wire  [23:0] v$OUT_14927_out0;
wire  [23:0] v$OUT_14928_out0;
wire  [23:0] v$OUT_14929_out0;
wire  [23:0] v$OUT_14930_out0;
wire  [23:0] v$OUT_14931_out0;
wire  [23:0] v$OUT_14932_out0;
wire  [23:0] v$OUT_14933_out0;
wire  [23:0] v$OUT_14934_out0;
wire  [23:0] v$OUT_14935_out0;
wire  [23:0] v$OUT_14936_out0;
wire  [23:0] v$OUT_14949_out0;
wire  [23:0] v$OUT_14950_out0;
wire  [23:0] v$OUT_14951_out0;
wire  [23:0] v$OUT_14952_out0;
wire  [23:0] v$OUT_14953_out0;
wire  [23:0] v$OUT_14954_out0;
wire  [23:0] v$OUT_14955_out0;
wire  [23:0] v$OUT_14956_out0;
wire  [23:0] v$OUT_14957_out0;
wire  [23:0] v$OUT_14958_out0;
wire  [23:0] v$OUT_14959_out0;
wire  [23:0] v$OUT_14960_out0;
wire  [23:0] v$OUT_14961_out0;
wire  [23:0] v$OUT_14962_out0;
wire  [23:0] v$OUT_14963_out0;
wire  [23:0] v$OUT_4913_out0;
wire  [23:0] v$OUT_4914_out0;
wire  [23:0] v$RESULT_5062_out0;
wire  [23:0] v$SEL6_5757_out0;
wire  [23:0] v$SUM$EXEC1_18543_out0;
wire  [23:0] v$SUM$HALF_2883_out0;
wire  [23:0] v$SUM1_12827_out0;
wire  [23:0] v$SUM1_12828_out0;
wire  [23:0] v$SUM1_12829_out0;
wire  [23:0] v$SUM1_12830_out0;
wire  [23:0] v$SUM1_12831_out0;
wire  [23:0] v$SUM1_5431_out0;
wire  [23:0] v$SUM_15166_out0;
wire  [23:0] v$SUM_15167_out0;
wire  [23:0] v$SUM_15168_out0;
wire  [23:0] v$SUM_15169_out0;
wire  [23:0] v$SUM_15170_out0;
wire  [23:0] v$SUM_15171_out0;
wire  [23:0] v$SUM_15172_out0;
wire  [23:0] v$SUM_15173_out0;
wire  [23:0] v$SUM_15174_out0;
wire  [23:0] v$SUM_15175_out0;
wire  [23:0] v$SUM_15176_out0;
wire  [23:0] v$SUM_15177_out0;
wire  [23:0] v$SUM_1905_out0;
wire  [23:0] v$SUM_1906_out0;
wire  [23:0] v$SUM_3466_out0;
wire  [23:0] v$SUM_3467_out0;
wire  [23:0] v$SUM_3468_out0;
wire  [23:0] v$SUM_3469_out0;
wire  [23:0] v$SUM_3470_out0;
wire  [23:0] v$SUM_3471_out0;
wire  [23:0] v$SUM_3472_out0;
wire  [23:0] v$SUM_3473_out0;
wire  [23:0] v$SUM_3474_out0;
wire  [23:0] v$SUM_3475_out0;
wire  [23:0] v$SUM_3476_out0;
wire  [23:0] v$SUM_3477_out0;
wire  [23:0] v$SUM_892_out0;
wire  [23:0] v$SUM_9362_out0;
wire  [23:0] v$SUM_9363_out0;
wire  [23:0] v$SUM_9364_out0;
wire  [23:0] v$SUM_9365_out0;
wire  [23:0] v$SUM_9366_out0;
wire  [23:0] v$XOR$IN_2245_out0;
wire  [23:0] v$XOR$IN_2246_out0;
wire  [23:0] v$XOR1_5399_out0;
wire  [23:0] v$XOR1_5400_out0;
wire  [23:0] v$XOR2_7849_out0;
wire  [23:0] v$XOR2_7850_out0;
wire  [23:0] v$_10038_out0;
wire  [23:0] v$_10039_out0;
wire  [23:0] v$_11015_out0;
wire  [23:0] v$_11016_out0;
wire  [23:0] v$_1158_out0;
wire  [23:0] v$_14091_out0;
wire  [23:0] v$_14092_out0;
wire  [23:0] v$_1510_out0;
wire  [23:0] v$_1511_out0;
wire  [23:0] v$_15349_out0;
wire  [23:0] v$_15350_out0;
wire  [23:0] v$_17770_out0;
wire  [23:0] v$_17771_out0;
wire  [23:0] v$_17993_out0;
wire  [23:0] v$_17994_out0;
wire  [23:0] v$_17995_out0;
wire  [23:0] v$_17996_out0;
wire  [23:0] v$_17997_out0;
wire  [23:0] v$_17998_out0;
wire  [23:0] v$_17999_out0;
wire  [23:0] v$_18000_out0;
wire  [23:0] v$_18001_out0;
wire  [23:0] v$_18002_out0;
wire  [23:0] v$_18003_out0;
wire  [23:0] v$_18004_out0;
wire  [23:0] v$_3759_out0;
wire  [23:0] v$_3760_out0;
wire  [23:0] v$_3761_out0;
wire  [23:0] v$_3762_out0;
wire  [23:0] v$_3763_out0;
wire  [23:0] v$_4245_out0;
wire  [23:0] v$_4246_out0;
wire  [23:0] v$_4247_out0;
wire  [23:0] v$_4248_out0;
wire  [23:0] v$_4249_out0;
wire  [23:0] v$_4250_out0;
wire  [23:0] v$_4251_out0;
wire  [23:0] v$_4252_out0;
wire  [23:0] v$_4253_out0;
wire  [23:0] v$_4254_out0;
wire  [23:0] v$_4255_out0;
wire  [23:0] v$_4256_out0;
wire  [23:0] v$_4257_out0;
wire  [23:0] v$_4258_out0;
wire  [23:0] v$_4259_out0;
wire  [23:0] v$_4260_out0;
wire  [23:0] v$_4261_out0;
wire  [23:0] v$_4262_out0;
wire  [23:0] v$_4263_out0;
wire  [23:0] v$_4264_out0;
wire  [23:0] v$_4265_out0;
wire  [23:0] v$_4266_out0;
wire  [23:0] v$_4267_out0;
wire  [23:0] v$_4268_out0;
wire  [23:0] v$_4269_out0;
wire  [23:0] v$_4270_out0;
wire  [23:0] v$_4271_out0;
wire  [23:0] v$_4272_out0;
wire  [23:0] v$_4273_out0;
wire  [23:0] v$_4274_out0;
wire  [23:0] v$_4275_out0;
wire  [23:0] v$_4276_out0;
wire  [23:0] v$_4277_out0;
wire  [23:0] v$_4278_out0;
wire  [23:0] v$_4279_out0;
wire  [23:0] v$_4280_out0;
wire  [23:0] v$_4293_out0;
wire  [23:0] v$_4294_out0;
wire  [23:0] v$_4295_out0;
wire  [23:0] v$_4296_out0;
wire  [23:0] v$_4297_out0;
wire  [23:0] v$_4298_out0;
wire  [23:0] v$_4299_out0;
wire  [23:0] v$_4300_out0;
wire  [23:0] v$_4301_out0;
wire  [23:0] v$_4302_out0;
wire  [23:0] v$_4303_out0;
wire  [23:0] v$_4304_out0;
wire  [23:0] v$_4305_out0;
wire  [23:0] v$_4306_out0;
wire  [23:0] v$_4307_out0;
wire  [23:0] v$_7380_out0;
wire  [23:0] v$_7418_out0;
wire  [23:0] v$_7419_out0;
wire  [23:0] v$_7615_out0;
wire  [23:0] v$_7616_out0;
wire  [23:0] v$_8980_out0;
wire  [23:0] v$_8981_out0;
wire  [23:0] v$_8982_out0;
wire  [23:0] v$_8983_out0;
wire  [23:0] v$_8984_out0;
wire  [23:0] v$_8985_out0;
wire  [23:0] v$_8986_out0;
wire  [23:0] v$_8987_out0;
wire  [23:0] v$_8988_out0;
wire  [23:0] v$_8989_out0;
wire  [23:0] v$_8990_out0;
wire  [23:0] v$_8991_out0;
wire  [23:0] v$_8992_out0;
wire  [23:0] v$_8993_out0;
wire  [23:0] v$_8994_out0;
wire  [23:0] v$_8995_out0;
wire  [23:0] v$_8996_out0;
wire  [23:0] v$_8997_out0;
wire  [23:0] v$_8998_out0;
wire  [23:0] v$_8999_out0;
wire  [23:0] v$_9000_out0;
wire  [23:0] v$_9001_out0;
wire  [23:0] v$_9002_out0;
wire  [23:0] v$_9003_out0;
wire  [23:0] v$_9004_out0;
wire  [23:0] v$_9005_out0;
wire  [23:0] v$_9006_out0;
wire  [23:0] v$_9007_out0;
wire  [23:0] v$_9008_out0;
wire  [23:0] v$_9009_out0;
wire  [23:0] v$_9010_out0;
wire  [23:0] v$_9011_out0;
wire  [23:0] v$_9012_out0;
wire  [23:0] v$_9013_out0;
wire  [23:0] v$_9014_out0;
wire  [23:0] v$_9015_out0;
wire  [23:0] v$_9028_out0;
wire  [23:0] v$_9029_out0;
wire  [23:0] v$_9030_out0;
wire  [23:0] v$_9031_out0;
wire  [23:0] v$_9032_out0;
wire  [23:0] v$_9033_out0;
wire  [23:0] v$_9034_out0;
wire  [23:0] v$_9035_out0;
wire  [23:0] v$_9036_out0;
wire  [23:0] v$_9037_out0;
wire  [23:0] v$_9038_out0;
wire  [23:0] v$_9039_out0;
wire  [23:0] v$_9040_out0;
wire  [23:0] v$_9041_out0;
wire  [23:0] v$_9042_out0;
wire  [23:0] v$_9906_out0;
wire  [23:0] v$_9907_out0;
wire  [23:0] v$_9908_out0;
wire  [23:0] v$_9909_out0;
wire  [23:0] v$_9910_out0;
wire  [24:0] v$_10453_out0;
wire  [24:0] v$_18087_out0;
wire  [25:0] v$_11764_out0;
wire  [25:0] v$_4910_out0;
wire  [26:0] v$_13990_out0;
wire  [26:0] v$_7621_out0;
wire  [27:0] v$_10037_out0;
wire  [27:0] v$_4158_out0;
wire  [27:0] v$_9931_out0;
wire  [27:0] v$_9932_out0;
wire  [28:0] v$_15111_out0;
wire  [28:0] v$_16351_out0;
wire  [29:0] v$_17404_out0;
wire  [29:0] v$_1971_out0;
wire  [2:0] v$9_14162_out0;
wire  [2:0] v$9_14163_out0;
wire  [2:0] v$ALU$OP_16826_out0;
wire  [2:0] v$ALU$OP_16827_out0;
wire  [2:0] v$C10_13540_out0;
wire  [2:0] v$C10_13541_out0;
wire  [2:0] v$C1_16842_out0;
wire  [2:0] v$C1_16843_out0;
wire  [2:0] v$C2_13325_out0;
wire  [2:0] v$C2_13326_out0;
wire  [2:0] v$C4_6625_out0;
wire  [2:0] v$C4_6626_out0;
wire  [2:0] v$IR1$OP_5519_out0;
wire  [2:0] v$IR1$OP_5520_out0;
wire  [2:0] v$IR2$OP_15861_out0;
wire  [2:0] v$IR2$OP_15862_out0;
wire  [2:0] v$IR2$OP_18020_out0;
wire  [2:0] v$IR2$OP_18021_out0;
wire  [2:0] v$MODE_1617_out0;
wire  [2:0] v$MODE_1618_out0;
wire  [2:0] v$MODE_9126_out0;
wire  [2:0] v$MODE_9127_out0;
wire  [2:0] v$MUX1_14693_out0;
wire  [2:0] v$MUX1_14694_out0;
wire  [2:0] v$MUX1_14695_out0;
wire  [2:0] v$MUX1_14696_out0;
wire  [2:0] v$MUX1_14697_out0;
wire  [2:0] v$MUX1_14698_out0;
wire  [2:0] v$MUX1_14699_out0;
wire  [2:0] v$MUX1_14700_out0;
wire  [2:0] v$Mode_10976_out0;
wire  [2:0] v$Mode_10977_out0;
wire  [2:0] v$Mode_13197_out0;
wire  [2:0] v$Mode_13198_out0;
wire  [2:0] v$NUPPER_17364_out0;
wire  [2:0] v$NUPPER_17365_out0;
wire  [2:0] v$NUPPER_17366_out0;
wire  [2:0] v$NUPPER_17367_out0;
wire  [2:0] v$OPCODE_7892_out0;
wire  [2:0] v$OPCODE_7893_out0;
wire  [2:0] v$OP_17642_out0;
wire  [2:0] v$OP_17643_out0;
wire  [2:0] v$OP_1872_out0;
wire  [2:0] v$OP_1873_out0;
wire  [2:0] v$SEL26_4837_out0;
wire  [2:0] v$SEL26_4838_out0;
wire  [2:0] v$SEL26_4839_out0;
wire  [2:0] v$SEL26_4840_out0;
wire  [2:0] v$Y_7756_out0;
wire  [2:0] v$Y_7757_out0;
wire  [2:0] v$Y_7758_out0;
wire  [2:0] v$Y_7759_out0;
wire  [2:0] v$Y_7760_out0;
wire  [2:0] v$Y_7761_out0;
wire  [2:0] v$Y_7762_out0;
wire  [2:0] v$Y_7763_out0;
wire  [2:0] v$_10048_out0;
wire  [2:0] v$_10048_out1;
wire  [2:0] v$_10049_out0;
wire  [2:0] v$_10049_out1;
wire  [2:0] v$_10050_out0;
wire  [2:0] v$_10050_out1;
wire  [2:0] v$_10051_out0;
wire  [2:0] v$_10051_out1;
wire  [2:0] v$_10052_out0;
wire  [2:0] v$_10052_out1;
wire  [2:0] v$_12987_out0;
wire  [2:0] v$_12987_out1;
wire  [2:0] v$_12988_out0;
wire  [2:0] v$_12988_out1;
wire  [2:0] v$_12989_out0;
wire  [2:0] v$_12989_out1;
wire  [2:0] v$_12990_out0;
wire  [2:0] v$_12990_out1;
wire  [2:0] v$_12991_out0;
wire  [2:0] v$_12991_out1;
wire  [2:0] v$_13741_out0;
wire  [2:0] v$_13741_out1;
wire  [2:0] v$_13742_out0;
wire  [2:0] v$_13742_out1;
wire  [2:0] v$_13743_out0;
wire  [2:0] v$_13743_out1;
wire  [2:0] v$_13744_out0;
wire  [2:0] v$_13744_out1;
wire  [2:0] v$_13745_out0;
wire  [2:0] v$_13745_out1;
wire  [2:0] v$_13770_out0;
wire  [2:0] v$_13770_out1;
wire  [2:0] v$_13771_out0;
wire  [2:0] v$_13771_out1;
wire  [2:0] v$_13772_out0;
wire  [2:0] v$_13772_out1;
wire  [2:0] v$_13773_out0;
wire  [2:0] v$_13773_out1;
wire  [2:0] v$_13774_out0;
wire  [2:0] v$_13774_out1;
wire  [2:0] v$_16682_out0;
wire  [2:0] v$_16683_out0;
wire  [2:0] v$_17732_out0;
wire  [2:0] v$_17732_out1;
wire  [2:0] v$_17733_out0;
wire  [2:0] v$_17733_out1;
wire  [2:0] v$_17734_out0;
wire  [2:0] v$_17734_out1;
wire  [2:0] v$_17735_out0;
wire  [2:0] v$_17735_out1;
wire  [2:0] v$_17736_out0;
wire  [2:0] v$_17736_out1;
wire  [2:0] v$_18420_out0;
wire  [2:0] v$_18420_out1;
wire  [2:0] v$_18421_out0;
wire  [2:0] v$_18421_out1;
wire  [2:0] v$_18422_out0;
wire  [2:0] v$_18422_out1;
wire  [2:0] v$_18423_out0;
wire  [2:0] v$_18423_out1;
wire  [2:0] v$_18424_out0;
wire  [2:0] v$_18424_out1;
wire  [2:0] v$_18544_out0;
wire  [2:0] v$_18545_out0;
wire  [2:0] v$_1863_out0;
wire  [2:0] v$_1863_out1;
wire  [2:0] v$_1864_out0;
wire  [2:0] v$_1864_out1;
wire  [2:0] v$_1865_out0;
wire  [2:0] v$_1865_out1;
wire  [2:0] v$_1866_out0;
wire  [2:0] v$_1866_out1;
wire  [2:0] v$_1867_out0;
wire  [2:0] v$_1867_out1;
wire  [2:0] v$_4896_out0;
wire  [2:0] v$_4897_out0;
wire  [2:0] v$_4997_out0;
wire  [2:0] v$_4998_out0;
wire  [2:0] v$_5466_out0;
wire  [2:0] v$_5467_out0;
wire  [2:0] v$_5468_out0;
wire  [2:0] v$_5469_out0;
wire  [2:0] v$_5470_out0;
wire  [2:0] v$_5471_out0;
wire  [2:0] v$_5472_out0;
wire  [2:0] v$_5473_out0;
wire  [2:0] v$_8101_out0;
wire  [2:0] v$_8102_out0;
wire  [2:0] v$_8148_out0;
wire  [2:0] v$_8149_out0;
wire  [2:0] v$_8150_out0;
wire  [2:0] v$_8151_out0;
wire  [2:0] v$_8152_out0;
wire  [2:0] v$_8153_out0;
wire  [2:0] v$_8154_out0;
wire  [2:0] v$_8155_out0;
wire  [2:0] v$_9933_out0;
wire  [2:0] v$_9933_out1;
wire  [2:0] v$_9934_out0;
wire  [2:0] v$_9934_out1;
wire  [2:0] v$_9935_out0;
wire  [2:0] v$_9935_out1;
wire  [2:0] v$_9936_out0;
wire  [2:0] v$_9936_out1;
wire  [2:0] v$_9937_out0;
wire  [2:0] v$_9937_out1;
wire  [30:0] v$C4_8257_out0;
wire  [30:0] v$C4_8259_out0;
wire  [30:0] v$MUX12_15140_out0;
wire  [30:0] v$MUX12_15141_out0;
wire  [30:0] v$MUX2_13631_out0;
wire  [30:0] v$MUX2_13633_out0;
wire  [30:0] v$MUX6_17434_out0;
wire  [30:0] v$MUX6_17435_out0;
wire  [30:0] v$SINGLE$MERGE_12120_out0;
wire  [30:0] v$SINGLE$MERGE_12121_out0;
wire  [30:0] v$_11831_out0;
wire  [30:0] v$_11832_out0;
wire  [30:0] v$_12651_out0;
wire  [30:0] v$_15351_out0;
wire  [30:0] v$_15352_out0;
wire  [30:0] v$_15847_out0;
wire  [30:0] v$_15849_out0;
wire  [30:0] v$_56_out0;
wire  [30:0] v$_57_out0;
wire  [30:0] v$_7021_out0;
wire  [30:0] v$_7022_out0;
wire  [30:0] v$_8260_out0;
wire  [31:0] v$A$32$BIT$MUL_3783_out0;
wire  [31:0] v$A$32$BIT$MUL_3784_out0;
wire  [31:0] v$A$32$BIT_16831_out0;
wire  [31:0] v$A$32$BIT_18440_out0;
wire  [31:0] v$A$32BIT_2990_out0;
wire  [31:0] v$A$32BIT_2991_out0;
wire  [31:0] v$A$FPU$ADDER$32$BIT_15887_out0;
wire  [31:0] v$A$FPU$ADDER$32$BIT_15888_out0;
wire  [31:0] v$A_13812_out0;
wire  [31:0] v$A_13814_out0;
wire  [31:0] v$A_13816_out0;
wire  [31:0] v$A_13818_out0;
wire  [31:0] v$B$32$BIT$FPU$ADDER_10189_out0;
wire  [31:0] v$B$32$BIT$FPU$ADDER_10190_out0;
wire  [31:0] v$B$32$BIT_17689_out0;
wire  [31:0] v$B$32$BIT_1896_out0;
wire  [31:0] v$B$32$MUL_13254_out0;
wire  [31:0] v$B$32$MUL_13255_out0;
wire  [31:0] v$B$32BIT_18471_out0;
wire  [31:0] v$B$32BIT_18472_out0;
wire  [31:0] v$B_4826_out0;
wire  [31:0] v$B_4828_out0;
wire  [31:0] v$B_4830_out0;
wire  [31:0] v$B_4832_out0;
wire  [31:0] v$C1_15226_out0;
wire  [31:0] v$C1_15227_out0;
wire  [31:0] v$C1_5997_out0;
wire  [31:0] v$C1_6003_out0;
wire  [31:0] v$C2_139_out0;
wire  [31:0] v$C2_145_out0;
wire  [31:0] v$C4_14026_out0;
wire  [31:0] v$C4_14027_out0;
wire  [31:0] v$C5_4112_out0;
wire  [31:0] v$C5_4113_out0;
wire  [31:0] v$FPU$ADDER$OUT_4009_out0;
wire  [31:0] v$FPU$ADDER$OUT_4010_out0;
wire  [31:0] v$FPU$ADDER$OUT_5784_out0;
wire  [31:0] v$FPU$ADDER$OUT_5785_out0;
wire  [31:0] v$FPU$MULTIPLIER$OUT_10921_out0;
wire  [31:0] v$FPU$MULTIPLIER$OUT_10922_out0;
wire  [31:0] v$HALF$PRECISION$32$BIT_14802_out0;
wire  [31:0] v$HALF$PRECISION$32$BIT_14803_out0;
wire  [31:0] v$HALF$PRECISION_10311_out0;
wire  [31:0] v$HALF$PRECISION_10312_out0;
wire  [31:0] v$MUX12_16796_out0;
wire  [31:0] v$MUX12_16797_out0;
wire  [31:0] v$MUX13_10727_out0;
wire  [31:0] v$MUX14_1189_out0;
wire  [31:0] v$MUX1_13555_out0;
wire  [31:0] v$MUX1_13556_out0;
wire  [31:0] v$MUX2_16229_out0;
wire  [31:0] v$MUX2_16230_out0;
wire  [31:0] v$MUX3_8965_out0;
wire  [31:0] v$MUX3_8966_out0;
wire  [31:0] v$MUX4_1257_out0;
wire  [31:0] v$MUX4_1258_out0;
wire  [31:0] v$MUX7_4863_out0;
wire  [31:0] v$MUX7_4864_out0;
wire  [31:0] v$OUT1_17809_out0;
wire  [31:0] v$OUT1_17810_out0;
wire  [31:0] v$OUT_12479_out0;
wire  [31:0] v$OUT_12481_out0;
wire  [31:0] v$OUT_3364_out0;
wire  [31:0] v$OUT_3365_out0;
wire  [31:0] v$SEL1_15425_out0;
wire  [31:0] v$SEL1_15431_out0;
wire  [31:0] v$SEL1_8734_out0;
wire  [31:0] v$SEL1_8740_out0;
wire  [31:0] v$SINGLE$PRECISION$32$BITS_13705_out0;
wire  [31:0] v$SINGLE$PRECISION_7900_out0;
wire  [31:0] v$SINGLE$PRECISION_7901_out0;
wire  [31:0] v$_12523_out0;
wire  [31:0] v$_12524_out0;
wire  [31:0] v$_15826_out0;
wire  [31:0] v$_15827_out0;
wire  [31:0] v$_16096_out0;
wire  [31:0] v$_16507_out0;
wire  [31:0] v$_16508_out0;
wire  [31:0] v$_16799_out0;
wire  [31:0] v$_16800_out0;
wire  [31:0] v$_17036_out0;
wire  [31:0] v$_17037_out0;
wire  [31:0] v$_18260_out0;
wire  [31:0] v$_18261_out0;
wire  [31:0] v$_18417_out0;
wire  [31:0] v$_18419_out0;
wire  [31:0] v$_1852_out0;
wire  [31:0] v$_1853_out0;
wire  [31:0] v$_5491_out0;
wire  [32:0] v$_12992_out0;
wire  [32:0] v$_9488_out0;
wire  [33:0] v$_15860_out0;
wire  [33:0] v$_16504_out0;
wire  [34:0] v$_16340_out0;
wire  [34:0] v$_1828_out0;
wire  [35:0] v$MULTIPLIER$TO$SAVE_16746_out0;
wire  [35:0] v$SAVED_14656_out0;
wire  [35:0] v$SAVED_15383_out0;
wire  [35:0] v$_13316_out0;
wire  [35:0] v$_1606_out0;
wire  [39:0] v$SEL1_15423_out0;
wire  [39:0] v$SEL1_15429_out0;
wire  [39:0] v$SEL1_8732_out0;
wire  [39:0] v$SEL1_8738_out0;
wire  [3:0] v$3_13396_out0;
wire  [3:0] v$3_13397_out0;
wire  [3:0] v$9_14315_out0;
wire  [3:0] v$9_14316_out0;
wire  [3:0] v$ADDRMSB_15028_out0;
wire  [3:0] v$ADDRMSB_15029_out0;
wire  [3:0] v$A_11316_out0;
wire  [3:0] v$A_11318_out0;
wire  [3:0] v$A_11319_out0;
wire  [3:0] v$A_11320_out0;
wire  [3:0] v$A_11322_out0;
wire  [3:0] v$A_11323_out0;
wire  [3:0] v$A_11326_out0;
wire  [3:0] v$A_11327_out0;
wire  [3:0] v$A_11330_out0;
wire  [3:0] v$A_11331_out0;
wire  [3:0] v$A_11334_out0;
wire  [3:0] v$A_11335_out0;
wire  [3:0] v$A_11336_out0;
wire  [3:0] v$A_11338_out0;
wire  [3:0] v$A_11339_out0;
wire  [3:0] v$A_11340_out0;
wire  [3:0] v$A_11342_out0;
wire  [3:0] v$A_11343_out0;
wire  [3:0] v$A_11346_out0;
wire  [3:0] v$A_11347_out0;
wire  [3:0] v$B_13212_out0;
wire  [3:0] v$B_13213_out0;
wire  [3:0] v$B_14424_out0;
wire  [3:0] v$B_14426_out0;
wire  [3:0] v$B_14427_out0;
wire  [3:0] v$B_14428_out0;
wire  [3:0] v$B_14430_out0;
wire  [3:0] v$B_14431_out0;
wire  [3:0] v$B_14434_out0;
wire  [3:0] v$B_14435_out0;
wire  [3:0] v$B_14438_out0;
wire  [3:0] v$B_14439_out0;
wire  [3:0] v$B_14442_out0;
wire  [3:0] v$B_14443_out0;
wire  [3:0] v$B_14444_out0;
wire  [3:0] v$B_14446_out0;
wire  [3:0] v$B_14447_out0;
wire  [3:0] v$B_14448_out0;
wire  [3:0] v$B_14450_out0;
wire  [3:0] v$B_14451_out0;
wire  [3:0] v$B_14454_out0;
wire  [3:0] v$B_14455_out0;
wire  [3:0] v$B_14623_out0;
wire  [3:0] v$B_14624_out0;
wire  [3:0] v$B_3704_out0;
wire  [3:0] v$B_3705_out0;
wire  [3:0] v$B_8316_out0;
wire  [3:0] v$B_8317_out0;
wire  [3:0] v$C0_204_out0;
wire  [3:0] v$C0_205_out0;
wire  [3:0] v$C12_3282_out0;
wire  [3:0] v$C12_3283_out0;
wire  [3:0] v$C1_12825_out0;
wire  [3:0] v$C1_12826_out0;
wire  [3:0] v$C1_5412_out0;
wire  [3:0] v$C1_5413_out0;
wire  [3:0] v$C1_5964_out0;
wire  [3:0] v$C1_5969_out0;
wire  [3:0] v$C1_5974_out0;
wire  [3:0] v$C1_5978_out0;
wire  [3:0] v$C1_5984_out0;
wire  [3:0] v$C1_5988_out0;
wire  [3:0] v$C1_5995_out0;
wire  [3:0] v$C1_6002_out0;
wire  [3:0] v$C1_6008_out0;
wire  [3:0] v$C1_6012_out0;
wire  [3:0] v$C1_6017_out0;
wire  [3:0] v$C1_6022_out0;
wire  [3:0] v$C1_7973_out0;
wire  [3:0] v$C1_7977_out0;
wire  [3:0] v$C2_106_out0;
wire  [3:0] v$C2_111_out0;
wire  [3:0] v$C2_116_out0;
wire  [3:0] v$C2_120_out0;
wire  [3:0] v$C2_126_out0;
wire  [3:0] v$C2_130_out0;
wire  [3:0] v$C2_137_out0;
wire  [3:0] v$C2_144_out0;
wire  [3:0] v$C2_150_out0;
wire  [3:0] v$C2_154_out0;
wire  [3:0] v$C2_159_out0;
wire  [3:0] v$C2_164_out0;
wire  [3:0] v$C4_10778_out0;
wire  [3:0] v$C4_10779_out0;
wire  [3:0] v$C8_7281_out0;
wire  [3:0] v$C8_7282_out0;
wire  [3:0] v$C8_8325_out0;
wire  [3:0] v$C8_8326_out0;
wire  [3:0] v$IN_15057_out0;
wire  [3:0] v$IN_15058_out0;
wire  [3:0] v$IN_15059_out0;
wire  [3:0] v$IN_15060_out0;
wire  [3:0] v$IN_15061_out0;
wire  [3:0] v$IN_15062_out0;
wire  [3:0] v$IN_15063_out0;
wire  [3:0] v$IN_15064_out0;
wire  [3:0] v$IN_15065_out0;
wire  [3:0] v$IN_15066_out0;
wire  [3:0] v$IN_15067_out0;
wire  [3:0] v$IN_15068_out0;
wire  [3:0] v$IN_15069_out0;
wire  [3:0] v$IN_15070_out0;
wire  [3:0] v$IN_15071_out0;
wire  [3:0] v$IN_15072_out0;
wire  [3:0] v$IN_15073_out0;
wire  [3:0] v$IN_15074_out0;
wire  [3:0] v$IN_15075_out0;
wire  [3:0] v$IN_15076_out0;
wire  [3:0] v$IN_15077_out0;
wire  [3:0] v$IN_15078_out0;
wire  [3:0] v$IN_15079_out0;
wire  [3:0] v$IN_15080_out0;
wire  [3:0] v$IN_15081_out0;
wire  [3:0] v$IN_15082_out0;
wire  [3:0] v$IN_15083_out0;
wire  [3:0] v$IN_15084_out0;
wire  [3:0] v$IN_15085_out0;
wire  [3:0] v$IN_15086_out0;
wire  [3:0] v$IN_15087_out0;
wire  [3:0] v$IN_15088_out0;
wire  [3:0] v$IN_15089_out0;
wire  [3:0] v$IN_15090_out0;
wire  [3:0] v$IN_15091_out0;
wire  [3:0] v$IN_15092_out0;
wire  [3:0] v$IN_15093_out0;
wire  [3:0] v$IN_15094_out0;
wire  [3:0] v$IN_15095_out0;
wire  [3:0] v$IN_15096_out0;
wire  [3:0] v$IN_15097_out0;
wire  [3:0] v$IN_15098_out0;
wire  [3:0] v$IN_15099_out0;
wire  [3:0] v$IN_15100_out0;
wire  [3:0] v$IN_15101_out0;
wire  [3:0] v$IN_15102_out0;
wire  [3:0] v$IN_15103_out0;
wire  [3:0] v$IN_15104_out0;
wire  [3:0] v$IR1$FULL$OP$CODE_17055_out0;
wire  [3:0] v$IR1$FULL$OP$CODE_17056_out0;
wire  [3:0] v$IR1$N_15765_out0;
wire  [3:0] v$IR1$N_15766_out0;
wire  [3:0] v$IR1$OPCODE_2895_out0;
wire  [3:0] v$IR1$OPCODE_2896_out0;
wire  [3:0] v$IR1$OPCODE_9564_out0;
wire  [3:0] v$IR1$OPCODE_9565_out0;
wire  [3:0] v$IR2$FULL$OP$CODE_11820_out0;
wire  [3:0] v$IR2$FULL$OP$CODE_11821_out0;
wire  [3:0] v$IR2$N_2984_out0;
wire  [3:0] v$IR2$N_2985_out0;
wire  [3:0] v$IR2$OPCODE_2569_out0;
wire  [3:0] v$IR2$OPCODE_2570_out0;
wire  [3:0] v$LSBS_15316_out0;
wire  [3:0] v$LSBS_15317_out0;
wire  [3:0] v$MUX3_17470_out0;
wire  [3:0] v$MUX3_17471_out0;
wire  [3:0] v$MUX3_17472_out0;
wire  [3:0] v$MUX3_17473_out0;
wire  [3:0] v$MUX3_17474_out0;
wire  [3:0] v$MUX3_17475_out0;
wire  [3:0] v$MUX3_17476_out0;
wire  [3:0] v$MUX3_17477_out0;
wire  [3:0] v$MUX4_2871_out0;
wire  [3:0] v$MUX4_2872_out0;
wire  [3:0] v$MUX4_2874_out0;
wire  [3:0] v$MUX4_2875_out0;
wire  [3:0] v$MUX4_2876_out0;
wire  [3:0] v$MUX4_2878_out0;
wire  [3:0] v$MUX4_2879_out0;
wire  [3:0] v$MUX4_2880_out0;
wire  [3:0] v$MUX5_14489_out0;
wire  [3:0] v$MUX5_14490_out0;
wire  [3:0] v$MUX5_4054_out0;
wire  [3:0] v$MUX5_4056_out0;
wire  [3:0] v$MUX5_4058_out0;
wire  [3:0] v$MUX5_4059_out0;
wire  [3:0] v$MUX5_4060_out0;
wire  [3:0] v$MUX5_4062_out0;
wire  [3:0] v$MUX5_4063_out0;
wire  [3:0] v$MUX5_4064_out0;
wire  [3:0] v$MUX6_2847_out0;
wire  [3:0] v$MUX6_2848_out0;
wire  [3:0] v$OPCODE_18050_out0;
wire  [3:0] v$OPCODE_18051_out0;
wire  [3:0] v$OP_10992_out0;
wire  [3:0] v$OP_10993_out0;
wire  [3:0] v$OP_14780_out0;
wire  [3:0] v$OP_14781_out0;
wire  [3:0] v$OP_17803_out0;
wire  [3:0] v$OP_17804_out0;
wire  [3:0] v$OP_3690_out0;
wire  [3:0] v$OP_3691_out0;
wire  [3:0] v$OP_5038_out0;
wire  [3:0] v$OP_5039_out0;
wire  [3:0] v$OUT_8952_out0;
wire  [3:0] v$OUT_8954_out0;
wire  [3:0] v$OUT_8956_out0;
wire  [3:0] v$OUT_8957_out0;
wire  [3:0] v$OUT_8958_out0;
wire  [3:0] v$OUT_8960_out0;
wire  [3:0] v$OUT_8961_out0;
wire  [3:0] v$OUT_8962_out0;
wire  [3:0] v$QP_18537_out0;
wire  [3:0] v$QP_18538_out0;
wire  [3:0] v$Q_12980_out0;
wire  [3:0] v$Q_12981_out0;
wire  [3:0] v$Q_6153_out0;
wire  [3:0] v$Q_6154_out0;
wire  [3:0] v$RXFSMQP_10030_out0;
wire  [3:0] v$RXFSMQP_10031_out0;
wire  [3:0] v$RXFSMQ_10814_out0;
wire  [3:0] v$RXFSMQ_10815_out0;
wire  [3:0] v$SEL12_12802_out0;
wire  [3:0] v$SEL12_12803_out0;
wire  [3:0] v$SEL1_10290_out0;
wire  [3:0] v$SEL1_10291_out0;
wire  [3:0] v$SEL1_10292_out0;
wire  [3:0] v$SEL1_10293_out0;
wire  [3:0] v$SEL1_10294_out0;
wire  [3:0] v$SEL1_10295_out0;
wire  [3:0] v$SEL1_10296_out0;
wire  [3:0] v$SEL1_10297_out0;
wire  [3:0] v$SEL1_16455_out0;
wire  [3:0] v$SEL1_16456_out0;
wire  [3:0] v$SEL1_16457_out0;
wire  [3:0] v$SEL1_16458_out0;
wire  [3:0] v$SEL1_16459_out0;
wire  [3:0] v$SEL1_16460_out0;
wire  [3:0] v$SEL1_16461_out0;
wire  [3:0] v$SEL1_16462_out0;
wire  [3:0] v$SEL1_16685_out0;
wire  [3:0] v$SEL1_16687_out0;
wire  [3:0] v$SEL1_16689_out0;
wire  [3:0] v$SEL1_16690_out0;
wire  [3:0] v$SEL1_16691_out0;
wire  [3:0] v$SEL1_16693_out0;
wire  [3:0] v$SEL1_16694_out0;
wire  [3:0] v$SEL1_16695_out0;
wire  [3:0] v$SEL1_18247_out0;
wire  [3:0] v$SEL1_18248_out0;
wire  [3:0] v$SEL1_8796_out0;
wire  [3:0] v$SEL1_8797_out0;
wire  [3:0] v$SEL2_13850_out0;
wire  [3:0] v$SEL2_13851_out0;
wire  [3:0] v$SEL2_13853_out0;
wire  [3:0] v$SEL2_13854_out0;
wire  [3:0] v$SEL2_13855_out0;
wire  [3:0] v$SEL2_13857_out0;
wire  [3:0] v$SEL2_13858_out0;
wire  [3:0] v$SEL2_13859_out0;
wire  [3:0] v$SEL2_17438_out0;
wire  [3:0] v$SEL2_17439_out0;
wire  [3:0] v$SEL2_17440_out0;
wire  [3:0] v$SEL2_17441_out0;
wire  [3:0] v$SEL2_17442_out0;
wire  [3:0] v$SEL2_17443_out0;
wire  [3:0] v$SEL2_17444_out0;
wire  [3:0] v$SEL2_17445_out0;
wire  [3:0] v$SEL2_2434_out0;
wire  [3:0] v$SEL2_2435_out0;
wire  [3:0] v$SEL2_3024_out0;
wire  [3:0] v$SEL2_3025_out0;
wire  [3:0] v$SEL2_3026_out0;
wire  [3:0] v$SEL2_3027_out0;
wire  [3:0] v$SEL2_3028_out0;
wire  [3:0] v$SEL2_3029_out0;
wire  [3:0] v$SEL2_3030_out0;
wire  [3:0] v$SEL2_3031_out0;
wire  [3:0] v$SEL3_16650_out0;
wire  [3:0] v$SEL3_16651_out0;
wire  [3:0] v$SEL3_18618_out0;
wire  [3:0] v$SEL3_18619_out0;
wire  [3:0] v$SEL3_18620_out0;
wire  [3:0] v$SEL3_18621_out0;
wire  [3:0] v$SEL3_7364_out0;
wire  [3:0] v$SEL3_7365_out0;
wire  [3:0] v$SEL3_7367_out0;
wire  [3:0] v$SEL3_7368_out0;
wire  [3:0] v$SEL3_7369_out0;
wire  [3:0] v$SEL3_7371_out0;
wire  [3:0] v$SEL3_7372_out0;
wire  [3:0] v$SEL3_7373_out0;
wire  [3:0] v$SEL3_9047_out0;
wire  [3:0] v$SEL3_9048_out0;
wire  [3:0] v$SEL3_9049_out0;
wire  [3:0] v$SEL3_9050_out0;
wire  [3:0] v$SEL3_9051_out0;
wire  [3:0] v$SEL3_9052_out0;
wire  [3:0] v$SEL3_9053_out0;
wire  [3:0] v$SEL3_9054_out0;
wire  [3:0] v$SEL4_17330_out0;
wire  [3:0] v$SEL4_17331_out0;
wire  [3:0] v$SEL4_17332_out0;
wire  [3:0] v$SEL4_17333_out0;
wire  [3:0] v$SEL4_17334_out0;
wire  [3:0] v$SEL4_17335_out0;
wire  [3:0] v$SEL4_17336_out0;
wire  [3:0] v$SEL4_17337_out0;
wire  [3:0] v$SEL4_3368_out0;
wire  [3:0] v$SEL4_3369_out0;
wire  [3:0] v$SEL4_3370_out0;
wire  [3:0] v$SEL4_3371_out0;
wire  [3:0] v$SEL4_3372_out0;
wire  [3:0] v$SEL4_3373_out0;
wire  [3:0] v$SEL4_3374_out0;
wire  [3:0] v$SEL4_3375_out0;
wire  [3:0] v$SEL4_9574_out0;
wire  [3:0] v$SEL4_9575_out0;
wire  [3:0] v$SEL4_9576_out0;
wire  [3:0] v$SEL4_9577_out0;
wire  [3:0] v$TXFSMQP_8772_out0;
wire  [3:0] v$TXFSMQP_8773_out0;
wire  [3:0] v$TXFSMQ_6207_out0;
wire  [3:0] v$TXFSMQ_6208_out0;
wire  [3:0] v$USELESS_15483_out0;
wire  [3:0] v$_10250_out0;
wire  [3:0] v$_10251_out0;
wire  [3:0] v$_10349_out0;
wire  [3:0] v$_10350_out0;
wire  [3:0] v$_10351_out0;
wire  [3:0] v$_10352_out0;
wire  [3:0] v$_10353_out0;
wire  [3:0] v$_10355_out0;
wire  [3:0] v$_10356_out0;
wire  [3:0] v$_10357_out0;
wire  [3:0] v$_10358_out0;
wire  [3:0] v$_10359_out0;
wire  [3:0] v$_1231_out0;
wire  [3:0] v$_1232_out0;
wire  [3:0] v$_1242_out0;
wire  [3:0] v$_1243_out0;
wire  [3:0] v$_1244_out0;
wire  [3:0] v$_1245_out0;
wire  [3:0] v$_1246_out0;
wire  [3:0] v$_12860_out0;
wire  [3:0] v$_12860_out1;
wire  [3:0] v$_12861_out0;
wire  [3:0] v$_12861_out1;
wire  [3:0] v$_12862_out0;
wire  [3:0] v$_12862_out1;
wire  [3:0] v$_12863_out0;
wire  [3:0] v$_12863_out1;
wire  [3:0] v$_12864_out0;
wire  [3:0] v$_12864_out1;
wire  [3:0] v$_12865_out0;
wire  [3:0] v$_12865_out1;
wire  [3:0] v$_12866_out0;
wire  [3:0] v$_12866_out1;
wire  [3:0] v$_12867_out0;
wire  [3:0] v$_12867_out1;
wire  [3:0] v$_12868_out0;
wire  [3:0] v$_12868_out1;
wire  [3:0] v$_12869_out0;
wire  [3:0] v$_12869_out1;
wire  [3:0] v$_12870_out0;
wire  [3:0] v$_12870_out1;
wire  [3:0] v$_12871_out0;
wire  [3:0] v$_12871_out1;
wire  [3:0] v$_12902_out0;
wire  [3:0] v$_12903_out0;
wire  [3:0] v$_13013_out0;
wire  [3:0] v$_13014_out0;
wire  [3:0] v$_13270_out0;
wire  [3:0] v$_13273_out0;
wire  [3:0] v$_13732_out0;
wire  [3:0] v$_13733_out0;
wire  [3:0] v$_13734_out0;
wire  [3:0] v$_13735_out0;
wire  [3:0] v$_13736_out0;
wire  [3:0] v$_14024_out1;
wire  [3:0] v$_14025_out1;
wire  [3:0] v$_14293_out0;
wire  [3:0] v$_14294_out0;
wire  [3:0] v$_14295_out0;
wire  [3:0] v$_14296_out0;
wire  [3:0] v$_14297_out0;
wire  [3:0] v$_1557_out0;
wire  [3:0] v$_1558_out0;
wire  [3:0] v$_1559_out0;
wire  [3:0] v$_1560_out0;
wire  [3:0] v$_1561_out0;
wire  [3:0] v$_16041_out0;
wire  [3:0] v$_16042_out0;
wire  [3:0] v$_16127_out0;
wire  [3:0] v$_16128_out0;
wire  [3:0] v$_16256_out0;
wire  [3:0] v$_16257_out0;
wire  [3:0] v$_16258_out0;
wire  [3:0] v$_16259_out0;
wire  [3:0] v$_16260_out0;
wire  [3:0] v$_16886_out0;
wire  [3:0] v$_16887_out0;
wire  [3:0] v$_17409_out0;
wire  [3:0] v$_17410_out0;
wire  [3:0] v$_17964_out0;
wire  [3:0] v$_17965_out0;
wire  [3:0] v$_17966_out0;
wire  [3:0] v$_17967_out0;
wire  [3:0] v$_17968_out0;
wire  [3:0] v$_18249_out0;
wire  [3:0] v$_18250_out0;
wire  [3:0] v$_18303_out0;
wire  [3:0] v$_18304_out0;
wire  [3:0] v$_18305_out0;
wire  [3:0] v$_18306_out0;
wire  [3:0] v$_18307_out0;
wire  [3:0] v$_1838_out0;
wire  [3:0] v$_1839_out0;
wire  [3:0] v$_18459_out0;
wire  [3:0] v$_18459_out1;
wire  [3:0] v$_18460_out0;
wire  [3:0] v$_18460_out1;
wire  [3:0] v$_18607_out0;
wire  [3:0] v$_18608_out0;
wire  [3:0] v$_2345_out0;
wire  [3:0] v$_2345_out1;
wire  [3:0] v$_2346_out0;
wire  [3:0] v$_2346_out1;
wire  [3:0] v$_258_out0;
wire  [3:0] v$_259_out0;
wire  [3:0] v$_2897_out0;
wire  [3:0] v$_2897_out1;
wire  [3:0] v$_2898_out0;
wire  [3:0] v$_2898_out1;
wire  [3:0] v$_304_out0;
wire  [3:0] v$_305_out0;
wire  [3:0] v$_3706_out0;
wire  [3:0] v$_3707_out0;
wire  [3:0] v$_3799_out0;
wire  [3:0] v$_3800_out0;
wire  [3:0] v$_3977_out0;
wire  [3:0] v$_3978_out0;
wire  [3:0] v$_3979_out0;
wire  [3:0] v$_3980_out0;
wire  [3:0] v$_3981_out0;
wire  [3:0] v$_3982_out0;
wire  [3:0] v$_3983_out0;
wire  [3:0] v$_3984_out0;
wire  [3:0] v$_4164_out0;
wire  [3:0] v$_4165_out0;
wire  [3:0] v$_5090_out0;
wire  [3:0] v$_5092_out0;
wire  [3:0] v$_5094_out0;
wire  [3:0] v$_5095_out0;
wire  [3:0] v$_5096_out0;
wire  [3:0] v$_5098_out0;
wire  [3:0] v$_5099_out0;
wire  [3:0] v$_5100_out0;
wire  [3:0] v$_5232_out0;
wire  [3:0] v$_5233_out0;
wire  [3:0] v$_5474_out0;
wire  [3:0] v$_5475_out0;
wire  [3:0] v$_5517_out0;
wire  [3:0] v$_5518_out0;
wire  [3:0] v$_6343_out0;
wire  [3:0] v$_6344_out0;
wire  [3:0] v$_6461_out0;
wire  [3:0] v$_6461_out1;
wire  [3:0] v$_6462_out0;
wire  [3:0] v$_6462_out1;
wire  [3:0] v$_683_out0;
wire  [3:0] v$_684_out0;
wire  [3:0] v$_6990_out0;
wire  [3:0] v$_6991_out0;
wire  [3:0] v$_7023_out0;
wire  [3:0] v$_7024_out0;
wire  [3:0] v$_7253_out0;
wire  [3:0] v$_7254_out0;
wire  [3:0] v$_7255_out0;
wire  [3:0] v$_7256_out0;
wire  [3:0] v$_7257_out0;
wire  [3:0] v$_7277_out0;
wire  [3:0] v$_7378_out0;
wire  [3:0] v$_7379_out0;
wire  [3:0] v$_7404_out0;
wire  [3:0] v$_7405_out0;
wire  [3:0] v$_7406_out0;
wire  [3:0] v$_7407_out0;
wire  [3:0] v$_7408_out0;
wire  [3:0] v$_7550_out0;
wire  [3:0] v$_7551_out0;
wire  [3:0] v$_8213_out0;
wire  [3:0] v$_8213_out1;
wire  [3:0] v$_8214_out0;
wire  [3:0] v$_8214_out1;
wire  [3:0] v$_8408_out0;
wire  [3:0] v$_8408_out1;
wire  [3:0] v$_8409_out0;
wire  [3:0] v$_8409_out1;
wire  [3:0] v$_8691_out0;
wire  [3:0] v$_8692_out0;
wire  [3:0] v$_8781_out0;
wire  [3:0] v$_8783_out0;
wire  [3:0] v$_8785_out0;
wire  [3:0] v$_8786_out0;
wire  [3:0] v$_8787_out0;
wire  [3:0] v$_8789_out0;
wire  [3:0] v$_8790_out0;
wire  [3:0] v$_8791_out0;
wire  [3:0] v$_8896_out0;
wire  [3:0] v$_8897_out0;
wire  [3:0] v$_8899_out0;
wire  [3:0] v$_8900_out0;
wire  [3:0] v$_8901_out0;
wire  [3:0] v$_8903_out0;
wire  [3:0] v$_8904_out0;
wire  [3:0] v$_8905_out0;
wire  [3:0] v$_8935_out0;
wire  [3:0] v$_8936_out0;
wire  [3:0] v$_9432_out0;
wire  [3:0] v$_9433_out0;
wire  [3:0] v$_9491_out0;
wire  [3:0] v$_9492_out0;
wire  [3:0] v$_9493_out0;
wire  [3:0] v$_9494_out0;
wire  [3:0] v$_9495_out0;
wire  [43:0] v$AROM1_16158_out0;
wire  [43:0] v$AROM1_16159_out0;
wire  [43:0] v$SEL1_15427_out0;
wire  [43:0] v$SEL1_15433_out0;
wire  [43:0] v$SEL1_8736_out0;
wire  [43:0] v$SEL1_8742_out0;
wire  [45:0] v$SEL1_15424_out0;
wire  [45:0] v$SEL1_15430_out0;
wire  [45:0] v$SEL1_8733_out0;
wire  [45:0] v$SEL1_8739_out0;
wire  [46:0] v$SEL1_15426_out0;
wire  [46:0] v$SEL1_15432_out0;
wire  [46:0] v$SEL1_8735_out0;
wire  [46:0] v$SEL1_8741_out0;
wire  [47:0] v$IN_11073_out0;
wire  [47:0] v$IN_11074_out0;
wire  [47:0] v$IN_11644_out0;
wire  [47:0] v$IN_11645_out0;
wire  [47:0] v$IN_11788_out0;
wire  [47:0] v$IN_11789_out0;
wire  [47:0] v$IN_13566_out0;
wire  [47:0] v$IN_13570_out0;
wire  [47:0] v$IN_15610_out0;
wire  [47:0] v$IN_15611_out0;
wire  [47:0] v$IN_18264_out0;
wire  [47:0] v$IN_18265_out0;
wire  [47:0] v$IN_3866_out0;
wire  [47:0] v$IN_3867_out0;
wire  [47:0] v$IN_3868_out0;
wire  [47:0] v$IN_3869_out0;
wire  [47:0] v$IN_3870_out0;
wire  [47:0] v$IN_3871_out0;
wire  [47:0] v$IN_4192_out0;
wire  [47:0] v$IN_4193_out0;
wire  [47:0] v$IN_5030_out0;
wire  [47:0] v$IN_5031_out0;
wire  [47:0] v$IN_5183_out0;
wire  [47:0] v$IN_5184_out0;
wire  [47:0] v$IN_5185_out0;
wire  [47:0] v$IN_5186_out0;
wire  [47:0] v$IN_5187_out0;
wire  [47:0] v$IN_5188_out0;
wire  [47:0] v$IN_5189_out0;
wire  [47:0] v$IN_5190_out0;
wire  [47:0] v$IN_5191_out0;
wire  [47:0] v$IN_5192_out0;
wire  [47:0] v$IN_5193_out0;
wire  [47:0] v$IN_5194_out0;
wire  [47:0] v$IN_8296_out0;
wire  [47:0] v$IN_8297_out0;
wire  [47:0] v$MULTIPLIER$OUT_5788_out0;
wire  [47:0] v$MULTIPLIER$OUT_9344_out0;
wire  [47:0] v$MUX1_2385_out0;
wire  [47:0] v$MUX1_2386_out0;
wire  [47:0] v$MUX1_2387_out0;
wire  [47:0] v$MUX1_2388_out0;
wire  [47:0] v$MUX1_2389_out0;
wire  [47:0] v$MUX1_2390_out0;
wire  [47:0] v$MUX1_2391_out0;
wire  [47:0] v$MUX1_2392_out0;
wire  [47:0] v$MUX1_2393_out0;
wire  [47:0] v$MUX1_2394_out0;
wire  [47:0] v$MUX1_2395_out0;
wire  [47:0] v$MUX1_2396_out0;
wire  [47:0] v$MUX2_15241_out0;
wire  [47:0] v$MUX2_15242_out0;
wire  [47:0] v$MUX2_18580_out0;
wire  [47:0] v$MUX2_18581_out0;
wire  [47:0] v$MUX2_18582_out0;
wire  [47:0] v$MUX2_18583_out0;
wire  [47:0] v$MUX2_18584_out0;
wire  [47:0] v$MUX2_18585_out0;
wire  [47:0] v$MUX2_2482_out0;
wire  [47:0] v$MUX2_2483_out0;
wire  [47:0] v$MUX2_2504_out0;
wire  [47:0] v$MUX2_2505_out0;
wire  [47:0] v$OUT_14937_out0;
wire  [47:0] v$OUT_14938_out0;
wire  [47:0] v$OUT_14939_out0;
wire  [47:0] v$OUT_14940_out0;
wire  [47:0] v$OUT_14941_out0;
wire  [47:0] v$OUT_14942_out0;
wire  [47:0] v$OUT_14943_out0;
wire  [47:0] v$OUT_14944_out0;
wire  [47:0] v$OUT_14945_out0;
wire  [47:0] v$OUT_14946_out0;
wire  [47:0] v$OUT_14947_out0;
wire  [47:0] v$OUT_14948_out0;
wire  [47:0] v$OUT_4915_out0;
wire  [47:0] v$OUT_4916_out0;
wire  [47:0] v$OUT_8212_out0;
wire  [47:0] v$_2533_out0;
wire  [47:0] v$_4281_out0;
wire  [47:0] v$_4282_out0;
wire  [47:0] v$_4283_out0;
wire  [47:0] v$_4284_out0;
wire  [47:0] v$_4285_out0;
wire  [47:0] v$_4286_out0;
wire  [47:0] v$_4287_out0;
wire  [47:0] v$_4288_out0;
wire  [47:0] v$_4289_out0;
wire  [47:0] v$_4290_out0;
wire  [47:0] v$_4291_out0;
wire  [47:0] v$_4292_out0;
wire  [47:0] v$_9016_out0;
wire  [47:0] v$_9017_out0;
wire  [47:0] v$_9018_out0;
wire  [47:0] v$_9019_out0;
wire  [47:0] v$_9020_out0;
wire  [47:0] v$_9021_out0;
wire  [47:0] v$_9022_out0;
wire  [47:0] v$_9023_out0;
wire  [47:0] v$_9024_out0;
wire  [47:0] v$_9025_out0;
wire  [47:0] v$_9026_out0;
wire  [47:0] v$_9027_out0;
wire  [4:0] v$A$EXP_284_out0;
wire  [4:0] v$A$EXP_286_out0;
wire  [4:0] v$A$EXP_288_out0;
wire  [4:0] v$A$EXP_290_out0;
wire  [4:0] v$A1_11802_out0;
wire  [4:0] v$A1_11803_out0;
wire  [4:0] v$A1_2662_out0;
wire  [4:0] v$A1_2664_out0;
wire  [4:0] v$A1_2938_out0;
wire  [4:0] v$A1_5789_out0;
wire  [4:0] v$A1_5791_out0;
wire  [4:0] v$A1_5793_out0;
wire  [4:0] v$A1_5795_out0;
wire  [4:0] v$A1_7730_out0;
wire  [4:0] v$A1_7731_out0;
wire  [4:0] v$A2_10044_out0;
wire  [4:0] v$A2_10046_out0;
wire  [4:0] v$AMOUNT$OF$SHIFT_9459_out0;
wire  [4:0] v$AMOUNT$OF$SHIFT_9460_out0;
wire  [4:0] v$A_11324_out0;
wire  [4:0] v$A_11328_out0;
wire  [4:0] v$A_11332_out0;
wire  [4:0] v$A_11344_out0;
wire  [4:0] v$B$EXP_16672_out0;
wire  [4:0] v$B$EXP_16674_out0;
wire  [4:0] v$B$EXP_16676_out0;
wire  [4:0] v$B$EXP_16678_out0;
wire  [4:0] v$B_14432_out0;
wire  [4:0] v$B_14436_out0;
wire  [4:0] v$B_14440_out0;
wire  [4:0] v$B_14452_out0;
wire  [4:0] v$C1_13574_out0;
wire  [4:0] v$C1_13576_out0;
wire  [4:0] v$C1_13578_out0;
wire  [4:0] v$C1_13580_out0;
wire  [4:0] v$C1_15678_out0;
wire  [4:0] v$C1_15734_out0;
wire  [4:0] v$C1_15735_out0;
wire  [4:0] v$C1_5239_out0;
wire  [4:0] v$C1_5955_out0;
wire  [4:0] v$C1_5957_out0;
wire  [4:0] v$C1_7424_out0;
wire  [4:0] v$C1_7425_out0;
wire  [4:0] v$C3_7014_out0;
wire  [4:0] v$C4_14657_out0;
wire  [4:0] v$DIFF_9087_out0;
wire  [4:0] v$DIFF_9089_out0;
wire  [4:0] v$DIFF_9091_out0;
wire  [4:0] v$DIFF_9093_out0;
wire  [4:0] v$D_5727_out0;
wire  [4:0] v$EXPONENT_16011_out0;
wire  [4:0] v$EXPONENT_16012_out0;
wire  [4:0] v$EXPONENT_16395_out0;
wire  [4:0] v$EXPONENT_16396_out0;
wire  [4:0] v$EXPONENT_18076_out0;
wire  [4:0] v$EXPONENT_18077_out0;
wire  [4:0] v$HALF$PRECISION$EXPONENT$DENORM_6129_out0;
wire  [4:0] v$HALF$PRECISION$EXPONENT$DENORM_6130_out0;
wire  [4:0] v$HALF$PRECISION$EXPONENT_14671_out0;
wire  [4:0] v$HALF$PRECISION$EXPONENT_14672_out0;
wire  [4:0] v$HALF$PRECISION$EXPONENT_6382_out0;
wire  [4:0] v$HALF$PRECISION$EXPONENT_6383_out0;
wire  [4:0] v$HALF$PRECISSION$ADDITION$IN_1147_out0;
wire  [4:0] v$HALF$PRECISSION$ADDITION$IN_1148_out0;
wire  [4:0] v$K_301_out0;
wire  [4:0] v$K_302_out0;
wire  [4:0] v$LARGER$EXP_10274_out0;
wire  [4:0] v$LARGER$EXP_10276_out0;
wire  [4:0] v$MUX1_15287_out0;
wire  [4:0] v$MUX1_15288_out0;
wire  [4:0] v$MUX1_17923_out0;
wire  [4:0] v$MUX1_17925_out0;
wire  [4:0] v$MUX1_17927_out0;
wire  [4:0] v$MUX1_17929_out0;
wire  [4:0] v$MUX1_18598_out0;
wire  [4:0] v$MUX1_5137_out0;
wire  [4:0] v$MUX2_13544_out0;
wire  [4:0] v$MUX2_13545_out0;
wire  [4:0] v$MUX3_3391_out0;
wire  [4:0] v$MUX3_3393_out0;
wire  [4:0] v$MUX3_3395_out0;
wire  [4:0] v$MUX3_3397_out0;
wire  [4:0] v$MUX5_4053_out0;
wire  [4:0] v$MUX5_4055_out0;
wire  [4:0] v$NORMALIZATION$SHIFT_1824_out0;
wire  [4:0] v$NORMALIZATION$SHIFT_1825_out0;
wire  [4:0] v$NORMALIZATION$SHIFT_4397_out0;
wire  [4:0] v$NORMALIZATION$SHIFT_4398_out0;
wire  [4:0] v$N_16246_out0;
wire  [4:0] v$N_16247_out0;
wire  [4:0] v$N_16248_out0;
wire  [4:0] v$N_16249_out0;
wire  [4:0] v$OUT_170_out0;
wire  [4:0] v$OUT_171_out0;
wire  [4:0] v$OUT_5002_out0;
wire  [4:0] v$OUT_6193_out0;
wire  [4:0] v$OUT_6194_out0;
wire  [4:0] v$OUT_8923_out0;
wire  [4:0] v$OUT_8924_out0;
wire  [4:0] v$OUT_8951_out0;
wire  [4:0] v$OUT_8953_out0;
wire  [4:0] v$SEL10_3010_out0;
wire  [4:0] v$SEL10_3011_out0;
wire  [4:0] v$SEL14_9100_out0;
wire  [4:0] v$SEL14_9101_out0;
wire  [4:0] v$SEL18_18251_out0;
wire  [4:0] v$SEL18_18252_out0;
wire  [4:0] v$SEL1_7529_out0;
wire  [4:0] v$SEL1_7531_out0;
wire  [4:0] v$SEL1_7533_out0;
wire  [4:0] v$SEL1_7535_out0;
wire  [4:0] v$SEL1_9465_out0;
wire  [4:0] v$SEL1_9466_out0;
wire  [4:0] v$SEL25_13454_out0;
wire  [4:0] v$SEL25_13455_out0;
wire  [4:0] v$SEL25_13456_out0;
wire  [4:0] v$SEL25_13457_out0;
wire  [4:0] v$SEL2_6968_out0;
wire  [4:0] v$SEL2_6970_out0;
wire  [4:0] v$SEL2_6972_out0;
wire  [4:0] v$SEL2_6974_out0;
wire  [4:0] v$SEL9_3773_out0;
wire  [4:0] v$SEL9_3774_out0;
wire  [4:0] v$SMALLER$EXP_2941_out0;
wire  [4:0] v$SMALLER$EXP_2943_out0;
wire  [4:0] v$XOR1_10930_out0;
wire  [4:0] v$XOR1_10931_out0;
wire  [4:0] v$XOR1_3954_out0;
wire  [4:0] v$XOR1_7589_out0;
wire  [4:0] v$XOR1_7591_out0;
wire  [4:0] v$XOR1_7593_out0;
wire  [4:0] v$XOR1_7595_out0;
wire  [4:0] v$_1325_out0;
wire  [4:0] v$_1326_out0;
wire  [4:0] v$_2675_out0;
wire  [4:0] v$_2676_out0;
wire  [4:0] v$_3328_out0;
wire  [4:0] v$_3329_out0;
wire  [4:0] v$_5089_out0;
wire  [4:0] v$_5091_out0;
wire  [4:0] v$_6341_out0;
wire  [4:0] v$_6342_out0;
wire  [4:0] v$_7273_out0;
wire  [4:0] v$_7274_out0;
wire  [4:0] v$_8780_out0;
wire  [4:0] v$_8782_out0;
wire  [5:0] v$A1_4011_out0;
wire  [5:0] v$A1_4012_out0;
wire  [5:0] v$A2_14825_out0;
wire  [5:0] v$A2_14826_out0;
wire  [5:0] v$ADDRESS_14580_out0;
wire  [5:0] v$ADDRESS_14581_out0;
wire  [5:0] v$AMOUNT$OF$SHIFT_9461_out0;
wire  [5:0] v$AMOUNT$OF$SHIFT_9462_out0;
wire  [5:0] v$C2_15986_out0;
wire  [5:0] v$C2_15987_out0;
wire  [5:0] v$C3_13163_out0;
wire  [5:0] v$C3_13164_out0;
wire  [5:0] v$C6_8046_out0;
wire  [5:0] v$C6_8047_out0;
wire  [5:0] v$MUX1_9915_out0;
wire  [5:0] v$MUX1_9916_out0;
wire  [5:0] v$MUX4_2873_out0;
wire  [5:0] v$MUX4_2877_out0;
wire  [5:0] v$MUX5_4057_out0;
wire  [5:0] v$MUX5_4061_out0;
wire  [5:0] v$OUT_8955_out0;
wire  [5:0] v$OUT_8959_out0;
wire  [5:0] v$_1218_out0;
wire  [5:0] v$_1218_out1;
wire  [5:0] v$_1219_out0;
wire  [5:0] v$_1219_out1;
wire  [5:0] v$_1220_out0;
wire  [5:0] v$_1220_out1;
wire  [5:0] v$_1221_out0;
wire  [5:0] v$_1221_out1;
wire  [5:0] v$_1222_out0;
wire  [5:0] v$_1222_out1;
wire  [5:0] v$_1523_out0;
wire  [5:0] v$_1523_out1;
wire  [5:0] v$_1524_out0;
wire  [5:0] v$_1524_out1;
wire  [5:0] v$_1525_out0;
wire  [5:0] v$_1525_out1;
wire  [5:0] v$_1526_out0;
wire  [5:0] v$_1526_out1;
wire  [5:0] v$_1527_out0;
wire  [5:0] v$_1527_out1;
wire  [5:0] v$_16111_out0;
wire  [5:0] v$_16111_out1;
wire  [5:0] v$_16112_out0;
wire  [5:0] v$_16112_out1;
wire  [5:0] v$_16113_out0;
wire  [5:0] v$_16113_out1;
wire  [5:0] v$_16114_out0;
wire  [5:0] v$_16114_out1;
wire  [5:0] v$_16115_out0;
wire  [5:0] v$_16115_out1;
wire  [5:0] v$_17028_out0;
wire  [5:0] v$_17028_out1;
wire  [5:0] v$_17029_out0;
wire  [5:0] v$_17029_out1;
wire  [5:0] v$_17030_out0;
wire  [5:0] v$_17030_out1;
wire  [5:0] v$_17031_out0;
wire  [5:0] v$_17031_out1;
wire  [5:0] v$_17032_out0;
wire  [5:0] v$_17032_out1;
wire  [5:0] v$_5093_out0;
wire  [5:0] v$_5097_out0;
wire  [5:0] v$_8784_out0;
wire  [5:0] v$_8788_out0;
wire  [5:0] v$_8898_out0;
wire  [5:0] v$_8902_out0;
wire  [7:0] v$8LSB_7606_out0;
wire  [7:0] v$8LSB_7607_out0;
wire  [7:0] v$A$EXP_285_out0;
wire  [7:0] v$A$EXP_287_out0;
wire  [7:0] v$A$EXP_289_out0;
wire  [7:0] v$A$EXP_291_out0;
wire  [7:0] v$A1_15763_out0;
wire  [7:0] v$A1_15764_out0;
wire  [7:0] v$A1_2663_out0;
wire  [7:0] v$A1_2665_out0;
wire  [7:0] v$A1_5790_out0;
wire  [7:0] v$A1_5792_out0;
wire  [7:0] v$A1_5794_out0;
wire  [7:0] v$A1_5796_out0;
wire  [7:0] v$A1_638_out0;
wire  [7:0] v$A1_639_out0;
wire  [7:0] v$A2_10045_out0;
wire  [7:0] v$A2_10047_out0;
wire  [7:0] v$A_11317_out0;
wire  [7:0] v$A_11321_out0;
wire  [7:0] v$A_11325_out0;
wire  [7:0] v$A_11329_out0;
wire  [7:0] v$A_11333_out0;
wire  [7:0] v$A_11337_out0;
wire  [7:0] v$A_11341_out0;
wire  [7:0] v$A_11345_out0;
wire  [7:0] v$B$EXP_16673_out0;
wire  [7:0] v$B$EXP_16675_out0;
wire  [7:0] v$B$EXP_16677_out0;
wire  [7:0] v$B$EXP_16679_out0;
wire  [7:0] v$B_14425_out0;
wire  [7:0] v$B_14429_out0;
wire  [7:0] v$B_14433_out0;
wire  [7:0] v$B_14437_out0;
wire  [7:0] v$B_14441_out0;
wire  [7:0] v$B_14445_out0;
wire  [7:0] v$B_14449_out0;
wire  [7:0] v$B_14453_out0;
wire  [7:0] v$C1_13448_out0;
wire  [7:0] v$C1_13449_out0;
wire  [7:0] v$C1_13575_out0;
wire  [7:0] v$C1_13577_out0;
wire  [7:0] v$C1_13579_out0;
wire  [7:0] v$C1_13581_out0;
wire  [7:0] v$C1_13991_out0;
wire  [7:0] v$C1_13992_out0;
wire  [7:0] v$C1_14812_out0;
wire  [7:0] v$C1_14813_out0;
wire  [7:0] v$C1_1555_out0;
wire  [7:0] v$C1_1556_out0;
wire  [7:0] v$C1_5956_out0;
wire  [7:0] v$C1_5958_out0;
wire  [7:0] v$C1_5962_out0;
wire  [7:0] v$C1_5967_out0;
wire  [7:0] v$C1_5972_out0;
wire  [7:0] v$C1_5977_out0;
wire  [7:0] v$C1_5982_out0;
wire  [7:0] v$C1_5987_out0;
wire  [7:0] v$C1_5993_out0;
wire  [7:0] v$C1_5998_out0;
wire  [7:0] v$C1_6004_out0;
wire  [7:0] v$C1_6010_out0;
wire  [7:0] v$C1_6015_out0;
wire  [7:0] v$C1_6020_out0;
wire  [7:0] v$C1_7974_out0;
wire  [7:0] v$C1_7978_out0;
wire  [7:0] v$C2_104_out0;
wire  [7:0] v$C2_109_out0;
wire  [7:0] v$C2_114_out0;
wire  [7:0] v$C2_119_out0;
wire  [7:0] v$C2_124_out0;
wire  [7:0] v$C2_129_out0;
wire  [7:0] v$C2_135_out0;
wire  [7:0] v$C2_140_out0;
wire  [7:0] v$C2_146_out0;
wire  [7:0] v$C2_152_out0;
wire  [7:0] v$C2_157_out0;
wire  [7:0] v$C2_162_out0;
wire  [7:0] v$DIFF$VIEW$MANTISA$ADDER_12723_out0;
wire  [7:0] v$DIFF$VIEW$MANTISA$ADDER_12724_out0;
wire  [7:0] v$DIFF_12660_out0;
wire  [7:0] v$DIFF_12661_out0;
wire  [7:0] v$DIFF_15930_out0;
wire  [7:0] v$DIFF_15931_out0;
wire  [7:0] v$DIFF_17503_out0;
wire  [7:0] v$DIFF_17504_out0;
wire  [7:0] v$DIFF_17505_out0;
wire  [7:0] v$DIFF_17506_out0;
wire  [7:0] v$DIFF_2820_out0;
wire  [7:0] v$DIFF_2821_out0;
wire  [7:0] v$DIFF_292_out0;
wire  [7:0] v$DIFF_293_out0;
wire  [7:0] v$DIFF_9088_out0;
wire  [7:0] v$DIFF_9090_out0;
wire  [7:0] v$DIFF_9092_out0;
wire  [7:0] v$DIFF_9094_out0;
wire  [7:0] v$EDGEMODE_2886_out0;
wire  [7:0] v$EDGEMODE_2887_out0;
wire  [7:0] v$END_12712_out0;
wire  [7:0] v$END_12713_out0;
wire  [7:0] v$EXP$DIFF_12470_out0;
wire  [7:0] v$EXP$DIFF_12471_out0;
wire  [7:0] v$EXP$DIFF_13788_out0;
wire  [7:0] v$EXP$DIFF_13789_out0;
wire  [7:0] v$EXP$DIFF_14330_out0;
wire  [7:0] v$EXP$DIFF_14331_out0;
wire  [7:0] v$EXP$DIFF_17679_out0;
wire  [7:0] v$EXP$DIFF_17680_out0;
wire  [7:0] v$EXPONENT_1358_out0;
wire  [7:0] v$EXPONENT_1359_out0;
wire  [7:0] v$EXPONENT_13686_out0;
wire  [7:0] v$EXPONENT_13687_out0;
wire  [7:0] v$IN_14854_out0;
wire  [7:0] v$IN_14855_out0;
wire  [7:0] v$IN_14856_out0;
wire  [7:0] v$IN_14857_out0;
wire  [7:0] v$IN_14858_out0;
wire  [7:0] v$IN_14859_out0;
wire  [7:0] v$IN_14860_out0;
wire  [7:0] v$IN_14861_out0;
wire  [7:0] v$LARGER$EXP_10275_out0;
wire  [7:0] v$LARGER$EXP_10277_out0;
wire  [7:0] v$LSBS_7937_out0;
wire  [7:0] v$LSBS_7938_out0;
wire  [7:0] v$MODEIN_5780_out0;
wire  [7:0] v$MODEIN_5781_out0;
wire  [7:0] v$MODE_10801_out0;
wire  [7:0] v$MODE_10802_out0;
wire  [7:0] v$MODE_17842_out0;
wire  [7:0] v$MODE_17843_out0;
wire  [7:0] v$MODE_48_out0;
wire  [7:0] v$MODE_49_out0;
wire  [7:0] v$MUX13_10363_out0;
wire  [7:0] v$MUX13_10364_out0;
wire  [7:0] v$MUX1_17924_out0;
wire  [7:0] v$MUX1_17926_out0;
wire  [7:0] v$MUX1_17928_out0;
wire  [7:0] v$MUX1_17930_out0;
wire  [7:0] v$MUX2_17760_out0;
wire  [7:0] v$MUX2_17761_out0;
wire  [7:0] v$MUX3_3392_out0;
wire  [7:0] v$MUX3_3394_out0;
wire  [7:0] v$MUX3_3396_out0;
wire  [7:0] v$MUX3_3398_out0;
wire  [7:0] v$MUX5_13175_out0;
wire  [7:0] v$MUX5_13176_out0;
wire  [7:0] v$MUX6_13706_out0;
wire  [7:0] v$MUX6_13707_out0;
wire  [7:0] v$MUX6_7948_out0;
wire  [7:0] v$MUX6_7949_out0;
wire  [7:0] v$NORMALIZATION$SHIFT$WHOLE_6672_out0;
wire  [7:0] v$NORMALIZATION$SHIFT$WHOLE_6673_out0;
wire  [7:0] v$NORMALIZATION$SHIFT_10742_out0;
wire  [7:0] v$NORMALIZATION$SHIFT_10743_out0;
wire  [7:0] v$NORMALIZATION$SHIFT_1165_out0;
wire  [7:0] v$NORMALIZATION$SHIFT_1166_out0;
wire  [7:0] v$NORMALIZATION$SHIFT_18622_out0;
wire  [7:0] v$NORMALIZATION$SHIFT_18623_out0;
wire  [7:0] v$NORMALIZATION$SHIFT_3253_out0;
wire  [7:0] v$NORMALIZATION$SHIFT_3254_out0;
wire  [7:0] v$N_14070_out0;
wire  [7:0] v$N_14071_out0;
wire  [7:0] v$N_14072_out0;
wire  [7:0] v$N_14073_out0;
wire  [7:0] v$OUT_14778_out0;
wire  [7:0] v$OUT_14779_out0;
wire  [7:0] v$OUT_16097_out0;
wire  [7:0] v$OUT_16098_out0;
wire  [7:0] v$PIN_6634_out0;
wire  [7:0] v$PIN_6635_out0;
wire  [7:0] v$PIN_6636_out0;
wire  [7:0] v$PIN_6637_out0;
wire  [7:0] v$PIN_6638_out0;
wire  [7:0] v$PIN_6639_out0;
wire  [7:0] v$PIN_6640_out0;
wire  [7:0] v$PIN_6641_out0;
wire  [7:0] v$PIN_6642_out0;
wire  [7:0] v$PIN_6643_out0;
wire  [7:0] v$PIN_6644_out0;
wire  [7:0] v$PIN_6645_out0;
wire  [7:0] v$POUT_10361_out0;
wire  [7:0] v$POUT_10362_out0;
wire  [7:0] v$POut_13688_out0;
wire  [7:0] v$POut_13689_out0;
wire  [7:0] v$RXBYTE_18390_out0;
wire  [7:0] v$RXBYTE_18391_out0;
wire  [7:0] v$RXBYTE_9628_out0;
wire  [7:0] v$RXBYTE_9629_out0;
wire  [7:0] v$SEL17_5388_out0;
wire  [7:0] v$SEL17_5389_out0;
wire  [7:0] v$SEL1_15386_out0;
wire  [7:0] v$SEL1_15391_out0;
wire  [7:0] v$SEL1_15396_out0;
wire  [7:0] v$SEL1_15404_out0;
wire  [7:0] v$SEL1_15406_out0;
wire  [7:0] v$SEL1_15414_out0;
wire  [7:0] v$SEL1_15417_out0;
wire  [7:0] v$SEL1_15434_out0;
wire  [7:0] v$SEL1_15439_out0;
wire  [7:0] v$SEL1_15444_out0;
wire  [7:0] v$SEL1_16684_out0;
wire  [7:0] v$SEL1_16686_out0;
wire  [7:0] v$SEL1_17423_out0;
wire  [7:0] v$SEL1_17424_out0;
wire  [7:0] v$SEL1_351_out0;
wire  [7:0] v$SEL1_352_out0;
wire  [7:0] v$SEL1_7530_out0;
wire  [7:0] v$SEL1_7532_out0;
wire  [7:0] v$SEL1_7534_out0;
wire  [7:0] v$SEL1_7536_out0;
wire  [7:0] v$SEL1_8083_out0;
wire  [7:0] v$SEL1_8084_out0;
wire  [7:0] v$SEL1_8085_out0;
wire  [7:0] v$SEL1_8086_out0;
wire  [7:0] v$SEL1_8695_out0;
wire  [7:0] v$SEL1_8700_out0;
wire  [7:0] v$SEL1_8705_out0;
wire  [7:0] v$SEL1_8713_out0;
wire  [7:0] v$SEL1_8715_out0;
wire  [7:0] v$SEL1_8723_out0;
wire  [7:0] v$SEL1_8726_out0;
wire  [7:0] v$SEL1_8743_out0;
wire  [7:0] v$SEL1_8748_out0;
wire  [7:0] v$SEL1_8753_out0;
wire  [7:0] v$SEL2_17370_out0;
wire  [7:0] v$SEL2_17371_out0;
wire  [7:0] v$SEL2_17517_out0;
wire  [7:0] v$SEL2_17518_out0;
wire  [7:0] v$SEL2_17519_out0;
wire  [7:0] v$SEL2_17520_out0;
wire  [7:0] v$SEL2_6969_out0;
wire  [7:0] v$SEL2_6971_out0;
wire  [7:0] v$SEL2_6973_out0;
wire  [7:0] v$SEL2_6975_out0;
wire  [7:0] v$SEL3_17773_out0;
wire  [7:0] v$SEL3_17774_out0;
wire  [7:0] v$SEL3_17817_out0;
wire  [7:0] v$SEL3_17818_out0;
wire  [7:0] v$SEL4_11854_out0;
wire  [7:0] v$SEL4_11855_out0;
wire  [7:0] v$SEL4_12199_out0;
wire  [7:0] v$SEL4_12200_out0;
wire  [7:0] v$SHIFT$AMOUNT_7387_out0;
wire  [7:0] v$SHIFT$AMOUNT_7388_out0;
wire  [7:0] v$SHIFT$AMOUNT_7389_out0;
wire  [7:0] v$SHIFT$AMOUNT_7390_out0;
wire  [7:0] v$SHIFT$AMOUNT_7391_out0;
wire  [7:0] v$SHIFT$AMOUNT_7392_out0;
wire  [7:0] v$SHIFT$AMOUNT_7393_out0;
wire  [7:0] v$SHIFT$AMOUNT_7394_out0;
wire  [7:0] v$SINGLE$EXPONENT_7086_out0;
wire  [7:0] v$SINGLE$EXPONENT_7087_out0;
wire  [7:0] v$SINGLE$PRECISION$EXPONENT_11046_out0;
wire  [7:0] v$SINGLE$PRECISION$EXPONENT_11047_out0;
wire  [7:0] v$SMALLER$EXP_2942_out0;
wire  [7:0] v$SMALLER$EXP_2944_out0;
wire  [7:0] v$STATUS_31_out0;
wire  [7:0] v$STATUS_32_out0;
wire  [7:0] v$STATUS_8810_out0;
wire  [7:0] v$STATUS_8811_out0;
wire  [7:0] v$Status_3791_out0;
wire  [7:0] v$Status_3792_out0;
wire  [7:0] v$XOR1_14547_out0;
wire  [7:0] v$XOR1_14548_out0;
wire  [7:0] v$XOR1_7590_out0;
wire  [7:0] v$XOR1_7592_out0;
wire  [7:0] v$XOR1_7594_out0;
wire  [7:0] v$XOR1_7596_out0;
wire  [7:0] v$_10370_out0;
wire  [7:0] v$_10371_out0;
wire  [7:0] v$_1173_out0;
wire  [7:0] v$_1174_out0;
wire  [7:0] v$_1175_out0;
wire  [7:0] v$_1176_out0;
wire  [7:0] v$_1177_out0;
wire  [7:0] v$_12902_out1;
wire  [7:0] v$_12903_out1;
wire  [7:0] v$_13271_out0;
wire  [7:0] v$_13274_out0;
wire  [7:0] v$_14093_out0;
wire  [7:0] v$_14094_out0;
wire  [7:0] v$_14313_out0;
wire  [7:0] v$_14314_out0;
wire  [7:0] v$_14602_out0;
wire  [7:0] v$_14606_out0;
wire  [7:0] v$_14636_out0;
wire  [7:0] v$_14640_out0;
wire  [7:0] v$_14651_out0;
wire  [7:0] v$_14652_out0;
wire  [7:0] v$_1528_out0;
wire  [7:0] v$_1528_out1;
wire  [7:0] v$_1529_out0;
wire  [7:0] v$_1529_out1;
wire  [7:0] v$_15670_out0;
wire  [7:0] v$_15671_out0;
wire  [7:0] v$_16169_out0;
wire  [7:0] v$_16170_out0;
wire  [7:0] v$_1669_out0;
wire  [7:0] v$_1670_out0;
wire  [7:0] v$_1671_out0;
wire  [7:0] v$_1671_out1;
wire  [7:0] v$_1672_out0;
wire  [7:0] v$_1672_out1;
wire  [7:0] v$_16750_out0;
wire  [7:0] v$_16754_out0;
wire  [7:0] v$_16760_out0;
wire  [7:0] v$_16760_out1;
wire  [7:0] v$_16761_out0;
wire  [7:0] v$_16761_out1;
wire  [7:0] v$_17353_out0;
wire  [7:0] v$_17354_out0;
wire  [7:0] v$_17355_out0;
wire  [7:0] v$_17356_out0;
wire  [7:0] v$_17357_out0;
wire  [7:0] v$_17405_out0;
wire  [7:0] v$_17406_out0;
wire  [7:0] v$_17748_out0;
wire  [7:0] v$_17749_out0;
wire  [7:0] v$_17750_out0;
wire  [7:0] v$_17751_out0;
wire  [7:0] v$_17752_out0;
wire  [7:0] v$_3687_out0;
wire  [7:0] v$_3688_out0;
wire  [7:0] v$_4092_out0;
wire  [7:0] v$_4093_out0;
wire  [7:0] v$_4094_out0;
wire  [7:0] v$_4095_out0;
wire  [7:0] v$_4096_out0;
wire  [7:0] v$_4803_out0;
wire  [7:0] v$_4807_out0;
wire  [7:0] v$_6658_out0;
wire  [7:0] v$_6659_out0;
wire  [7:0] v$_6660_out0;
wire  [7:0] v$_6661_out0;
wire  [7:0] v$_6662_out0;
wire  [7:0] v$_7277_out1;
wire  [7:0] v$_7610_out0;
wire  [7:0] v$_7611_out0;
wire  [7:0] v$_7790_out0;
wire  [7:0] v$_7791_out0;
wire  [7:0] v$_7792_out0;
wire  [7:0] v$_7793_out0;
wire  [7:0] v$_7794_out0;
wire  [7:0] v$_7902_out0;
wire  [7:0] v$_7902_out1;
wire  [7:0] v$_7903_out0;
wire  [7:0] v$_7903_out1;
wire  [7:0] v$_8976_out0;
wire  [7:0] v$_8976_out1;
wire  [7:0] v$_8977_out0;
wire  [7:0] v$_8977_out1;
wire  [7:0] v$_9043_out0;
wire  [7:0] v$_9044_out0;
wire  [9:0] v$HALF$PRECISION$MANTISA$DENORM_14497_out0;
wire  [9:0] v$HALF$PRECISION$MANTISA$DENORM_14498_out0;
wire  [9:0] v$SEL10_3207_out0;
wire  [9:0] v$SEL10_3208_out0;
wire  [9:0] v$SEL12_16_out0;
wire  [9:0] v$SEL12_17_out0;
wire  [9:0] v$SEL2_8098_out0;
wire  [9:0] v$SEL2_8099_out0;
wire  [9:0] v$SEL5_7812_out0;
wire  [9:0] v$SEL5_7813_out0;
wire  [9:0] v$SEL7_12476_out0;
wire  [9:0] v$SEL7_12477_out0;
wire  [9:0] v$SEL7_3274_out0;
wire  [9:0] v$SEL7_3275_out0;
wire  [9:0] v$SEL9_9969_out0;
wire  [9:0] v$SEL9_9970_out0;
wire v$1_1533_out0;
wire v$1_1534_out0;
wire v$2StopBits_3484_out0;
wire v$2StopBits_3485_out0;
wire v$32$BIT$INPUT_203_out0;
wire v$32$BIT$VIEWER$IN$FPU_4384_out0;
wire v$32BIT_10932_out0;
wire v$32BIT_10933_out0;
wire v$32BIT_15872_out0;
wire v$32BIT_15873_out0;
wire v$4_15164_out0;
wire v$4_15165_out0;
wire v$5_12290_out0;
wire v$5_12291_out0;
wire v$6_1948_out0;
wire v$6_1949_out0;
wire v$6_9868_out0;
wire v$6_9869_out0;
wire v$7_15358_out0;
wire v$7_15359_out0;
wire v$8_15540_out0;
wire v$8_15541_out0;
wire v$A$EXP$LARGER_17482_out0;
wire v$A$EXP$LARGER_17483_out0;
wire v$A$EXP$LARGER_18245_out0;
wire v$A$EXP$LARGER_18246_out0;
wire v$A$EXP$LARGER_9441_out0;
wire v$A$EXP$LARGER_9442_out0;
wire v$A$IS$OP1_5005_out0;
wire v$A$IS$OP1_5006_out0;
wire v$A$MANTISA$LARGER_14712_out0;
wire v$A$MANTISA$LARGER_14713_out0;
wire v$A$MANTISA$LARGER_16027_out0;
wire v$A$MANTISA$LARGER_16028_out0;
wire v$A0$COMP$B0_7986_out0;
wire v$A0$COMP$B0_7987_out0;
wire v$A0$COMP$B0_7988_out0;
wire v$A0$COMP$B0_7989_out0;
wire v$A0$COMP$B0_7990_out0;
wire v$A0$COMP$B0_7991_out0;
wire v$A0$COMP$B0_7992_out0;
wire v$A0$COMP$B0_7993_out0;
wire v$A0$COMP$B0_7994_out0;
wire v$A0$COMP$B0_7995_out0;
wire v$A0$COMP$B0_7996_out0;
wire v$A0$COMP$B0_7997_out0;
wire v$A0$COMP$B0_7998_out0;
wire v$A0$COMP$B0_7999_out0;
wire v$A0$COMP$B0_8000_out0;
wire v$A0$COMP$B0_8001_out0;
wire v$A0$COMP$B0_8002_out0;
wire v$A0$COMP$B0_8003_out0;
wire v$A0$COMP$B0_8004_out0;
wire v$A0$COMP$B0_8005_out0;
wire v$A0$COMP$B0_8006_out0;
wire v$A0$COMP$B0_8007_out0;
wire v$A0$COMP$B0_8008_out0;
wire v$A0$COMP$B0_8009_out0;
wire v$A0XNORB0_1432_out0;
wire v$A0XNORB0_1433_out0;
wire v$A0XNORB0_1434_out0;
wire v$A0XNORB0_1435_out0;
wire v$A0XNORB0_1436_out0;
wire v$A0XNORB0_1437_out0;
wire v$A0XNORB0_1438_out0;
wire v$A0XNORB0_1439_out0;
wire v$A0XNORB0_1440_out0;
wire v$A0XNORB0_1441_out0;
wire v$A0XNORB0_1442_out0;
wire v$A0XNORB0_1443_out0;
wire v$A0XNORB0_1444_out0;
wire v$A0XNORB0_1445_out0;
wire v$A0XNORB0_1446_out0;
wire v$A0XNORB0_1447_out0;
wire v$A0XNORB0_1448_out0;
wire v$A0XNORB0_1449_out0;
wire v$A0XNORB0_1450_out0;
wire v$A0XNORB0_1451_out0;
wire v$A0XNORB0_1452_out0;
wire v$A0XNORB0_1453_out0;
wire v$A0XNORB0_1454_out0;
wire v$A0XNORB0_1455_out0;
wire v$A0_1725_out0;
wire v$A0_1726_out0;
wire v$A0_1727_out0;
wire v$A0_1728_out0;
wire v$A0_1729_out0;
wire v$A0_1730_out0;
wire v$A0_1731_out0;
wire v$A0_1732_out0;
wire v$A0_1733_out0;
wire v$A0_1734_out0;
wire v$A0_1735_out0;
wire v$A0_1736_out0;
wire v$A0_1737_out0;
wire v$A0_1738_out0;
wire v$A0_1739_out0;
wire v$A0_1740_out0;
wire v$A0_1741_out0;
wire v$A0_1742_out0;
wire v$A0_1743_out0;
wire v$A0_1744_out0;
wire v$A0_1745_out0;
wire v$A0_1746_out0;
wire v$A0_1747_out0;
wire v$A0_1748_out0;
wire v$A0_4308_out0;
wire v$A0_4309_out0;
wire v$A0_4310_out0;
wire v$A0_4311_out0;
wire v$A0_4312_out0;
wire v$A1$COMP$B1_12486_out0;
wire v$A1$COMP$B1_12487_out0;
wire v$A1$COMP$B1_12488_out0;
wire v$A1$COMP$B1_12489_out0;
wire v$A1$COMP$B1_12490_out0;
wire v$A1$COMP$B1_12491_out0;
wire v$A1$COMP$B1_12492_out0;
wire v$A1$COMP$B1_12493_out0;
wire v$A1$COMP$B1_12494_out0;
wire v$A1$COMP$B1_12495_out0;
wire v$A1$COMP$B1_12496_out0;
wire v$A1$COMP$B1_12497_out0;
wire v$A1$COMP$B1_12498_out0;
wire v$A1$COMP$B1_12499_out0;
wire v$A1$COMP$B1_12500_out0;
wire v$A1$COMP$B1_12501_out0;
wire v$A1$COMP$B1_12502_out0;
wire v$A1$COMP$B1_12503_out0;
wire v$A1$COMP$B1_12504_out0;
wire v$A1$COMP$B1_12505_out0;
wire v$A1$COMP$B1_12506_out0;
wire v$A1$COMP$B1_12507_out0;
wire v$A1$COMP$B1_12508_out0;
wire v$A1$COMP$B1_12509_out0;
wire v$A10A_16002_out0;
wire v$A10A_16002_out1;
wire v$A10A_16003_out0;
wire v$A10A_16003_out1;
wire v$A10A_16004_out0;
wire v$A10A_16004_out1;
wire v$A10A_16005_out0;
wire v$A10A_16005_out1;
wire v$A10A_16006_out0;
wire v$A10A_16006_out1;
wire v$A10_1548_out0;
wire v$A10_1549_out0;
wire v$A10_1550_out0;
wire v$A10_1551_out0;
wire v$A10_1552_out0;
wire v$A11_17874_out0;
wire v$A11_17874_out1;
wire v$A11_17875_out0;
wire v$A11_17875_out1;
wire v$A11_17876_out0;
wire v$A11_17876_out1;
wire v$A11_17877_out0;
wire v$A11_17877_out1;
wire v$A11_17878_out0;
wire v$A11_17878_out1;
wire v$A11_9962_out0;
wire v$A11_9963_out0;
wire v$A11_9964_out0;
wire v$A11_9965_out0;
wire v$A11_9966_out0;
wire v$A12A_4445_out0;
wire v$A12A_4445_out1;
wire v$A12A_4446_out0;
wire v$A12A_4446_out1;
wire v$A12A_4447_out0;
wire v$A12A_4447_out1;
wire v$A12A_4448_out0;
wire v$A12A_4448_out1;
wire v$A12A_4449_out0;
wire v$A12A_4449_out1;
wire v$A12_3138_out0;
wire v$A12_3139_out0;
wire v$A12_3140_out0;
wire v$A12_3141_out0;
wire v$A12_3142_out0;
wire v$A13_13862_out0;
wire v$A13_13863_out0;
wire v$A13_13864_out0;
wire v$A13_13865_out0;
wire v$A13_13866_out0;
wire v$A13_7240_out0;
wire v$A13_7240_out1;
wire v$A13_7241_out0;
wire v$A13_7241_out1;
wire v$A13_7242_out0;
wire v$A13_7242_out1;
wire v$A13_7243_out0;
wire v$A13_7243_out1;
wire v$A13_7244_out0;
wire v$A13_7244_out1;
wire v$A14_15353_out0;
wire v$A14_15353_out1;
wire v$A14_15354_out0;
wire v$A14_15354_out1;
wire v$A14_15355_out0;
wire v$A14_15355_out1;
wire v$A14_15356_out0;
wire v$A14_15356_out1;
wire v$A14_15357_out0;
wire v$A14_15357_out1;
wire v$A14_676_out0;
wire v$A14_677_out0;
wire v$A14_678_out0;
wire v$A14_679_out0;
wire v$A14_680_out0;
wire v$A15_13216_out0;
wire v$A15_13216_out1;
wire v$A15_13217_out0;
wire v$A15_13217_out1;
wire v$A15_13218_out0;
wire v$A15_13218_out1;
wire v$A15_13219_out0;
wire v$A15_13219_out1;
wire v$A15_13220_out0;
wire v$A15_13220_out1;
wire v$A15_17318_out0;
wire v$A15_17319_out0;
wire v$A15_17320_out0;
wire v$A15_17321_out0;
wire v$A15_17322_out0;
wire v$A16A_14559_out0;
wire v$A16A_14559_out1;
wire v$A16A_14560_out0;
wire v$A16A_14560_out1;
wire v$A16A_14561_out0;
wire v$A16A_14561_out1;
wire v$A16A_14562_out0;
wire v$A16A_14562_out1;
wire v$A16A_14563_out0;
wire v$A16A_14563_out1;
wire v$A16_13614_out0;
wire v$A16_13615_out0;
wire v$A16_13616_out0;
wire v$A16_13617_out0;
wire v$A16_13618_out0;
wire v$A17A_2487_out0;
wire v$A17A_2487_out1;
wire v$A17A_2488_out0;
wire v$A17A_2488_out1;
wire v$A17A_2489_out0;
wire v$A17A_2489_out1;
wire v$A17A_2490_out0;
wire v$A17A_2490_out1;
wire v$A17A_2491_out0;
wire v$A17A_2491_out1;
wire v$A17_16722_out0;
wire v$A17_16723_out0;
wire v$A17_16724_out0;
wire v$A17_16725_out0;
wire v$A17_16726_out0;
wire v$A18_10032_out0;
wire v$A18_10032_out1;
wire v$A18_10033_out0;
wire v$A18_10033_out1;
wire v$A18_10034_out0;
wire v$A18_10034_out1;
wire v$A18_10035_out0;
wire v$A18_10035_out1;
wire v$A18_10036_out0;
wire v$A18_10036_out1;
wire v$A18_17695_out0;
wire v$A18_17696_out0;
wire v$A18_17697_out0;
wire v$A18_17698_out0;
wire v$A18_17699_out0;
wire v$A19_1213_out0;
wire v$A19_1214_out0;
wire v$A19_1215_out0;
wire v$A19_1216_out0;
wire v$A19_1217_out0;
wire v$A19_15908_out0;
wire v$A19_15908_out1;
wire v$A19_15909_out0;
wire v$A19_15909_out1;
wire v$A19_15910_out0;
wire v$A19_15910_out1;
wire v$A19_15911_out0;
wire v$A19_15911_out1;
wire v$A19_15912_out0;
wire v$A19_15912_out1;
wire v$A1A_11660_out0;
wire v$A1A_11660_out1;
wire v$A1A_11661_out0;
wire v$A1A_11661_out1;
wire v$A1A_11662_out0;
wire v$A1A_11662_out1;
wire v$A1A_11663_out0;
wire v$A1A_11663_out1;
wire v$A1A_11664_out0;
wire v$A1A_11664_out1;
wire v$A1XNORB1_16045_out0;
wire v$A1XNORB1_16046_out0;
wire v$A1XNORB1_16047_out0;
wire v$A1XNORB1_16048_out0;
wire v$A1XNORB1_16049_out0;
wire v$A1XNORB1_16050_out0;
wire v$A1XNORB1_16051_out0;
wire v$A1XNORB1_16052_out0;
wire v$A1XNORB1_16053_out0;
wire v$A1XNORB1_16054_out0;
wire v$A1XNORB1_16055_out0;
wire v$A1XNORB1_16056_out0;
wire v$A1XNORB1_16057_out0;
wire v$A1XNORB1_16058_out0;
wire v$A1XNORB1_16059_out0;
wire v$A1XNORB1_16060_out0;
wire v$A1XNORB1_16061_out0;
wire v$A1XNORB1_16062_out0;
wire v$A1XNORB1_16063_out0;
wire v$A1XNORB1_16064_out0;
wire v$A1XNORB1_16065_out0;
wire v$A1XNORB1_16066_out0;
wire v$A1XNORB1_16067_out0;
wire v$A1XNORB1_16068_out0;
wire v$A1_11802_out1;
wire v$A1_11803_out1;
wire v$A1_13701_out1;
wire v$A1_13702_out1;
wire v$A1_14339_out0;
wire v$A1_14340_out0;
wire v$A1_14341_out0;
wire v$A1_14342_out0;
wire v$A1_14343_out0;
wire v$A1_14344_out0;
wire v$A1_14345_out0;
wire v$A1_14346_out0;
wire v$A1_14347_out0;
wire v$A1_14348_out0;
wire v$A1_14349_out0;
wire v$A1_14350_out0;
wire v$A1_14351_out0;
wire v$A1_14352_out0;
wire v$A1_14353_out0;
wire v$A1_14354_out0;
wire v$A1_14355_out0;
wire v$A1_14356_out0;
wire v$A1_14357_out0;
wire v$A1_14358_out0;
wire v$A1_14359_out0;
wire v$A1_14360_out0;
wire v$A1_14361_out0;
wire v$A1_14362_out0;
wire v$A1_14820_out1;
wire v$A1_14821_out1;
wire v$A1_15214_out1;
wire v$A1_15215_out1;
wire v$A1_15216_out1;
wire v$A1_15217_out1;
wire v$A1_15218_out1;
wire v$A1_15219_out1;
wire v$A1_15220_out1;
wire v$A1_15221_out1;
wire v$A1_15222_out1;
wire v$A1_15223_out1;
wire v$A1_15224_out1;
wire v$A1_15225_out1;
wire v$A1_15763_out1;
wire v$A1_15764_out1;
wire v$A1_1710_out0;
wire v$A1_1711_out0;
wire v$A1_1712_out0;
wire v$A1_1713_out0;
wire v$A1_1714_out0;
wire v$A1_2662_out1;
wire v$A1_2663_out1;
wire v$A1_2664_out1;
wire v$A1_2665_out1;
wire v$A1_2938_out1;
wire v$A1_4011_out1;
wire v$A1_4012_out1;
wire v$A1_5789_out1;
wire v$A1_5790_out1;
wire v$A1_5791_out1;
wire v$A1_5792_out1;
wire v$A1_5793_out1;
wire v$A1_5794_out1;
wire v$A1_5795_out1;
wire v$A1_5796_out1;
wire v$A1_638_out1;
wire v$A1_639_out1;
wire v$A1_6409_out1;
wire v$A1_6410_out1;
wire v$A1_7730_out1;
wire v$A1_7731_out1;
wire v$A1_9430_out1;
wire v$A1_9431_out1;
wire v$A2$COMP$B2_1972_out0;
wire v$A2$COMP$B2_1973_out0;
wire v$A2$COMP$B2_1974_out0;
wire v$A2$COMP$B2_1975_out0;
wire v$A2$COMP$B2_1976_out0;
wire v$A2$COMP$B2_1977_out0;
wire v$A2$COMP$B2_1978_out0;
wire v$A2$COMP$B2_1979_out0;
wire v$A2$COMP$B2_1980_out0;
wire v$A2$COMP$B2_1981_out0;
wire v$A2$COMP$B2_1982_out0;
wire v$A2$COMP$B2_1983_out0;
wire v$A2$COMP$B2_1984_out0;
wire v$A2$COMP$B2_1985_out0;
wire v$A2$COMP$B2_1986_out0;
wire v$A2$COMP$B2_1987_out0;
wire v$A2$COMP$B2_1988_out0;
wire v$A2$COMP$B2_1989_out0;
wire v$A2$COMP$B2_1990_out0;
wire v$A2$COMP$B2_1991_out0;
wire v$A2$COMP$B2_1992_out0;
wire v$A2$COMP$B2_1993_out0;
wire v$A2$COMP$B2_1994_out0;
wire v$A2$COMP$B2_1995_out0;
wire v$A20_16374_out0;
wire v$A20_16374_out1;
wire v$A20_16375_out0;
wire v$A20_16375_out1;
wire v$A20_16376_out0;
wire v$A20_16376_out1;
wire v$A20_16377_out0;
wire v$A20_16377_out1;
wire v$A20_16378_out0;
wire v$A20_16378_out1;
wire v$A20_4436_out0;
wire v$A20_4437_out0;
wire v$A20_4438_out0;
wire v$A20_4439_out0;
wire v$A20_4440_out0;
wire v$A21_18568_out0;
wire v$A21_18568_out1;
wire v$A21_18569_out0;
wire v$A21_18569_out1;
wire v$A21_18570_out0;
wire v$A21_18570_out1;
wire v$A21_18571_out0;
wire v$A21_18571_out1;
wire v$A21_18572_out0;
wire v$A21_18572_out1;
wire v$A21_2598_out0;
wire v$A21_2599_out0;
wire v$A21_2600_out0;
wire v$A21_2601_out0;
wire v$A21_2602_out0;
wire v$A22_17488_out0;
wire v$A22_17488_out1;
wire v$A22_17489_out0;
wire v$A22_17489_out1;
wire v$A22_17490_out0;
wire v$A22_17490_out1;
wire v$A22_17491_out0;
wire v$A22_17491_out1;
wire v$A22_17492_out0;
wire v$A22_17492_out1;
wire v$A22_4424_out0;
wire v$A22_4425_out0;
wire v$A22_4426_out0;
wire v$A22_4427_out0;
wire v$A22_4428_out0;
wire v$A23_5063_out0;
wire v$A23_5064_out0;
wire v$A23_5065_out0;
wire v$A23_5066_out0;
wire v$A23_5067_out0;
wire v$A23_9546_out0;
wire v$A23_9546_out1;
wire v$A23_9547_out0;
wire v$A23_9547_out1;
wire v$A23_9548_out0;
wire v$A23_9548_out1;
wire v$A23_9549_out0;
wire v$A23_9549_out1;
wire v$A23_9550_out0;
wire v$A23_9550_out1;
wire v$A24_16973_out0;
wire v$A24_16973_out1;
wire v$A24_16974_out0;
wire v$A24_16974_out1;
wire v$A24_16975_out0;
wire v$A24_16975_out1;
wire v$A24_16976_out0;
wire v$A24_16976_out1;
wire v$A24_16977_out0;
wire v$A24_16977_out1;
wire v$A2A_1631_out0;
wire v$A2A_1631_out1;
wire v$A2A_1632_out0;
wire v$A2A_1632_out1;
wire v$A2A_1633_out0;
wire v$A2A_1633_out1;
wire v$A2A_1634_out0;
wire v$A2A_1634_out1;
wire v$A2A_1635_out0;
wire v$A2A_1635_out1;
wire v$A2XNORB2_4490_out0;
wire v$A2XNORB2_4491_out0;
wire v$A2XNORB2_4492_out0;
wire v$A2XNORB2_4493_out0;
wire v$A2XNORB2_4494_out0;
wire v$A2XNORB2_4495_out0;
wire v$A2XNORB2_4496_out0;
wire v$A2XNORB2_4497_out0;
wire v$A2XNORB2_4498_out0;
wire v$A2XNORB2_4499_out0;
wire v$A2XNORB2_4500_out0;
wire v$A2XNORB2_4501_out0;
wire v$A2XNORB2_4502_out0;
wire v$A2XNORB2_4503_out0;
wire v$A2XNORB2_4504_out0;
wire v$A2XNORB2_4505_out0;
wire v$A2XNORB2_4506_out0;
wire v$A2XNORB2_4507_out0;
wire v$A2XNORB2_4508_out0;
wire v$A2XNORB2_4509_out0;
wire v$A2XNORB2_4510_out0;
wire v$A2XNORB2_4511_out0;
wire v$A2XNORB2_4512_out0;
wire v$A2XNORB2_4513_out0;
wire v$A2_10044_out1;
wire v$A2_10045_out1;
wire v$A2_10046_out1;
wire v$A2_10047_out1;
wire v$A2_14825_out1;
wire v$A2_14826_out1;
wire v$A2_18266_out0;
wire v$A2_18267_out0;
wire v$A2_18268_out0;
wire v$A2_18269_out0;
wire v$A2_18270_out0;
wire v$A2_8057_out0;
wire v$A2_8058_out0;
wire v$A2_8059_out0;
wire v$A2_8060_out0;
wire v$A2_8061_out0;
wire v$A2_8062_out0;
wire v$A2_8063_out0;
wire v$A2_8064_out0;
wire v$A2_8065_out0;
wire v$A2_8066_out0;
wire v$A2_8067_out0;
wire v$A2_8068_out0;
wire v$A2_8069_out0;
wire v$A2_8070_out0;
wire v$A2_8071_out0;
wire v$A2_8072_out0;
wire v$A2_8073_out0;
wire v$A2_8074_out0;
wire v$A2_8075_out0;
wire v$A2_8076_out0;
wire v$A2_8077_out0;
wire v$A2_8078_out0;
wire v$A2_8079_out0;
wire v$A2_8080_out0;
wire v$A3$COMP$B3_4945_out0;
wire v$A3$COMP$B3_4946_out0;
wire v$A3$COMP$B3_4947_out0;
wire v$A3$COMP$B3_4948_out0;
wire v$A3$COMP$B3_4949_out0;
wire v$A3$COMP$B3_4950_out0;
wire v$A3$COMP$B3_4951_out0;
wire v$A3$COMP$B3_4952_out0;
wire v$A3$COMP$B3_4953_out0;
wire v$A3$COMP$B3_4954_out0;
wire v$A3$COMP$B3_4955_out0;
wire v$A3$COMP$B3_4956_out0;
wire v$A3$COMP$B3_4957_out0;
wire v$A3$COMP$B3_4958_out0;
wire v$A3$COMP$B3_4959_out0;
wire v$A3$COMP$B3_4960_out0;
wire v$A3$COMP$B3_4961_out0;
wire v$A3$COMP$B3_4962_out0;
wire v$A3$COMP$B3_4963_out0;
wire v$A3$COMP$B3_4964_out0;
wire v$A3$COMP$B3_4965_out0;
wire v$A3$COMP$B3_4966_out0;
wire v$A3$COMP$B3_4967_out0;
wire v$A3$COMP$B3_4968_out0;
wire v$A3A_11951_out0;
wire v$A3A_11951_out1;
wire v$A3A_11952_out0;
wire v$A3A_11952_out1;
wire v$A3A_11953_out0;
wire v$A3A_11953_out1;
wire v$A3A_11954_out0;
wire v$A3A_11954_out1;
wire v$A3A_11955_out0;
wire v$A3A_11955_out1;
wire v$A3XNORB3_14716_out0;
wire v$A3XNORB3_14717_out0;
wire v$A3XNORB3_14718_out0;
wire v$A3XNORB3_14719_out0;
wire v$A3XNORB3_14720_out0;
wire v$A3XNORB3_14721_out0;
wire v$A3XNORB3_14722_out0;
wire v$A3XNORB3_14723_out0;
wire v$A3XNORB3_14724_out0;
wire v$A3XNORB3_14725_out0;
wire v$A3XNORB3_14726_out0;
wire v$A3XNORB3_14727_out0;
wire v$A3XNORB3_14728_out0;
wire v$A3XNORB3_14729_out0;
wire v$A3XNORB3_14730_out0;
wire v$A3XNORB3_14731_out0;
wire v$A3XNORB3_14732_out0;
wire v$A3XNORB3_14733_out0;
wire v$A3XNORB3_14734_out0;
wire v$A3XNORB3_14735_out0;
wire v$A3XNORB3_14736_out0;
wire v$A3XNORB3_14737_out0;
wire v$A3XNORB3_14738_out0;
wire v$A3XNORB3_14739_out0;
wire v$A3_10702_out0;
wire v$A3_10703_out0;
wire v$A3_10704_out0;
wire v$A3_10705_out0;
wire v$A3_10706_out0;
wire v$A3_10707_out0;
wire v$A3_10708_out0;
wire v$A3_10709_out0;
wire v$A3_10710_out0;
wire v$A3_10711_out0;
wire v$A3_10712_out0;
wire v$A3_10713_out0;
wire v$A3_10714_out0;
wire v$A3_10715_out0;
wire v$A3_10716_out0;
wire v$A3_10717_out0;
wire v$A3_10718_out0;
wire v$A3_10719_out0;
wire v$A3_10720_out0;
wire v$A3_10721_out0;
wire v$A3_10722_out0;
wire v$A3_10723_out0;
wire v$A3_10724_out0;
wire v$A3_10725_out0;
wire v$A3_14607_out0;
wire v$A3_14608_out0;
wire v$A3_14609_out0;
wire v$A3_14610_out0;
wire v$A3_14611_out0;
wire v$A4$COMP$B4_7409_out0;
wire v$A4$COMP$B4_7410_out0;
wire v$A4$COMP$B4_7411_out0;
wire v$A4$COMP$B4_7412_out0;
wire v$A4A_13154_out0;
wire v$A4A_13154_out1;
wire v$A4A_13155_out0;
wire v$A4A_13155_out1;
wire v$A4A_13156_out0;
wire v$A4A_13156_out1;
wire v$A4A_13157_out0;
wire v$A4A_13157_out1;
wire v$A4A_13158_out0;
wire v$A4A_13158_out1;
wire v$A4XNORB4_1372_out0;
wire v$A4XNORB4_1373_out0;
wire v$A4XNORB4_1374_out0;
wire v$A4XNORB4_1375_out0;
wire v$A4_15007_out0;
wire v$A4_15008_out0;
wire v$A4_15009_out0;
wire v$A4_15010_out0;
wire v$A4_17498_out0;
wire v$A4_17499_out0;
wire v$A4_17500_out0;
wire v$A4_17501_out0;
wire v$A4_17502_out0;
wire v$A5A_16099_out0;
wire v$A5A_16099_out1;
wire v$A5A_16100_out0;
wire v$A5A_16100_out1;
wire v$A5A_16101_out0;
wire v$A5A_16101_out1;
wire v$A5A_16102_out0;
wire v$A5A_16102_out1;
wire v$A5A_16103_out0;
wire v$A5A_16103_out1;
wire v$A5_6665_out0;
wire v$A5_6666_out0;
wire v$A5_6667_out0;
wire v$A5_6668_out0;
wire v$A5_6669_out0;
wire v$A6A_3121_out0;
wire v$A6A_3121_out1;
wire v$A6A_3122_out0;
wire v$A6A_3122_out1;
wire v$A6A_3123_out0;
wire v$A6A_3123_out1;
wire v$A6A_3124_out0;
wire v$A6A_3124_out1;
wire v$A6A_3125_out0;
wire v$A6A_3125_out1;
wire v$A6_308_out0;
wire v$A6_309_out0;
wire v$A6_310_out0;
wire v$A6_311_out0;
wire v$A6_312_out0;
wire v$A7A_1657_out0;
wire v$A7A_1657_out1;
wire v$A7A_1658_out0;
wire v$A7A_1658_out1;
wire v$A7A_1659_out0;
wire v$A7A_1659_out1;
wire v$A7A_1660_out0;
wire v$A7A_1660_out1;
wire v$A7A_1661_out0;
wire v$A7A_1661_out1;
wire v$A7_15307_out0;
wire v$A7_15308_out0;
wire v$A7_15309_out0;
wire v$A7_15310_out0;
wire v$A7_15311_out0;
wire v$A8A_1505_out0;
wire v$A8A_1505_out1;
wire v$A8A_1506_out0;
wire v$A8A_1506_out1;
wire v$A8A_1507_out0;
wire v$A8A_1507_out1;
wire v$A8A_1508_out0;
wire v$A8A_1508_out1;
wire v$A8A_1509_out0;
wire v$A8A_1509_out1;
wire v$A8_18090_out0;
wire v$A8_18091_out0;
wire v$A8_18092_out0;
wire v$A8_18093_out0;
wire v$A8_18094_out0;
wire v$A9A_10411_out0;
wire v$A9A_10411_out1;
wire v$A9A_10412_out0;
wire v$A9A_10412_out1;
wire v$A9A_10413_out0;
wire v$A9A_10413_out1;
wire v$A9A_10414_out0;
wire v$A9A_10414_out1;
wire v$A9A_10415_out0;
wire v$A9A_10415_out1;
wire v$A9_3435_out0;
wire v$A9_3436_out0;
wire v$A9_3437_out0;
wire v$A9_3438_out0;
wire v$A9_3439_out0;
wire v$AD3$EQUALS$AD2_14557_out0;
wire v$AD3$EQUALS$AD2_14558_out0;
wire v$ADD_8219_out0;
wire v$ADD_8220_out0;
wire v$ARBHALT0_2908_out0;
wire v$ARBHALT1_5453_out0;
wire v$ARR0_10978_out0;
wire v$ARR1_9067_out0;
wire v$AUTODISABLE_18213_out0;
wire v$AUTODISABLE_18214_out0;
wire v$AWR0_1798_out0;
wire v$AWR1_15889_out0;
wire v$A_7101_out0;
wire v$A_7102_out0;
wire v$A_7103_out0;
wire v$A_7104_out0;
wire v$A_7105_out0;
wire v$A_7106_out0;
wire v$A_7107_out0;
wire v$A_7108_out0;
wire v$A_7109_out0;
wire v$A_7110_out0;
wire v$A_7111_out0;
wire v$A_7112_out0;
wire v$A_7113_out0;
wire v$A_7114_out0;
wire v$A_7115_out0;
wire v$A_7116_out0;
wire v$A_7117_out0;
wire v$A_7118_out0;
wire v$A_7119_out0;
wire v$A_7120_out0;
wire v$A_7121_out0;
wire v$A_7122_out0;
wire v$A_7123_out0;
wire v$A_7124_out0;
wire v$A_7125_out0;
wire v$A_7126_out0;
wire v$A_7127_out0;
wire v$A_7128_out0;
wire v$A_7129_out0;
wire v$A_7130_out0;
wire v$A_7131_out0;
wire v$A_7132_out0;
wire v$A_7133_out0;
wire v$A_7134_out0;
wire v$A_7135_out0;
wire v$A_7136_out0;
wire v$A_7137_out0;
wire v$A_7138_out0;
wire v$A_7139_out0;
wire v$A_7140_out0;
wire v$A_7141_out0;
wire v$A_7142_out0;
wire v$A_7143_out0;
wire v$A_7144_out0;
wire v$A_7145_out0;
wire v$A_7146_out0;
wire v$A_7147_out0;
wire v$A_7148_out0;
wire v$A_7149_out0;
wire v$A_7150_out0;
wire v$A_7151_out0;
wire v$A_7152_out0;
wire v$A_7153_out0;
wire v$A_7154_out0;
wire v$A_7155_out0;
wire v$A_7156_out0;
wire v$A_7157_out0;
wire v$A_7158_out0;
wire v$A_7159_out0;
wire v$A_7160_out0;
wire v$A_7161_out0;
wire v$A_7162_out0;
wire v$A_7163_out0;
wire v$A_7164_out0;
wire v$A_7165_out0;
wire v$A_7166_out0;
wire v$A_7167_out0;
wire v$A_7168_out0;
wire v$A_7169_out0;
wire v$A_7170_out0;
wire v$A_7171_out0;
wire v$A_7172_out0;
wire v$A_7173_out0;
wire v$A_7174_out0;
wire v$A_7175_out0;
wire v$A_7176_out0;
wire v$A_7177_out0;
wire v$A_7178_out0;
wire v$A_7179_out0;
wire v$A_7180_out0;
wire v$A_7181_out0;
wire v$A_7182_out0;
wire v$A_7183_out0;
wire v$A_7184_out0;
wire v$A_7185_out0;
wire v$A_7186_out0;
wire v$A_7187_out0;
wire v$A_7188_out0;
wire v$A_7189_out0;
wire v$A_7190_out0;
wire v$A_7191_out0;
wire v$A_7192_out0;
wire v$A_7193_out0;
wire v$A_7194_out0;
wire v$A_7195_out0;
wire v$A_7196_out0;
wire v$A_7197_out0;
wire v$A_7198_out0;
wire v$A_7199_out0;
wire v$A_7200_out0;
wire v$A_7201_out0;
wire v$A_7202_out0;
wire v$A_7203_out0;
wire v$A_7204_out0;
wire v$A_7205_out0;
wire v$A_7206_out0;
wire v$A_7207_out0;
wire v$A_7208_out0;
wire v$A_7209_out0;
wire v$A_7210_out0;
wire v$A_7211_out0;
wire v$A_7212_out0;
wire v$A_7213_out0;
wire v$A_7214_out0;
wire v$A_7215_out0;
wire v$A_7216_out0;
wire v$A_7217_out0;
wire v$A_7218_out0;
wire v$A_7219_out0;
wire v$A_7220_out0;
wire v$B$IS$RD_14084_out0;
wire v$B$IS$RD_14085_out0;
wire v$B0_3200_out0;
wire v$B0_3201_out0;
wire v$B0_3202_out0;
wire v$B0_3203_out0;
wire v$B0_3204_out0;
wire v$B0_3645_out0;
wire v$B0_3646_out0;
wire v$B0_3647_out0;
wire v$B0_3648_out0;
wire v$B0_3649_out0;
wire v$B0_3650_out0;
wire v$B0_3651_out0;
wire v$B0_3652_out0;
wire v$B0_3653_out0;
wire v$B0_3654_out0;
wire v$B0_3655_out0;
wire v$B0_3656_out0;
wire v$B0_3657_out0;
wire v$B0_3658_out0;
wire v$B0_3659_out0;
wire v$B0_3660_out0;
wire v$B0_3661_out0;
wire v$B0_3662_out0;
wire v$B0_3663_out0;
wire v$B0_3664_out0;
wire v$B0_3665_out0;
wire v$B0_3666_out0;
wire v$B0_3667_out0;
wire v$B0_3668_out0;
wire v$B10_9877_out0;
wire v$B10_9878_out0;
wire v$B10_9879_out0;
wire v$B10_9880_out0;
wire v$B10_9881_out0;
wire v$B11_9116_out0;
wire v$B11_9117_out0;
wire v$B11_9118_out0;
wire v$B11_9119_out0;
wire v$B11_9120_out0;
wire v$B12_1950_out0;
wire v$B12_1951_out0;
wire v$B12_1952_out0;
wire v$B12_1953_out0;
wire v$B12_1954_out0;
wire v$B13_8675_out0;
wire v$B13_8676_out0;
wire v$B13_8677_out0;
wire v$B13_8678_out0;
wire v$B13_8679_out0;
wire v$B14_4002_out0;
wire v$B14_4003_out0;
wire v$B14_4004_out0;
wire v$B14_4005_out0;
wire v$B14_4006_out0;
wire v$B15_10021_out0;
wire v$B15_10022_out0;
wire v$B15_10023_out0;
wire v$B15_10024_out0;
wire v$B15_10025_out0;
wire v$B16_16414_out0;
wire v$B16_16415_out0;
wire v$B16_16416_out0;
wire v$B16_16417_out0;
wire v$B16_16418_out0;
wire v$B17_15535_out0;
wire v$B17_15536_out0;
wire v$B17_15537_out0;
wire v$B17_15538_out0;
wire v$B17_15539_out0;
wire v$B18_10867_out0;
wire v$B18_10868_out0;
wire v$B18_10869_out0;
wire v$B18_10870_out0;
wire v$B18_10871_out0;
wire v$B19_16789_out0;
wire v$B19_16790_out0;
wire v$B19_16791_out0;
wire v$B19_16792_out0;
wire v$B19_16793_out0;
wire v$B1_14220_out0;
wire v$B1_14221_out0;
wire v$B1_14222_out0;
wire v$B1_14223_out0;
wire v$B1_14224_out0;
wire v$B1_14225_out0;
wire v$B1_14226_out0;
wire v$B1_14227_out0;
wire v$B1_14228_out0;
wire v$B1_14229_out0;
wire v$B1_14230_out0;
wire v$B1_14231_out0;
wire v$B1_14232_out0;
wire v$B1_14233_out0;
wire v$B1_14234_out0;
wire v$B1_14235_out0;
wire v$B1_14236_out0;
wire v$B1_14237_out0;
wire v$B1_14238_out0;
wire v$B1_14239_out0;
wire v$B1_14240_out0;
wire v$B1_14241_out0;
wire v$B1_14242_out0;
wire v$B1_14243_out0;
wire v$B1_8123_out0;
wire v$B1_8124_out0;
wire v$B1_8125_out0;
wire v$B1_8126_out0;
wire v$B1_8127_out0;
wire v$B20_3943_out0;
wire v$B20_3944_out0;
wire v$B20_3945_out0;
wire v$B20_3946_out0;
wire v$B20_3947_out0;
wire v$B21_18082_out0;
wire v$B21_18083_out0;
wire v$B21_18084_out0;
wire v$B21_18085_out0;
wire v$B21_18086_out0;
wire v$B22_10805_out0;
wire v$B22_10806_out0;
wire v$B22_10807_out0;
wire v$B22_10808_out0;
wire v$B22_10809_out0;
wire v$B23_1283_out0;
wire v$B23_1284_out0;
wire v$B23_1285_out0;
wire v$B23_1286_out0;
wire v$B23_1287_out0;
wire v$B2_16624_out0;
wire v$B2_16625_out0;
wire v$B2_16626_out0;
wire v$B2_16627_out0;
wire v$B2_16628_out0;
wire v$B2_16629_out0;
wire v$B2_16630_out0;
wire v$B2_16631_out0;
wire v$B2_16632_out0;
wire v$B2_16633_out0;
wire v$B2_16634_out0;
wire v$B2_16635_out0;
wire v$B2_16636_out0;
wire v$B2_16637_out0;
wire v$B2_16638_out0;
wire v$B2_16639_out0;
wire v$B2_16640_out0;
wire v$B2_16641_out0;
wire v$B2_16642_out0;
wire v$B2_16643_out0;
wire v$B2_16644_out0;
wire v$B2_16645_out0;
wire v$B2_16646_out0;
wire v$B2_16647_out0;
wire v$B2_3113_out0;
wire v$B2_3114_out0;
wire v$B2_3115_out0;
wire v$B2_3116_out0;
wire v$B2_3117_out0;
wire v$B3_17850_out0;
wire v$B3_17851_out0;
wire v$B3_17852_out0;
wire v$B3_17853_out0;
wire v$B3_17854_out0;
wire v$B3_17855_out0;
wire v$B3_17856_out0;
wire v$B3_17857_out0;
wire v$B3_17858_out0;
wire v$B3_17859_out0;
wire v$B3_17860_out0;
wire v$B3_17861_out0;
wire v$B3_17862_out0;
wire v$B3_17863_out0;
wire v$B3_17864_out0;
wire v$B3_17865_out0;
wire v$B3_17866_out0;
wire v$B3_17867_out0;
wire v$B3_17868_out0;
wire v$B3_17869_out0;
wire v$B3_17870_out0;
wire v$B3_17871_out0;
wire v$B3_17872_out0;
wire v$B3_17873_out0;
wire v$B3_9471_out0;
wire v$B3_9472_out0;
wire v$B3_9473_out0;
wire v$B3_9474_out0;
wire v$B3_9475_out0;
wire v$B4_14663_out0;
wire v$B4_14664_out0;
wire v$B4_14665_out0;
wire v$B4_14666_out0;
wire v$B4_14667_out0;
wire v$B4_16926_out0;
wire v$B4_16927_out0;
wire v$B4_16928_out0;
wire v$B4_16929_out0;
wire v$B5_18374_out0;
wire v$B5_18375_out0;
wire v$B5_18376_out0;
wire v$B5_18377_out0;
wire v$B5_18378_out0;
wire v$B6_13298_out0;
wire v$B6_13299_out0;
wire v$B6_13300_out0;
wire v$B6_13301_out0;
wire v$B6_13302_out0;
wire v$B7_17040_out0;
wire v$B7_17041_out0;
wire v$B7_17042_out0;
wire v$B7_17043_out0;
wire v$B7_17044_out0;
wire v$B8_13138_out0;
wire v$B8_13139_out0;
wire v$B8_13140_out0;
wire v$B8_13141_out0;
wire v$B8_13142_out0;
wire v$B9_4065_out0;
wire v$B9_4066_out0;
wire v$B9_4067_out0;
wire v$B9_4068_out0;
wire v$B9_4069_out0;
wire v$B_2696_out0;
wire v$B_2697_out0;
wire v$B_2698_out0;
wire v$B_2699_out0;
wire v$B_2700_out0;
wire v$B_2701_out0;
wire v$B_2702_out0;
wire v$B_2703_out0;
wire v$B_2704_out0;
wire v$B_2705_out0;
wire v$B_2706_out0;
wire v$B_2707_out0;
wire v$B_2708_out0;
wire v$B_2709_out0;
wire v$B_2710_out0;
wire v$B_2711_out0;
wire v$B_2712_out0;
wire v$B_2713_out0;
wire v$B_2714_out0;
wire v$B_2715_out0;
wire v$B_2716_out0;
wire v$B_2717_out0;
wire v$B_2718_out0;
wire v$B_2719_out0;
wire v$B_2720_out0;
wire v$B_2721_out0;
wire v$B_2722_out0;
wire v$B_2723_out0;
wire v$B_2724_out0;
wire v$B_2725_out0;
wire v$B_2726_out0;
wire v$B_2727_out0;
wire v$B_2728_out0;
wire v$B_2729_out0;
wire v$B_2730_out0;
wire v$B_2731_out0;
wire v$B_2732_out0;
wire v$B_2733_out0;
wire v$B_2734_out0;
wire v$B_2735_out0;
wire v$B_2736_out0;
wire v$B_2737_out0;
wire v$B_2738_out0;
wire v$B_2739_out0;
wire v$B_2740_out0;
wire v$B_2741_out0;
wire v$B_2742_out0;
wire v$B_2743_out0;
wire v$B_2744_out0;
wire v$B_2745_out0;
wire v$B_2746_out0;
wire v$B_2747_out0;
wire v$B_2748_out0;
wire v$B_2749_out0;
wire v$B_2750_out0;
wire v$B_2751_out0;
wire v$B_2752_out0;
wire v$B_2753_out0;
wire v$B_2754_out0;
wire v$B_2755_out0;
wire v$B_2756_out0;
wire v$B_2757_out0;
wire v$B_2758_out0;
wire v$B_2759_out0;
wire v$B_2760_out0;
wire v$B_2761_out0;
wire v$B_2762_out0;
wire v$B_2763_out0;
wire v$B_2764_out0;
wire v$B_2765_out0;
wire v$B_2766_out0;
wire v$B_2767_out0;
wire v$B_2768_out0;
wire v$B_2769_out0;
wire v$B_2770_out0;
wire v$B_2771_out0;
wire v$B_2772_out0;
wire v$B_2773_out0;
wire v$B_2774_out0;
wire v$B_2775_out0;
wire v$B_2776_out0;
wire v$B_2777_out0;
wire v$B_2778_out0;
wire v$B_2779_out0;
wire v$B_2780_out0;
wire v$B_2781_out0;
wire v$B_2782_out0;
wire v$B_2783_out0;
wire v$B_2784_out0;
wire v$B_2785_out0;
wire v$B_2786_out0;
wire v$B_2787_out0;
wire v$B_2788_out0;
wire v$B_2789_out0;
wire v$B_2790_out0;
wire v$B_2791_out0;
wire v$B_2792_out0;
wire v$B_2793_out0;
wire v$B_2794_out0;
wire v$B_2795_out0;
wire v$B_2796_out0;
wire v$B_2797_out0;
wire v$B_2798_out0;
wire v$B_2799_out0;
wire v$B_2800_out0;
wire v$B_2801_out0;
wire v$B_2802_out0;
wire v$B_2803_out0;
wire v$B_2804_out0;
wire v$B_2805_out0;
wire v$B_2806_out0;
wire v$B_2807_out0;
wire v$B_2808_out0;
wire v$B_2809_out0;
wire v$B_2810_out0;
wire v$B_2811_out0;
wire v$B_2812_out0;
wire v$B_2813_out0;
wire v$B_2814_out0;
wire v$B_2815_out0;
wire v$C0_10692_out0;
wire v$C0_10693_out0;
wire v$C0_10694_out0;
wire v$C0_10695_out0;
wire v$C0_10696_out0;
wire v$C0_9374_out0;
wire v$C0_9375_out0;
wire v$C0_9376_out0;
wire v$C0_9377_out0;
wire v$C0_9378_out0;
wire v$C10_12732_out0;
wire v$C10_12733_out0;
wire v$C10_12734_out0;
wire v$C10_12735_out0;
wire v$C10_12736_out0;
wire v$C10_1940_out0;
wire v$C10_1941_out0;
wire v$C10_1942_out0;
wire v$C10_1943_out0;
wire v$C10_1944_out0;
wire v$C11_14796_out0;
wire v$C11_14797_out0;
wire v$C11_14798_out0;
wire v$C11_14799_out0;
wire v$C11_14800_out0;
wire v$C11_3632_out0;
wire v$C11_3633_out0;
wire v$C11_9510_out0;
wire v$C11_9511_out0;
wire v$C11_9512_out0;
wire v$C11_9513_out0;
wire v$C11_9514_out0;
wire v$C12_13520_out0;
wire v$C12_13521_out0;
wire v$C12_13522_out0;
wire v$C12_13523_out0;
wire v$C12_13524_out0;
wire v$C12_9394_out0;
wire v$C12_9395_out0;
wire v$C12_9396_out0;
wire v$C12_9397_out0;
wire v$C12_9398_out0;
wire v$C13_11776_out0;
wire v$C13_11777_out0;
wire v$C13_11778_out0;
wire v$C13_11779_out0;
wire v$C13_11780_out0;
wire v$C13_18589_out0;
wire v$C13_18590_out0;
wire v$C13_18591_out0;
wire v$C13_18592_out0;
wire v$C13_18593_out0;
wire v$C14_279_out0;
wire v$C14_280_out0;
wire v$C14_281_out0;
wire v$C14_282_out0;
wire v$C14_283_out0;
wire v$C14_325_out0;
wire v$C14_326_out0;
wire v$C14_327_out0;
wire v$C14_328_out0;
wire v$C14_329_out0;
wire v$C15_13131_out0;
wire v$C15_13132_out0;
wire v$C15_13133_out0;
wire v$C15_13134_out0;
wire v$C15_13135_out0;
wire v$C15_8143_out0;
wire v$C15_8144_out0;
wire v$C15_8145_out0;
wire v$C15_8146_out0;
wire v$C15_8147_out0;
wire v$C16_1268_out0;
wire v$C16_1269_out0;
wire v$C16_1270_out0;
wire v$C16_1271_out0;
wire v$C16_1272_out0;
wire v$C16_15157_out0;
wire v$C16_15158_out0;
wire v$C16_15159_out0;
wire v$C16_15160_out0;
wire v$C16_15161_out0;
wire v$C17_2520_out0;
wire v$C17_2521_out0;
wire v$C17_2522_out0;
wire v$C17_2523_out0;
wire v$C17_2524_out0;
wire v$C17_6066_out0;
wire v$C17_6067_out0;
wire v$C17_6068_out0;
wire v$C17_6069_out0;
wire v$C17_6070_out0;
wire v$C18_16289_out0;
wire v$C18_16290_out0;
wire v$C18_16291_out0;
wire v$C18_16292_out0;
wire v$C18_16293_out0;
wire v$C18_18005_out0;
wire v$C18_18006_out0;
wire v$C18_18007_out0;
wire v$C18_18008_out0;
wire v$C18_18009_out0;
wire v$C19_13833_out0;
wire v$C19_13834_out0;
wire v$C19_13835_out0;
wire v$C19_13836_out0;
wire v$C19_13837_out0;
wire v$C19_8160_out0;
wire v$C19_8161_out0;
wire v$C19_8162_out0;
wire v$C19_8163_out0;
wire v$C19_8164_out0;
wire v$C1_11849_out0;
wire v$C1_11850_out0;
wire v$C1_11851_out0;
wire v$C1_11852_out0;
wire v$C1_11853_out0;
wire v$C1_12852_out0;
wire v$C1_12853_out0;
wire v$C1_14029_out0;
wire v$C1_1471_out0;
wire v$C1_1472_out0;
wire v$C1_1514_out0;
wire v$C1_1515_out0;
wire v$C1_15720_out0;
wire v$C1_15721_out0;
wire v$C1_15722_out0;
wire v$C1_15723_out0;
wire v$C1_15921_out0;
wire v$C1_15922_out0;
wire v$C1_16781_out0;
wire v$C1_16782_out0;
wire v$C1_16783_out0;
wire v$C1_16784_out0;
wire v$C1_16785_out0;
wire v$C1_17338_out0;
wire v$C1_17339_out0;
wire v$C1_17340_out0;
wire v$C1_17341_out0;
wire v$C1_17666_out0;
wire v$C1_17667_out0;
wire v$C1_17668_out0;
wire v$C1_17669_out0;
wire v$C1_17670_out0;
wire v$C1_17671_out0;
wire v$C1_17672_out0;
wire v$C1_17673_out0;
wire v$C1_2633_out0;
wire v$C1_2634_out0;
wire v$C1_2635_out0;
wire v$C1_2636_out0;
wire v$C1_2637_out0;
wire v$C1_2638_out0;
wire v$C1_2639_out0;
wire v$C1_2640_out0;
wire v$C1_2641_out0;
wire v$C1_2642_out0;
wire v$C1_2643_out0;
wire v$C1_2644_out0;
wire v$C1_4356_out0;
wire v$C1_4357_out0;
wire v$C1_4464_out0;
wire v$C1_4465_out0;
wire v$C1_4466_out0;
wire v$C1_4467_out0;
wire v$C1_4468_out0;
wire v$C1_5434_out0;
wire v$C1_5435_out0;
wire v$C1_5963_out0;
wire v$C1_5968_out0;
wire v$C1_5973_out0;
wire v$C1_5976_out0;
wire v$C1_5983_out0;
wire v$C1_5986_out0;
wire v$C1_5991_out0;
wire v$C1_5994_out0;
wire v$C1_6001_out0;
wire v$C1_6007_out0;
wire v$C1_6011_out0;
wire v$C1_6016_out0;
wire v$C1_6021_out0;
wire v$C1_6457_out0;
wire v$C1_6458_out0;
wire v$C1_7971_out0;
wire v$C1_7975_out0;
wire v$C20_14978_out0;
wire v$C20_14979_out0;
wire v$C20_14980_out0;
wire v$C20_14981_out0;
wire v$C20_14982_out0;
wire v$C20_15489_out0;
wire v$C20_15490_out0;
wire v$C20_15491_out0;
wire v$C20_15492_out0;
wire v$C20_15493_out0;
wire v$C21_10767_out0;
wire v$C21_10768_out0;
wire v$C21_10769_out0;
wire v$C21_10770_out0;
wire v$C21_10771_out0;
wire v$C21_6369_out0;
wire v$C21_6370_out0;
wire v$C21_6371_out0;
wire v$C21_6372_out0;
wire v$C21_6373_out0;
wire v$C22_10981_out0;
wire v$C22_10982_out0;
wire v$C22_10983_out0;
wire v$C22_10984_out0;
wire v$C22_10985_out0;
wire v$C22_8410_out0;
wire v$C22_8411_out0;
wire v$C22_8412_out0;
wire v$C22_8413_out0;
wire v$C22_8414_out0;
wire v$C23_16149_out0;
wire v$C23_16150_out0;
wire v$C23_16151_out0;
wire v$C23_16152_out0;
wire v$C23_16153_out0;
wire v$C23_4843_out0;
wire v$C23_4844_out0;
wire v$C23_4845_out0;
wire v$C23_4846_out0;
wire v$C23_4847_out0;
wire v$C2_105_out0;
wire v$C2_10701_out0;
wire v$C2_110_out0;
wire v$C2_115_out0;
wire v$C2_1171_out0;
wire v$C2_1172_out0;
wire v$C2_118_out0;
wire v$C2_125_out0;
wire v$C2_128_out0;
wire v$C2_133_out0;
wire v$C2_13509_out0;
wire v$C2_13510_out0;
wire v$C2_136_out0;
wire v$C2_143_out0;
wire v$C2_1456_out0;
wire v$C2_1457_out0;
wire v$C2_149_out0;
wire v$C2_15178_out0;
wire v$C2_15179_out0;
wire v$C2_15180_out0;
wire v$C2_15181_out0;
wire v$C2_153_out0;
wire v$C2_158_out0;
wire v$C2_16240_out0;
wire v$C2_16241_out0;
wire v$C2_16281_out0;
wire v$C2_16282_out0;
wire v$C2_16283_out0;
wire v$C2_16284_out0;
wire v$C2_16329_out0;
wire v$C2_16330_out0;
wire v$C2_16331_out0;
wire v$C2_16332_out0;
wire v$C2_163_out0;
wire v$C2_17020_out0;
wire v$C2_17021_out0;
wire v$C2_18179_out0;
wire v$C2_18180_out0;
wire v$C2_18181_out0;
wire v$C2_18182_out0;
wire v$C2_18183_out0;
wire v$C2_18320_out0;
wire v$C2_18321_out0;
wire v$C2_2666_out0;
wire v$C2_2667_out0;
wire v$C2_2686_out0;
wire v$C2_2687_out0;
wire v$C2_2688_out0;
wire v$C2_2689_out0;
wire v$C2_2690_out0;
wire v$C2_2975_out0;
wire v$C2_2976_out0;
wire v$C2_3628_out0;
wire v$C2_3629_out0;
wire v$C2_7624_out0;
wire v$C2_7625_out0;
wire v$C2_7626_out0;
wire v$C2_7627_out0;
wire v$C2_7628_out0;
wire v$C2_7629_out0;
wire v$C2_7630_out0;
wire v$C2_7631_out0;
wire v$C3_13516_out0;
wire v$C3_13517_out0;
wire v$C3_13518_out0;
wire v$C3_13519_out0;
wire v$C3_1362_out0;
wire v$C3_1363_out0;
wire v$C3_15726_out0;
wire v$C3_15727_out0;
wire v$C3_15728_out0;
wire v$C3_15729_out0;
wire v$C3_15730_out0;
wire v$C3_15817_out0;
wire v$C3_15818_out0;
wire v$C3_15819_out0;
wire v$C3_15820_out0;
wire v$C3_15821_out0;
wire v$C3_18128_out0;
wire v$C3_18129_out0;
wire v$C3_18130_out0;
wire v$C3_18552_out0;
wire v$C3_18553_out0;
wire v$C3_5386_out0;
wire v$C3_5387_out0;
wire v$C4_1259_out0;
wire v$C4_1260_out0;
wire v$C4_1261_out0;
wire v$C4_1262_out0;
wire v$C4_1263_out0;
wire v$C4_14830_out0;
wire v$C4_14831_out0;
wire v$C4_14832_out0;
wire v$C4_14833_out0;
wire v$C4_1876_out0;
wire v$C4_1877_out0;
wire v$C4_1878_out0;
wire v$C4_1879_out0;
wire v$C4_1880_out0;
wire v$C4_2920_out0;
wire v$C4_2921_out0;
wire v$C4_3754_out0;
wire v$C4_3755_out0;
wire v$C4_6367_out0;
wire v$C4_6368_out0;
wire v$C5_11686_out0;
wire v$C5_11687_out0;
wire v$C5_11688_out0;
wire v$C5_11689_out0;
wire v$C5_11690_out0;
wire v$C5_15915_out0;
wire v$C5_15916_out0;
wire v$C5_15917_out0;
wire v$C5_15918_out0;
wire v$C5_15919_out0;
wire v$C5_16095_out0;
wire v$C5_16908_out0;
wire v$C5_16910_out0;
wire v$C5_8762_out0;
wire v$C5_8763_out0;
wire v$C5_8764_out0;
wire v$C5_8765_out0;
wire v$C6_11350_out0;
wire v$C6_11351_out0;
wire v$C6_11352_out0;
wire v$C6_11353_out0;
wire v$C6_11354_out0;
wire v$C6_11355_out0;
wire v$C6_11356_out0;
wire v$C6_11357_out0;
wire v$C6_11358_out0;
wire v$C6_11359_out0;
wire v$C6_11360_out0;
wire v$C6_11361_out0;
wire v$C6_12551_out0;
wire v$C6_12552_out0;
wire v$C6_1568_out0;
wire v$C6_1569_out0;
wire v$C6_2432_out0;
wire v$C6_2433_out0;
wire v$C6_7055_out0;
wire v$C6_7056_out0;
wire v$C6_7057_out0;
wire v$C6_7058_out0;
wire v$C6_7059_out0;
wire v$C6_8836_out0;
wire v$C6_9586_out0;
wire v$C6_9587_out0;
wire v$C6_9588_out0;
wire v$C6_9589_out0;
wire v$C6_9590_out0;
wire v$C7_10969_out0;
wire v$C7_10970_out0;
wire v$C7_10971_out0;
wire v$C7_10972_out0;
wire v$C7_10973_out0;
wire v$C7_16430_out0;
wire v$C7_16431_out0;
wire v$C7_16432_out0;
wire v$C7_16433_out0;
wire v$C7_16434_out0;
wire v$C7_338_out0;
wire v$C7_339_out0;
wire v$C7_9496_out0;
wire v$C8_18497_out0;
wire v$C8_18498_out0;
wire v$C8_18499_out0;
wire v$C8_18500_out0;
wire v$C8_18501_out0;
wire v$C8_7430_out0;
wire v$C8_7431_out0;
wire v$C8_7432_out0;
wire v$C8_7433_out0;
wire v$C8_7434_out0;
wire v$C9_12155_out0;
wire v$C9_12156_out0;
wire v$C9_12157_out0;
wire v$C9_12158_out0;
wire v$C9_12159_out0;
wire v$C9_5937_out0;
wire v$C9_5938_out0;
wire v$C9_5939_out0;
wire v$C9_5940_out0;
wire v$C9_5941_out0;
wire v$CALCULATING_1493_out0;
wire v$CALCULATING_7798_out0;
wire v$CAPTURE_242_out0;
wire v$CAPTURE_243_out0;
wire v$CARRY_10908_out0;
wire v$CARRY_10909_out0;
wire v$CARRY_13442_out0;
wire v$CARRY_13443_out0;
wire v$CARRY_5003_out0;
wire v$CARRY_5004_out0;
wire v$CARRY_6332_out0;
wire v$CARRY_6333_out0;
wire v$CARRY_6334_out0;
wire v$CARRY_6335_out0;
wire v$CARRY_6336_out0;
wire v$CHECKPARITY_1327_out0;
wire v$CHECKPARITY_1328_out0;
wire v$CIN$EXEC1_1591_out0;
wire v$CINA_8464_out0;
wire v$CINA_8465_out0;
wire v$CINA_8466_out0;
wire v$CINA_8467_out0;
wire v$CINA_8468_out0;
wire v$CINA_8469_out0;
wire v$CINA_8470_out0;
wire v$CINA_8471_out0;
wire v$CINA_8472_out0;
wire v$CINA_8473_out0;
wire v$CINA_8474_out0;
wire v$CINA_8475_out0;
wire v$CINA_8476_out0;
wire v$CINA_8477_out0;
wire v$CINA_8478_out0;
wire v$CINA_8479_out0;
wire v$CINA_8480_out0;
wire v$CINA_8481_out0;
wire v$CINA_8482_out0;
wire v$CINA_8483_out0;
wire v$CINA_8484_out0;
wire v$CINA_8485_out0;
wire v$CINA_8486_out0;
wire v$CINA_8487_out0;
wire v$CINA_8488_out0;
wire v$CINA_8489_out0;
wire v$CINA_8490_out0;
wire v$CINA_8491_out0;
wire v$CINA_8492_out0;
wire v$CINA_8493_out0;
wire v$CINA_8494_out0;
wire v$CINA_8495_out0;
wire v$CINA_8496_out0;
wire v$CINA_8497_out0;
wire v$CINA_8498_out0;
wire v$CINA_8499_out0;
wire v$CINA_8500_out0;
wire v$CINA_8501_out0;
wire v$CINA_8502_out0;
wire v$CINA_8503_out0;
wire v$CINA_8504_out0;
wire v$CINA_8505_out0;
wire v$CINA_8506_out0;
wire v$CINA_8507_out0;
wire v$CINA_8508_out0;
wire v$CINA_8509_out0;
wire v$CINA_8510_out0;
wire v$CINA_8511_out0;
wire v$CINA_8512_out0;
wire v$CINA_8513_out0;
wire v$CINA_8514_out0;
wire v$CINA_8515_out0;
wire v$CINA_8516_out0;
wire v$CINA_8517_out0;
wire v$CINA_8518_out0;
wire v$CINA_8519_out0;
wire v$CINA_8520_out0;
wire v$CINA_8521_out0;
wire v$CINA_8522_out0;
wire v$CINA_8523_out0;
wire v$CINA_8524_out0;
wire v$CINA_8525_out0;
wire v$CINA_8526_out0;
wire v$CINA_8527_out0;
wire v$CINA_8528_out0;
wire v$CINA_8529_out0;
wire v$CINA_8530_out0;
wire v$CINA_8531_out0;
wire v$CINA_8532_out0;
wire v$CINA_8533_out0;
wire v$CINA_8534_out0;
wire v$CINA_8535_out0;
wire v$CINA_8536_out0;
wire v$CINA_8537_out0;
wire v$CINA_8538_out0;
wire v$CINA_8539_out0;
wire v$CINA_8540_out0;
wire v$CINA_8541_out0;
wire v$CINA_8542_out0;
wire v$CINA_8543_out0;
wire v$CINA_8544_out0;
wire v$CINA_8545_out0;
wire v$CINA_8546_out0;
wire v$CINA_8547_out0;
wire v$CINA_8548_out0;
wire v$CINA_8549_out0;
wire v$CINA_8550_out0;
wire v$CINA_8551_out0;
wire v$CINA_8552_out0;
wire v$CINA_8553_out0;
wire v$CINA_8554_out0;
wire v$CINA_8555_out0;
wire v$CINA_8556_out0;
wire v$CINA_8557_out0;
wire v$CINA_8558_out0;
wire v$CINA_8559_out0;
wire v$CINA_8560_out0;
wire v$CINA_8561_out0;
wire v$CINA_8562_out0;
wire v$CINA_8563_out0;
wire v$CINA_8564_out0;
wire v$CINA_8565_out0;
wire v$CINA_8566_out0;
wire v$CINA_8567_out0;
wire v$CINA_8568_out0;
wire v$CINA_8569_out0;
wire v$CINA_8570_out0;
wire v$CINA_8571_out0;
wire v$CINA_8572_out0;
wire v$CINA_8573_out0;
wire v$CINA_8574_out0;
wire v$CINA_8575_out0;
wire v$CINA_8576_out0;
wire v$CINA_8577_out0;
wire v$CINA_8578_out0;
wire v$CINA_8579_out0;
wire v$CINA_8580_out0;
wire v$CINA_8581_out0;
wire v$CINA_8582_out0;
wire v$CINA_8583_out0;
wire v$CINA_8584_out0;
wire v$CINA_8585_out0;
wire v$CINA_8586_out0;
wire v$CINA_8587_out0;
wire v$CINA_8588_out0;
wire v$CINA_8589_out0;
wire v$CINA_8590_out0;
wire v$CINA_8591_out0;
wire v$CINA_8592_out0;
wire v$CINA_8593_out0;
wire v$CINA_8594_out0;
wire v$CINA_8595_out0;
wire v$CINA_8596_out0;
wire v$CINA_8597_out0;
wire v$CINA_8598_out0;
wire v$CINA_8599_out0;
wire v$CINA_8600_out0;
wire v$CINA_8601_out0;
wire v$CINA_8602_out0;
wire v$CINA_8603_out0;
wire v$CINA_8604_out0;
wire v$CINA_8605_out0;
wire v$CINA_8606_out0;
wire v$CINA_8607_out0;
wire v$CINA_8608_out0;
wire v$CINA_8609_out0;
wire v$CINA_8610_out0;
wire v$CINA_8611_out0;
wire v$CINA_8612_out0;
wire v$CINA_8613_out0;
wire v$CINA_8614_out0;
wire v$CINA_8615_out0;
wire v$CINA_8616_out0;
wire v$CINA_8617_out0;
wire v$CINA_8618_out0;
wire v$CINA_8619_out0;
wire v$CINA_8620_out0;
wire v$CINA_8621_out0;
wire v$CINA_8622_out0;
wire v$CINA_8623_out0;
wire v$CINA_8624_out0;
wire v$CINA_8625_out0;
wire v$CINA_8626_out0;
wire v$CINA_8627_out0;
wire v$CINA_8628_out0;
wire v$CINA_8629_out0;
wire v$CINA_8630_out0;
wire v$CINA_8631_out0;
wire v$CINA_8632_out0;
wire v$CINA_8633_out0;
wire v$CINA_8634_out0;
wire v$CINA_8635_out0;
wire v$CINA_8636_out0;
wire v$CINA_8637_out0;
wire v$CINA_8638_out0;
wire v$CINA_8639_out0;
wire v$CINA_8640_out0;
wire v$CINA_8641_out0;
wire v$CINA_8642_out0;
wire v$CINA_8643_out0;
wire v$CINA_8644_out0;
wire v$CINA_8645_out0;
wire v$CINA_8646_out0;
wire v$CINA_8647_out0;
wire v$CINA_8648_out0;
wire v$CINA_8649_out0;
wire v$CINA_8650_out0;
wire v$CINA_8651_out0;
wire v$CINA_8652_out0;
wire v$CINA_8653_out0;
wire v$CINA_8654_out0;
wire v$CINA_8655_out0;
wire v$CINA_8656_out0;
wire v$CINA_8657_out0;
wire v$CINA_8658_out0;
wire v$CINA_8659_out0;
wire v$CINA_8660_out0;
wire v$CINA_8661_out0;
wire v$CINA_8662_out0;
wire v$CINA_8663_out0;
wire v$CINA_8664_out0;
wire v$CINA_8665_out0;
wire v$CINA_8666_out0;
wire v$CINA_8667_out0;
wire v$CINA_8668_out0;
wire v$CIN_15050_out0;
wire v$CIN_15051_out0;
wire v$CIN_15052_out0;
wire v$CIN_15053_out0;
wire v$CIN_15054_out0;
wire v$CIN_16106_out0;
wire v$CIN_16107_out0;
wire v$CIN_16108_out0;
wire v$CIN_16109_out0;
wire v$CIN_16110_out0;
wire v$CIN_16812_out0;
wire v$CIN_16813_out0;
wire v$CIN_16814_out0;
wire v$CIN_16815_out0;
wire v$CIN_16816_out0;
wire v$CIN_16817_out0;
wire v$CIN_16818_out0;
wire v$CIN_16819_out0;
wire v$CIN_16820_out0;
wire v$CIN_16821_out0;
wire v$CIN_16822_out0;
wire v$CIN_16823_out0;
wire v$CIN_17342_out0;
wire v$CIN_17343_out0;
wire v$CIN_17344_out0;
wire v$CIN_17345_out0;
wire v$CIN_17346_out0;
wire v$CIN_18225_out0;
wire v$CIN_18226_out0;
wire v$CIN_18227_out0;
wire v$CIN_18228_out0;
wire v$CIN_18229_out0;
wire v$CIN_18230_out0;
wire v$CIN_18231_out0;
wire v$CIN_18232_out0;
wire v$CIN_3886_out0;
wire v$CIN_3887_out0;
wire v$CIN_3888_out0;
wire v$CIN_3889_out0;
wire v$CIN_3890_out0;
wire v$CIN_3891_out0;
wire v$CIN_3892_out0;
wire v$CIN_3893_out0;
wire v$CIN_3894_out0;
wire v$CIN_3895_out0;
wire v$CIN_3896_out0;
wire v$CIN_3897_out0;
wire v$CLEAR_18404_out0;
wire v$CLEAR_18405_out0;
wire v$CLK4_12213_out0;
wire v$CLK4_12214_out0;
wire v$CLK4_16733_out0;
wire v$CLK4_16734_out0;
wire v$CLK4_17983_out0;
wire v$CLK4_17984_out0;
wire v$CLK4_2531_out0;
wire v$CLK4_2532_out0;
wire v$CLK4_3694_out0;
wire v$CLK4_3695_out0;
wire v$CLK4_7060_out0;
wire v$CLK4_7061_out0;
wire v$CLK4_8834_out0;
wire v$CLK4_8835_out0;
wire v$CLRINTERRUPTS_340_out0;
wire v$CLRINTERRUPTS_341_out0;
wire v$CLR_4434_out0;
wire v$CLR_4435_out0;
wire v$COMP$H$OUT_6646_out0;
wire v$COMP$H$OUT_6647_out0;
wire v$COMP$L$OUT_11695_out0;
wire v$COMP$L$OUT_11696_out0;
wire v$CON1_4080_out0;
wire v$CON1_4081_out0;
wire v$CON1_4082_out0;
wire v$CON1_4083_out0;
wire v$CON1_4084_out0;
wire v$CON2_14367_out0;
wire v$CON2_14368_out0;
wire v$CON2_14369_out0;
wire v$CON2_14370_out0;
wire v$CON2_14371_out0;
wire v$CON3_7912_out0;
wire v$CON3_7913_out0;
wire v$CON3_7914_out0;
wire v$CON3_7915_out0;
wire v$CON3_7916_out0;
wire v$CON4_16435_out0;
wire v$CON4_16436_out0;
wire v$CON4_16437_out0;
wire v$CON4_16438_out0;
wire v$CON4_16439_out0;
wire v$CON5_10681_out0;
wire v$CON5_10682_out0;
wire v$CON5_10683_out0;
wire v$CON5_10684_out0;
wire v$CON5_10685_out0;
wire v$CON6_12997_out0;
wire v$CON6_12998_out0;
wire v$CON6_12999_out0;
wire v$CON6_13000_out0;
wire v$CON6_13001_out0;
wire v$CON7_2420_out0;
wire v$CON7_2421_out0;
wire v$CON7_2422_out0;
wire v$CON7_2423_out0;
wire v$CON7_2424_out0;
wire v$COUNTEREN_13450_out0;
wire v$COUNTEREN_13451_out0;
wire v$COUNTEREN_1625_out0;
wire v$COUNTEREN_1626_out0;
wire v$COUNTERINTERRUPT_14849_out0;
wire v$COUNTERINTERRUPT_14850_out0;
wire v$COUT$EXEC1_1594_out0;
wire v$COUT$HALF_72_out0;
wire v$COUT1_7469_out0;
wire v$COUTD_6693_out0;
wire v$COUTD_6694_out0;
wire v$COUTD_6695_out0;
wire v$COUTD_6696_out0;
wire v$COUTD_6697_out0;
wire v$COUTD_6698_out0;
wire v$COUTD_6699_out0;
wire v$COUTD_6700_out0;
wire v$COUTD_6701_out0;
wire v$COUTD_6702_out0;
wire v$COUTD_6703_out0;
wire v$COUTD_6704_out0;
wire v$COUTD_6705_out0;
wire v$COUTD_6706_out0;
wire v$COUTD_6707_out0;
wire v$COUTD_6708_out0;
wire v$COUTD_6709_out0;
wire v$COUTD_6710_out0;
wire v$COUTD_6711_out0;
wire v$COUTD_6712_out0;
wire v$COUTD_6713_out0;
wire v$COUTD_6714_out0;
wire v$COUTD_6715_out0;
wire v$COUTD_6716_out0;
wire v$COUTD_6717_out0;
wire v$COUTD_6718_out0;
wire v$COUTD_6719_out0;
wire v$COUTD_6720_out0;
wire v$COUTD_6721_out0;
wire v$COUTD_6722_out0;
wire v$COUTD_6723_out0;
wire v$COUTD_6724_out0;
wire v$COUTD_6725_out0;
wire v$COUTD_6726_out0;
wire v$COUTD_6727_out0;
wire v$COUTD_6728_out0;
wire v$COUTD_6729_out0;
wire v$COUTD_6730_out0;
wire v$COUTD_6731_out0;
wire v$COUTD_6732_out0;
wire v$COUTD_6733_out0;
wire v$COUTD_6734_out0;
wire v$COUTD_6735_out0;
wire v$COUTD_6736_out0;
wire v$COUTD_6737_out0;
wire v$COUTD_6738_out0;
wire v$COUTD_6739_out0;
wire v$COUTD_6740_out0;
wire v$COUTD_6741_out0;
wire v$COUTD_6742_out0;
wire v$COUTD_6743_out0;
wire v$COUTD_6744_out0;
wire v$COUTD_6745_out0;
wire v$COUTD_6746_out0;
wire v$COUTD_6747_out0;
wire v$COUTD_6748_out0;
wire v$COUTD_6749_out0;
wire v$COUTD_6750_out0;
wire v$COUTD_6751_out0;
wire v$COUTD_6752_out0;
wire v$COUTD_6753_out0;
wire v$COUTD_6754_out0;
wire v$COUTD_6755_out0;
wire v$COUTD_6756_out0;
wire v$COUTD_6757_out0;
wire v$COUTD_6758_out0;
wire v$COUTD_6759_out0;
wire v$COUTD_6760_out0;
wire v$COUTD_6761_out0;
wire v$COUTD_6762_out0;
wire v$COUTD_6763_out0;
wire v$COUTD_6764_out0;
wire v$COUTD_6765_out0;
wire v$COUTD_6766_out0;
wire v$COUTD_6767_out0;
wire v$COUTD_6768_out0;
wire v$COUTD_6769_out0;
wire v$COUTD_6770_out0;
wire v$COUTD_6771_out0;
wire v$COUTD_6772_out0;
wire v$COUTD_6773_out0;
wire v$COUTD_6774_out0;
wire v$COUTD_6775_out0;
wire v$COUTD_6776_out0;
wire v$COUTD_6777_out0;
wire v$COUTD_6778_out0;
wire v$COUTD_6779_out0;
wire v$COUTD_6780_out0;
wire v$COUTD_6781_out0;
wire v$COUTD_6782_out0;
wire v$COUTD_6783_out0;
wire v$COUTD_6784_out0;
wire v$COUTD_6785_out0;
wire v$COUTD_6786_out0;
wire v$COUTD_6787_out0;
wire v$COUTD_6788_out0;
wire v$COUTD_6789_out0;
wire v$COUTD_6790_out0;
wire v$COUTD_6791_out0;
wire v$COUTD_6792_out0;
wire v$COUTD_6793_out0;
wire v$COUTD_6794_out0;
wire v$COUTD_6795_out0;
wire v$COUTD_6796_out0;
wire v$COUTD_6797_out0;
wire v$COUTD_6798_out0;
wire v$COUTD_6799_out0;
wire v$COUTD_6800_out0;
wire v$COUTD_6801_out0;
wire v$COUTD_6802_out0;
wire v$COUTD_6803_out0;
wire v$COUTD_6804_out0;
wire v$COUTD_6805_out0;
wire v$COUTD_6806_out0;
wire v$COUTD_6807_out0;
wire v$COUTD_6808_out0;
wire v$COUTD_6809_out0;
wire v$COUTD_6810_out0;
wire v$COUTD_6811_out0;
wire v$COUTD_6812_out0;
wire v$COUTD_6813_out0;
wire v$COUTD_6814_out0;
wire v$COUTD_6815_out0;
wire v$COUTD_6816_out0;
wire v$COUTD_6817_out0;
wire v$COUTD_6818_out0;
wire v$COUTD_6819_out0;
wire v$COUTD_6820_out0;
wire v$COUTD_6821_out0;
wire v$COUTD_6822_out0;
wire v$COUTD_6823_out0;
wire v$COUTD_6824_out0;
wire v$COUTD_6825_out0;
wire v$COUTD_6826_out0;
wire v$COUTD_6827_out0;
wire v$COUTD_6828_out0;
wire v$COUTD_6829_out0;
wire v$COUTD_6830_out0;
wire v$COUTD_6831_out0;
wire v$COUTD_6832_out0;
wire v$COUTD_6833_out0;
wire v$COUTD_6834_out0;
wire v$COUTD_6835_out0;
wire v$COUTD_6836_out0;
wire v$COUTD_6837_out0;
wire v$COUTD_6838_out0;
wire v$COUTD_6839_out0;
wire v$COUTD_6840_out0;
wire v$COUTD_6841_out0;
wire v$COUTD_6842_out0;
wire v$COUTD_6843_out0;
wire v$COUTD_6844_out0;
wire v$COUTD_6845_out0;
wire v$COUTD_6846_out0;
wire v$COUTD_6847_out0;
wire v$COUTD_6848_out0;
wire v$COUTD_6849_out0;
wire v$COUTD_6850_out0;
wire v$COUTD_6851_out0;
wire v$COUTD_6852_out0;
wire v$COUTD_6853_out0;
wire v$COUTD_6854_out0;
wire v$COUTD_6855_out0;
wire v$COUTD_6856_out0;
wire v$COUTD_6857_out0;
wire v$COUTD_6858_out0;
wire v$COUTD_6859_out0;
wire v$COUTD_6860_out0;
wire v$COUTD_6861_out0;
wire v$COUTD_6862_out0;
wire v$COUTD_6863_out0;
wire v$COUTD_6864_out0;
wire v$COUTD_6865_out0;
wire v$COUTD_6866_out0;
wire v$COUTD_6867_out0;
wire v$COUTD_6868_out0;
wire v$COUTD_6869_out0;
wire v$COUTD_6870_out0;
wire v$COUTD_6871_out0;
wire v$COUTD_6872_out0;
wire v$COUTD_6873_out0;
wire v$COUTD_6874_out0;
wire v$COUTD_6875_out0;
wire v$COUTD_6876_out0;
wire v$COUTD_6877_out0;
wire v$COUTD_6878_out0;
wire v$COUTD_6879_out0;
wire v$COUTD_6880_out0;
wire v$COUTD_6881_out0;
wire v$COUTD_6882_out0;
wire v$COUTD_6883_out0;
wire v$COUTD_6884_out0;
wire v$COUTD_6885_out0;
wire v$COUTD_6886_out0;
wire v$COUTD_6887_out0;
wire v$COUTD_6888_out0;
wire v$COUTD_6889_out0;
wire v$COUTD_6890_out0;
wire v$COUTD_6891_out0;
wire v$COUTD_6892_out0;
wire v$COUTD_6893_out0;
wire v$COUTD_6894_out0;
wire v$COUTD_6895_out0;
wire v$COUTD_6896_out0;
wire v$COUTD_6897_out0;
wire v$COUT_10728_out0;
wire v$COUT_10729_out0;
wire v$COUT_10730_out0;
wire v$COUT_10731_out0;
wire v$COUT_10732_out0;
wire v$COUT_10733_out0;
wire v$COUT_10734_out0;
wire v$COUT_10735_out0;
wire v$COUT_10736_out0;
wire v$COUT_10737_out0;
wire v$COUT_10738_out0;
wire v$COUT_10739_out0;
wire v$COUT_13515_out0;
wire v$COUT_5015_out0;
wire v$COUT_8111_out0;
wire v$COUT_8112_out0;
wire v$COUT_8113_out0;
wire v$COUT_8114_out0;
wire v$COUT_8115_out0;
wire v$COUT_8116_out0;
wire v$COUT_8117_out0;
wire v$COUT_8118_out0;
wire v$COUT_8119_out0;
wire v$COUT_8120_out0;
wire v$COUT_8121_out0;
wire v$COUT_8122_out0;
wire v$COUT_8292_out0;
wire v$COUT_8293_out0;
wire v$C_15895_out0;
wire v$C_15896_out0;
wire v$C_3198_out0;
wire v$C_3199_out0;
wire v$C_3641_out0;
wire v$C_3642_out0;
wire v$C_6062_out0;
wire v$C_6063_out0;
wire v$C_9609_out0;
wire v$C_9610_out0;
wire v$CheckParity_18678_out0;
wire v$CheckParity_18679_out0;
wire v$Clear_12750_out0;
wire v$Clear_12751_out0;
wire v$Clear_14641_out0;
wire v$Clear_14642_out0;
wire v$D1_14097_out0;
wire v$D1_14097_out1;
wire v$D1_14097_out2;
wire v$D1_14097_out3;
wire v$D1_14098_out0;
wire v$D1_14098_out1;
wire v$D1_14098_out2;
wire v$D1_14098_out3;
wire v$DATA$DEPENDENCY_6157_out0;
wire v$DATA$DEPENDENCY_6158_out0;
wire v$DATA$PROCESS$WB_17832_out0;
wire v$DATA$PROCESS$WB_17833_out0;
wire v$DISABLEINTERRUPTS_14974_out0;
wire v$DISABLEINTERRUPTS_14975_out0;
wire v$DM1_16244_out0;
wire v$DM1_16244_out1;
wire v$EDGE0_3990_out0;
wire v$EDGE0_3991_out0;
wire v$EDGE0_5740_out0;
wire v$EDGE0_5741_out0;
wire v$EDGE1_15272_out0;
wire v$EDGE1_15273_out0;
wire v$EDGE1_17407_out0;
wire v$EDGE1_17408_out0;
wire v$EDGE2_18118_out0;
wire v$EDGE2_18119_out0;
wire v$EDGE2_6999_out0;
wire v$EDGE2_7000_out0;
wire v$EDGE3_11040_out0;
wire v$EDGE3_11041_out0;
wire v$EDGE3_2241_out0;
wire v$EDGE3_2242_out0;
wire v$ENABLEINTERRUPTS_12547_out0;
wire v$ENABLEINTERRUPTS_12548_out0;
wire v$ENABLEINTERRUPTS_17026_out0;
wire v$ENABLEINTERRUPTS_17027_out0;
wire v$ENCODED0_14022_out0;
wire v$ENCODED0_14023_out0;
wire v$ENCODED1_9520_out0;
wire v$ENCODED1_9521_out0;
wire v$END0_9352_out0;
wire v$END0_9353_out0;
wire v$END0_9354_out0;
wire v$END0_9355_out0;
wire v$END0_9356_out0;
wire v$END10_1151_out0;
wire v$END10_1152_out0;
wire v$END10_1153_out0;
wire v$END10_1154_out0;
wire v$END10_1155_out0;
wire v$END11_12090_out0;
wire v$END11_12091_out0;
wire v$END11_12092_out0;
wire v$END11_12093_out0;
wire v$END11_12094_out0;
wire v$END12_10780_out0;
wire v$END12_10781_out0;
wire v$END12_10782_out0;
wire v$END12_10783_out0;
wire v$END12_10784_out0;
wire v$END13_18067_out0;
wire v$END13_18068_out0;
wire v$END13_18069_out0;
wire v$END13_18070_out0;
wire v$END13_18071_out0;
wire v$END14_274_out0;
wire v$END14_275_out0;
wire v$END14_276_out0;
wire v$END14_277_out0;
wire v$END14_278_out0;
wire v$END15_7382_out0;
wire v$END15_7383_out0;
wire v$END15_7384_out0;
wire v$END15_7385_out0;
wire v$END15_7386_out0;
wire v$END16_216_out0;
wire v$END16_217_out0;
wire v$END16_218_out0;
wire v$END16_219_out0;
wire v$END16_220_out0;
wire v$END17_7637_out0;
wire v$END17_7638_out0;
wire v$END17_7639_out0;
wire v$END17_7640_out0;
wire v$END17_7641_out0;
wire v$END18_11946_out0;
wire v$END18_11947_out0;
wire v$END18_11948_out0;
wire v$END18_11949_out0;
wire v$END18_11950_out0;
wire v$END19_11655_out0;
wire v$END19_11656_out0;
wire v$END19_11657_out0;
wire v$END19_11658_out0;
wire v$END19_11659_out0;
wire v$END1_1291_out0;
wire v$END1_1292_out0;
wire v$END1_1293_out0;
wire v$END1_1294_out0;
wire v$END1_1295_out0;
wire v$END1_1543_out0;
wire v$END1_1544_out0;
wire v$END1_1545_out0;
wire v$END1_1546_out0;
wire v$END1_1547_out0;
wire v$END1_6960_out0;
wire v$END1_6961_out0;
wire v$END1_6986_out0;
wire v$END1_6987_out0;
wire v$END20_13264_out0;
wire v$END20_13265_out0;
wire v$END20_13266_out0;
wire v$END20_13267_out0;
wire v$END20_13268_out0;
wire v$END21_4340_out0;
wire v$END21_4341_out0;
wire v$END21_4342_out0;
wire v$END21_4343_out0;
wire v$END21_4344_out0;
wire v$END22_15484_out0;
wire v$END22_15485_out0;
wire v$END22_15486_out0;
wire v$END22_15487_out0;
wire v$END22_15488_out0;
wire v$END23_16717_out0;
wire v$END23_16718_out0;
wire v$END23_16719_out0;
wire v$END23_16720_out0;
wire v$END23_16721_out0;
wire v$END24_16403_out0;
wire v$END24_16404_out0;
wire v$END24_16405_out0;
wire v$END24_16406_out0;
wire v$END24_16407_out0;
wire v$END25_17070_out0;
wire v$END25_17071_out0;
wire v$END25_17072_out0;
wire v$END25_17073_out0;
wire v$END25_17074_out0;
wire v$END26_6435_out0;
wire v$END26_6436_out0;
wire v$END26_6437_out0;
wire v$END26_6438_out0;
wire v$END26_6439_out0;
wire v$END27_2210_out0;
wire v$END27_2211_out0;
wire v$END27_2212_out0;
wire v$END27_2213_out0;
wire v$END27_2214_out0;
wire v$END28_13669_out0;
wire v$END28_13670_out0;
wire v$END28_13671_out0;
wire v$END28_13672_out0;
wire v$END28_13673_out0;
wire v$END29_5885_out0;
wire v$END29_5886_out0;
wire v$END29_5887_out0;
wire v$END29_5888_out0;
wire v$END29_5889_out0;
wire v$END2_5234_out0;
wire v$END2_5235_out0;
wire v$END2_5236_out0;
wire v$END2_5237_out0;
wire v$END2_5238_out0;
wire v$END2_7751_out0;
wire v$END2_7752_out0;
wire v$END2_7753_out0;
wire v$END2_7754_out0;
wire v$END2_7755_out0;
wire v$END30_15713_out0;
wire v$END30_15714_out0;
wire v$END30_15715_out0;
wire v$END30_15716_out0;
wire v$END30_15717_out0;
wire v$END31_18520_out0;
wire v$END31_18521_out0;
wire v$END31_18522_out0;
wire v$END31_18523_out0;
wire v$END31_18524_out0;
wire v$END32_2470_out0;
wire v$END32_2471_out0;
wire v$END32_2472_out0;
wire v$END32_2473_out0;
wire v$END32_2474_out0;
wire v$END33_264_out0;
wire v$END33_265_out0;
wire v$END33_266_out0;
wire v$END33_267_out0;
wire v$END33_268_out0;
wire v$END3_3445_out0;
wire v$END3_3446_out0;
wire v$END3_3447_out0;
wire v$END3_3448_out0;
wire v$END3_3449_out0;
wire v$END3_7932_out0;
wire v$END3_7933_out0;
wire v$END3_7934_out0;
wire v$END3_7935_out0;
wire v$END3_7936_out0;
wire v$END40_5775_out0;
wire v$END40_5776_out0;
wire v$END40_5777_out0;
wire v$END40_5778_out0;
wire v$END40_5779_out0;
wire v$END41_16665_out0;
wire v$END41_16666_out0;
wire v$END41_16667_out0;
wire v$END41_16668_out0;
wire v$END41_16669_out0;
wire v$END42_18311_out0;
wire v$END42_18312_out0;
wire v$END42_18313_out0;
wire v$END42_18314_out0;
wire v$END42_18315_out0;
wire v$END43_13192_out0;
wire v$END43_13193_out0;
wire v$END43_13194_out0;
wire v$END43_13195_out0;
wire v$END43_13196_out0;
wire v$END44_15665_out0;
wire v$END44_15666_out0;
wire v$END44_15667_out0;
wire v$END44_15668_out0;
wire v$END44_15669_out0;
wire v$END45_9057_out0;
wire v$END45_9058_out0;
wire v$END45_9059_out0;
wire v$END45_9060_out0;
wire v$END45_9061_out0;
wire v$END46_15045_out0;
wire v$END46_15046_out0;
wire v$END46_15047_out0;
wire v$END46_15048_out0;
wire v$END46_15049_out0;
wire v$END47_2679_out0;
wire v$END47_2680_out0;
wire v$END47_2681_out0;
wire v$END47_2682_out0;
wire v$END47_2683_out0;
wire v$END48_10365_out0;
wire v$END48_10366_out0;
wire v$END48_10367_out0;
wire v$END48_10368_out0;
wire v$END48_10369_out0;
wire v$END49_18450_out0;
wire v$END49_18451_out0;
wire v$END49_18452_out0;
wire v$END49_18453_out0;
wire v$END49_18454_out0;
wire v$END4_3267_out0;
wire v$END4_3268_out0;
wire v$END4_5246_out0;
wire v$END4_5247_out0;
wire v$END4_5248_out0;
wire v$END4_5249_out0;
wire v$END4_5250_out0;
wire v$END4_8128_out0;
wire v$END4_8129_out0;
wire v$END4_9367_out0;
wire v$END4_9368_out0;
wire v$END4_9369_out0;
wire v$END4_9370_out0;
wire v$END4_9371_out0;
wire v$END50_7413_out0;
wire v$END50_7414_out0;
wire v$END50_7415_out0;
wire v$END50_7416_out0;
wire v$END50_7417_out0;
wire v$END51_11676_out0;
wire v$END51_11677_out0;
wire v$END51_11678_out0;
wire v$END51_11679_out0;
wire v$END51_11680_out0;
wire v$END52_11973_out0;
wire v$END52_11974_out0;
wire v$END52_11975_out0;
wire v$END52_11976_out0;
wire v$END52_11977_out0;
wire v$END53_317_out0;
wire v$END53_318_out0;
wire v$END53_319_out0;
wire v$END53_320_out0;
wire v$END53_321_out0;
wire v$END5_4143_out0;
wire v$END5_4144_out0;
wire v$END5_4145_out0;
wire v$END5_4146_out0;
wire v$END5_4147_out0;
wire v$END60_15132_out0;
wire v$END60_15133_out0;
wire v$END60_15134_out0;
wire v$END60_15135_out0;
wire v$END60_15136_out0;
wire v$END61_17956_out0;
wire v$END61_17957_out0;
wire v$END61_17958_out0;
wire v$END61_17959_out0;
wire v$END61_17960_out0;
wire v$END6_15249_out0;
wire v$END6_15250_out0;
wire v$END6_15251_out0;
wire v$END6_15252_out0;
wire v$END6_15253_out0;
wire v$END6_7544_out0;
wire v$END6_7545_out0;
wire v$END7_3359_out0;
wire v$END7_3360_out0;
wire v$END7_3361_out0;
wire v$END7_3362_out0;
wire v$END7_3363_out0;
wire v$END8_3901_out0;
wire v$END8_3902_out0;
wire v$END8_3903_out0;
wire v$END8_3904_out0;
wire v$END8_3905_out0;
wire v$END9_4233_out0;
wire v$END9_4234_out0;
wire v$END9_4235_out0;
wire v$END9_4236_out0;
wire v$END9_4237_out0;
wire v$END_15738_out0;
wire v$END_15739_out0;
wire v$END_17049_out0;
wire v$END_17050_out0;
wire v$END_18272_out0;
wire v$END_18273_out0;
wire v$END_18274_out0;
wire v$END_18275_out0;
wire v$END_18276_out0;
wire v$END_3319_out0;
wire v$END_3320_out0;
wire v$END_3321_out0;
wire v$END_3322_out0;
wire v$END_3323_out0;
wire v$END_8096_out0;
wire v$END_8097_out0;
wire v$ENDa_16564_out0;
wire v$ENDa_16565_out0;
wire v$ENDa_16566_out0;
wire v$ENDa_16567_out0;
wire v$ENDa_16568_out0;
wire v$ENDd_10832_out0;
wire v$ENDd_10833_out0;
wire v$ENDd_10834_out0;
wire v$ENDd_10835_out0;
wire v$ENDd_10836_out0;
wire v$ENDe_17892_out0;
wire v$ENDe_17893_out0;
wire v$ENDe_17894_out0;
wire v$ENDe_17895_out0;
wire v$ENDe_17896_out0;
wire v$ENDi_8682_out0;
wire v$ENDi_8683_out0;
wire v$ENDi_8684_out0;
wire v$ENDi_8685_out0;
wire v$ENDi_8686_out0;
wire v$ENDo_18692_out0;
wire v$ENDo_18693_out0;
wire v$ENDo_18694_out0;
wire v$ENDo_18695_out0;
wire v$ENDo_18696_out0;
wire v$ENDp_3189_out0;
wire v$ENDp_3190_out0;
wire v$ENDp_3191_out0;
wire v$ENDp_3192_out0;
wire v$ENDp_3193_out0;
wire v$ENDq_1458_out0;
wire v$ENDq_1459_out0;
wire v$ENDq_1460_out0;
wire v$ENDq_1461_out0;
wire v$ENDq_1462_out0;
wire v$ENDr_7522_out0;
wire v$ENDr_7523_out0;
wire v$ENDr_7524_out0;
wire v$ENDr_7525_out0;
wire v$ENDr_7526_out0;
wire v$ENDs_3213_out0;
wire v$ENDs_3214_out0;
wire v$ENDs_3215_out0;
wire v$ENDs_3216_out0;
wire v$ENDs_3217_out0;
wire v$ENDt_10258_out0;
wire v$ENDt_10259_out0;
wire v$ENDt_10260_out0;
wire v$ENDt_10261_out0;
wire v$ENDt_10262_out0;
wire v$ENDu_7029_out0;
wire v$ENDu_7030_out0;
wire v$ENDu_7031_out0;
wire v$ENDu_7032_out0;
wire v$ENDu_7033_out0;
wire v$ENDw_9551_out0;
wire v$ENDw_9552_out0;
wire v$ENDw_9553_out0;
wire v$ENDw_9554_out0;
wire v$ENDw_9555_out0;
wire v$ENDy_4114_out0;
wire v$ENDy_4115_out0;
wire v$ENDy_4116_out0;
wire v$ENDy_4117_out0;
wire v$ENDy_4118_out0;
wire v$ENMODE_14574_out0;
wire v$ENMODE_14575_out0;
wire v$ENMODE_7737_out0;
wire v$ENMODE_7738_out0;
wire v$EN_1331_out0;
wire v$EN_1332_out0;
wire v$EN_1333_out0;
wire v$EN_1334_out0;
wire v$EN_1335_out0;
wire v$EN_1336_out0;
wire v$EN_1337_out0;
wire v$EN_1338_out0;
wire v$EN_1339_out0;
wire v$EN_1340_out0;
wire v$EN_1341_out0;
wire v$EN_1342_out0;
wire v$EN_1343_out0;
wire v$EN_1344_out0;
wire v$EN_1345_out0;
wire v$EN_1346_out0;
wire v$EN_1347_out0;
wire v$EN_1348_out0;
wire v$EN_1349_out0;
wire v$EN_1350_out0;
wire v$EN_15897_out0;
wire v$EN_15898_out0;
wire v$EN_16385_out0;
wire v$EN_16386_out0;
wire v$EN_16387_out0;
wire v$EN_16388_out0;
wire v$EN_16389_out0;
wire v$EN_16390_out0;
wire v$EN_16391_out0;
wire v$EN_16392_out0;
wire v$EN_16965_out0;
wire v$EN_16966_out0;
wire v$EN_16967_out0;
wire v$EN_16968_out0;
wire v$EN_16969_out0;
wire v$EN_16970_out0;
wire v$EN_16971_out0;
wire v$EN_16972_out0;
wire v$EN_3875_out0;
wire v$EN_3876_out0;
wire v$EN_3877_out0;
wire v$EN_4751_out0;
wire v$EN_4752_out0;
wire v$EN_4753_out0;
wire v$EN_4754_out0;
wire v$EN_4755_out0;
wire v$EN_4756_out0;
wire v$EN_4757_out0;
wire v$EN_4758_out0;
wire v$EN_4759_out0;
wire v$EN_4760_out0;
wire v$EN_4761_out0;
wire v$EN_4762_out0;
wire v$EN_5210_out0;
wire v$EN_5211_out0;
wire v$EN_5212_out0;
wire v$EN_5213_out0;
wire v$EN_5214_out0;
wire v$EN_5215_out0;
wire v$EN_5216_out0;
wire v$EN_5217_out0;
wire v$EN_5218_out0;
wire v$EN_5219_out0;
wire v$EN_5220_out0;
wire v$EN_5221_out0;
wire v$EN_5222_out0;
wire v$EN_5223_out0;
wire v$EN_5224_out0;
wire v$EN_5225_out0;
wire v$EN_7873_out0;
wire v$EN_7874_out0;
wire v$EN_7875_out0;
wire v$EN_7876_out0;
wire v$EN_7877_out0;
wire v$EN_7878_out0;
wire v$EN_7879_out0;
wire v$EN_7880_out0;
wire v$EN_7881_out0;
wire v$EN_7882_out0;
wire v$EN_7883_out0;
wire v$EN_7884_out0;
wire v$EN_9080_out0;
wire v$EN_9081_out0;
wire v$EPARITY_18309_out0;
wire v$EPARITY_18310_out0;
wire v$EQ$LDST_17430_out0;
wire v$EQ$LDST_17431_out0;
wire v$EQ10_13408_out0;
wire v$EQ10_13409_out0;
wire v$EQ10_5892_out0;
wire v$EQ10_5893_out0;
wire v$EQ10_5894_out0;
wire v$EQ10_5895_out0;
wire v$EQ10_9866_out0;
wire v$EQ10_9867_out0;
wire v$EQ11_11882_out0;
wire v$EQ11_11883_out0;
wire v$EQ11_13605_out0;
wire v$EQ11_13606_out0;
wire v$EQ11_6143_out0;
wire v$EQ11_6144_out0;
wire v$EQ11_6145_out0;
wire v$EQ11_6146_out0;
wire v$EQ12_13260_out0;
wire v$EQ12_13261_out0;
wire v$EQ12_13838_out0;
wire v$EQ12_13839_out0;
wire v$EQ12_13840_out0;
wire v$EQ12_13841_out0;
wire v$EQ12_15107_out0;
wire v$EQ12_15108_out0;
wire v$EQ12_1539_out0;
wire v$EQ12_1540_out0;
wire v$EQ13_18548_out0;
wire v$EQ13_18549_out0;
wire v$EQ13_5251_out0;
wire v$EQ13_5252_out0;
wire v$EQ13_9341_out0;
wire v$EQ13_9342_out0;
wire v$EQ13_9515_out0;
wire v$EQ13_9516_out0;
wire v$EQ13_9517_out0;
wire v$EQ13_9518_out0;
wire v$EQ14_12122_out0;
wire v$EQ14_12123_out0;
wire v$EQ14_5401_out0;
wire v$EQ14_5402_out0;
wire v$EQ14_5403_out0;
wire v$EQ14_5404_out0;
wire v$EQ14_5487_out0;
wire v$EQ14_5488_out0;
wire v$EQ15_15790_out0;
wire v$EQ15_15965_out0;
wire v$EQ15_15966_out0;
wire v$EQ15_15967_out0;
wire v$EQ15_15968_out0;
wire v$EQ15_17047_out0;
wire v$EQ15_17048_out0;
wire v$EQ16_10749_out0;
wire v$EQ16_1582_out0;
wire v$EQ16_1583_out0;
wire v$EQ16_8286_out0;
wire v$EQ16_8287_out0;
wire v$EQ16_8288_out0;
wire v$EQ16_8289_out0;
wire v$EQ17_5879_out0;
wire v$EQ17_5880_out0;
wire v$EQ17_5881_out0;
wire v$EQ17_5882_out0;
wire v$EQ18_12806_out0;
wire v$EQ18_12807_out0;
wire v$EQ18_12808_out0;
wire v$EQ18_12809_out0;
wire v$EQ19_5442_out0;
wire v$EQ19_5443_out0;
wire v$EQ19_5444_out0;
wire v$EQ19_5445_out0;
wire v$EQ1_10409_out0;
wire v$EQ1_10410_out0;
wire v$EQ1_11626_out0;
wire v$EQ1_11627_out0;
wire v$EQ1_12945_out0;
wire v$EQ1_12946_out0;
wire v$EQ1_13353_out0;
wire v$EQ1_13354_out0;
wire v$EQ1_13414_out0;
wire v$EQ1_13415_out0;
wire v$EQ1_13416_out0;
wire v$EQ1_13417_out0;
wire v$EQ1_14322_out0;
wire v$EQ1_14323_out0;
wire v$EQ1_15289_out0;
wire v$EQ1_15290_out0;
wire v$EQ1_15322_out0;
wire v$EQ1_15323_out0;
wire v$EQ1_16122_out0;
wire v$EQ1_16123_out0;
wire v$EQ1_16219_out0;
wire v$EQ1_16220_out0;
wire v$EQ1_16270_out0;
wire v$EQ1_16271_out0;
wire v$EQ1_17399_out0;
wire v$EQ1_18594_out0;
wire v$EQ1_18595_out0;
wire v$EQ1_2516_out0;
wire v$EQ1_2517_out0;
wire v$EQ1_2818_out0;
wire v$EQ1_2819_out0;
wire v$EQ1_2953_out0;
wire v$EQ1_2954_out0;
wire v$EQ1_3211_out0;
wire v$EQ1_3212_out0;
wire v$EQ1_4110_out0;
wire v$EQ1_4111_out0;
wire v$EQ1_5072_out0;
wire v$EQ1_5073_out0;
wire v$EQ1_5080_out0;
wire v$EQ1_5081_out0;
wire v$EQ1_6932_out0;
wire v$EQ1_6933_out0;
wire v$EQ1_7437_out0;
wire v$EQ1_7438_out0;
wire v$EQ1_7789_out0;
wire v$EQ20_9946_out0;
wire v$EQ20_9947_out0;
wire v$EQ20_9948_out0;
wire v$EQ20_9949_out0;
wire v$EQ21_3324_out0;
wire v$EQ21_3325_out0;
wire v$EQ21_3326_out0;
wire v$EQ21_3327_out0;
wire v$EQ22_2836_out0;
wire v$EQ22_2837_out0;
wire v$EQ22_2838_out0;
wire v$EQ22_2839_out0;
wire v$EQ23_3194_out0;
wire v$EQ23_3195_out0;
wire v$EQ23_3196_out0;
wire v$EQ23_3197_out0;
wire v$EQ24_2536_out0;
wire v$EQ24_2537_out0;
wire v$EQ24_2538_out0;
wire v$EQ24_2539_out0;
wire v$EQ2_10797_out0;
wire v$EQ2_10798_out0;
wire v$EQ2_11605_out0;
wire v$EQ2_11606_out0;
wire v$EQ2_12874_out0;
wire v$EQ2_12875_out0;
wire v$EQ2_13623_out0;
wire v$EQ2_13624_out0;
wire v$EQ2_14208_out0;
wire v$EQ2_14209_out0;
wire v$EQ2_14210_out0;
wire v$EQ2_14211_out0;
wire v$EQ2_14300_out0;
wire v$EQ2_14301_out0;
wire v$EQ2_15802_out0;
wire v$EQ2_15803_out0;
wire v$EQ2_16156_out0;
wire v$EQ2_16157_out0;
wire v$EQ2_16393_out0;
wire v$EQ2_16394_out0;
wire v$EQ2_16902_out0;
wire v$EQ2_16903_out0;
wire v$EQ2_18657_out0;
wire v$EQ2_18658_out0;
wire v$EQ2_3209_out0;
wire v$EQ2_3210_out0;
wire v$EQ2_4229_out0;
wire v$EQ2_4230_out0;
wire v$EQ2_7952_out0;
wire v$EQ2_7953_out0;
wire v$EQ3_11712_out0;
wire v$EQ3_11713_out0;
wire v$EQ3_12136_out0;
wire v$EQ3_12137_out0;
wire v$EQ3_13793_out0;
wire v$EQ3_13794_out0;
wire v$EQ3_14302_out0;
wire v$EQ3_14303_out0;
wire v$EQ3_15281_out0;
wire v$EQ3_15282_out0;
wire v$EQ3_15504_out0;
wire v$EQ3_15505_out0;
wire v$EQ3_16544_out0;
wire v$EQ3_16545_out0;
wire v$EQ3_17921_out0;
wire v$EQ3_17922_out0;
wire v$EQ3_1816_out0;
wire v$EQ3_1817_out0;
wire v$EQ3_1818_out0;
wire v$EQ3_1819_out0;
wire v$EQ3_2613_out0;
wire v$EQ3_2614_out0;
wire v$EQ3_4203_out0;
wire v$EQ3_4204_out0;
wire v$EQ3_5436_out0;
wire v$EQ3_5437_out0;
wire v$EQ3_5731_out0;
wire v$EQ3_5732_out0;
wire v$EQ3_7234_out0;
wire v$EQ3_7235_out0;
wire v$EQ3_7898_out0;
wire v$EQ3_7899_out0;
wire v$EQ4_12725_out0;
wire v$EQ4_12726_out0;
wire v$EQ4_16505_out0;
wire v$EQ4_16506_out0;
wire v$EQ4_16578_out0;
wire v$EQ4_16579_out0;
wire v$EQ4_16701_out0;
wire v$EQ4_16702_out0;
wire v$EQ4_18599_out0;
wire v$EQ4_18600_out0;
wire v$EQ4_18601_out0;
wire v$EQ4_18602_out0;
wire v$EQ4_2617_out0;
wire v$EQ4_2618_out0;
wire v$EQ4_3006_out0;
wire v$EQ4_3007_out0;
wire v$EQ4_5414_out0;
wire v$EQ4_5415_out0;
wire v$EQ4_9358_out0;
wire v$EQ4_9359_out0;
wire v$EQ4_9625_out0;
wire v$EQ4_9626_out0;
wire v$EQ5_10028_out0;
wire v$EQ5_10029_out0;
wire v$EQ5_14374_out0;
wire v$EQ5_14375_out0;
wire v$EQ5_1503_out0;
wire v$EQ5_1504_out0;
wire v$EQ5_1911_out0;
wire v$EQ5_1912_out0;
wire v$EQ5_2968_out0;
wire v$EQ5_2969_out0;
wire v$EQ5_3315_out0;
wire v$EQ5_3316_out0;
wire v$EQ5_3317_out0;
wire v$EQ5_3318_out0;
wire v$EQ5_3551_out0;
wire v$EQ5_3552_out0;
wire v$EQ5_4856_out0;
wire v$EQ5_4857_out0;
wire v$EQ5_9106_out0;
wire v$EQ5_9107_out0;
wire v$EQ6_1566_out0;
wire v$EQ6_1567_out0;
wire v$EQ6_15876_out0;
wire v$EQ6_15877_out0;
wire v$EQ6_16172_out0;
wire v$EQ6_16250_out0;
wire v$EQ6_16251_out0;
wire v$EQ6_3957_out0;
wire v$EQ6_3958_out0;
wire v$EQ6_5425_out0;
wire v$EQ6_5426_out0;
wire v$EQ6_5427_out0;
wire v$EQ6_5428_out0;
wire v$EQ6_6411_out0;
wire v$EQ6_6412_out0;
wire v$EQ7_13602_out0;
wire v$EQ7_16898_out0;
wire v$EQ7_16899_out0;
wire v$EQ7_18631_out0;
wire v$EQ7_18632_out0;
wire v$EQ7_231_out0;
wire v$EQ7_232_out0;
wire v$EQ7_3506_out0;
wire v$EQ7_3507_out0;
wire v$EQ7_4085_out0;
wire v$EQ7_4086_out0;
wire v$EQ7_4087_out0;
wire v$EQ7_4088_out0;
wire v$EQ8_14328_out0;
wire v$EQ8_14329_out0;
wire v$EQ8_14414_out0;
wire v$EQ8_14415_out0;
wire v$EQ8_14416_out0;
wire v$EQ8_14417_out0;
wire v$EQ8_16018_out0;
wire v$EQ8_252_out0;
wire v$EQ8_253_out0;
wire v$EQ9_13775_out0;
wire v$EQ9_13776_out0;
wire v$EQ9_13777_out0;
wire v$EQ9_13778_out0;
wire v$EQ9_17768_out0;
wire v$EQ9_17769_out0;
wire v$EQ9_18283_out0;
wire v$EQ9_18284_out0;
wire v$EQ9_7979_out0;
wire v$EQ9_7980_out0;
wire v$EQUAL_11623_out0;
wire v$EQUAL_11624_out0;
wire v$EQUAL_15828_out0;
wire v$EQUAL_15829_out0;
wire v$EQ_13422_out0;
wire v$EQ_13423_out0;
wire v$EQ_14576_out0;
wire v$EQ_14577_out0;
wire v$EQ_3478_out0;
wire v$EQ_3479_out0;
wire v$EQ_3708_out0;
wire v$EQ_3709_out0;
wire v$EQ_431_out0;
wire v$EQ_4328_out0;
wire v$EQ_4329_out0;
wire v$EQ_432_out0;
wire v$EQ_6151_out0;
wire v$EQ_6152_out0;
wire v$ERR_12774_out0;
wire v$ERR_12775_out0;
wire v$EVENPARITY_13588_out0;
wire v$EVENPARITY_13589_out0;
wire v$EXEC1$FPU_13675_out0;
wire v$EXEC1$FPU_13676_out0;
wire v$EXEC1$VIEW$MULTIPLIER_16419_out0;
wire v$EXEC1_10256_out0;
wire v$EXEC1_10257_out0;
wire v$EXEC1_18224_out0;
wire v$EXEC1_18513_out0;
wire v$EXEC1_18719_out0;
wire v$EXEC1_3855_out0;
wire v$EXEC1_7960_out0;
wire v$EXEC1_7961_out0;
wire v$EXEC1_7962_out0;
wire v$EXEC1_7963_out0;
wire v$EXEC1_7964_out0;
wire v$EXEC1_7965_out0;
wire v$EXEC1_7966_out0;
wire v$EXEC1_7967_out0;
wire v$EXEC1_7968_out0;
wire v$EXEC1_7969_out0;
wire v$EXEC1_7970_out0;
wire v$EXEC2_1167_out0;
wire v$EXEC2_1168_out0;
wire v$EXEC2_1469_out0;
wire v$EXEC2_1470_out0;
wire v$EXEC2_15883_out0;
wire v$EXEC2_15884_out0;
wire v$EXEC2_16363_out0;
wire v$EXEC2_16364_out0;
wire v$EXEC2_17638_out0;
wire v$EXEC2_17639_out0;
wire v$EXEC2_1945_out0;
wire v$EXEC2_1946_out0;
wire v$EXEC2_3998_out0;
wire v$EXEC2_3999_out0;
wire v$EXEC2_429_out0;
wire v$EXEC2_430_out0;
wire v$EXEC2_4387_out0;
wire v$EXEC2_4388_out0;
wire v$EXEC2_8015_out0;
wire v$EXEC2_8016_out0;
wire v$EXEC2_8048_out0;
wire v$EXEC2_8049_out0;
wire v$EXEC2_9439_out0;
wire v$EXEC2_9440_out0;
wire v$EXEC2_9863_out0;
wire v$EXEC2_9864_out0;
wire v$EXP$SAME_16546_out0;
wire v$EXP$SAME_16547_out0;
wire v$EXP$SAME_3134_out0;
wire v$EXP$SAME_3135_out0;
wire v$EXP$SAME_903_out0;
wire v$EXP$SAME_904_out0;
wire v$EXTHALT_17883_out0;
wire v$EXTHALT_17884_out0;
wire v$EXTHALT_6459_out0;
wire v$EXTHALT_6460_out0;
wire v$E_17351_out0;
wire v$E_17352_out0;
wire v$Error_3767_out0;
wire v$Error_3768_out0;
wire v$F0_15834_out0;
wire v$F0_15835_out0;
wire v$F1_3488_out0;
wire v$F1_3489_out0;
wire v$F2_12096_out0;
wire v$F2_12097_out0;
wire v$F3_8247_out0;
wire v$F3_8248_out0;
wire v$FINISHED_10861_out0;
wire v$FINISHED_11641_out0;
wire v$FINISHED_13867_out0;
wire v$FINISHED_18669_out0;
wire v$FINISHED_2255_out0;
wire v$FINISHED_7003_out0;
wire v$FINISHED_8010_out0;
wire v$FMUL$FINISHED$VIEWER_3162_out0;
wire v$FMUL$FINISHED_14472_out0;
wire v$FMUL$FINISHED_200_out0;
wire v$FPU$32$BIT$DATAPATH_17727_out0;
wire v$FPU$32$BIT$MUL$PIPELINED_3512_out0;
wire v$FPU$A$EN_11671_out0;
wire v$FPU$LOAD$B_11741_out0;
wire v$FPU$LOAD$B_11742_out0;
wire v$FPU$LOAD$STORE_10979_out0;
wire v$FPU$LOAD$STORE_10980_out0;
wire v$F_1969_out0;
wire v$F_1970_out0;
wire v$G$AB_9136_out0;
wire v$G$AB_9137_out0;
wire v$G$AB_9138_out0;
wire v$G$AB_9139_out0;
wire v$G$AB_9140_out0;
wire v$G$AB_9141_out0;
wire v$G$AB_9142_out0;
wire v$G$AB_9143_out0;
wire v$G$AB_9144_out0;
wire v$G$AB_9145_out0;
wire v$G$AB_9146_out0;
wire v$G$AB_9147_out0;
wire v$G$AB_9148_out0;
wire v$G$AB_9149_out0;
wire v$G$AB_9150_out0;
wire v$G$AB_9151_out0;
wire v$G$AB_9152_out0;
wire v$G$AB_9153_out0;
wire v$G$AB_9154_out0;
wire v$G$AB_9155_out0;
wire v$G$AB_9156_out0;
wire v$G$AB_9157_out0;
wire v$G$AB_9158_out0;
wire v$G$AB_9159_out0;
wire v$G$AB_9160_out0;
wire v$G$AB_9161_out0;
wire v$G$AB_9162_out0;
wire v$G$AB_9163_out0;
wire v$G$AB_9164_out0;
wire v$G$AB_9165_out0;
wire v$G$AB_9166_out0;
wire v$G$AB_9167_out0;
wire v$G$AB_9168_out0;
wire v$G$AB_9169_out0;
wire v$G$AB_9170_out0;
wire v$G$AB_9171_out0;
wire v$G$AB_9172_out0;
wire v$G$AB_9173_out0;
wire v$G$AB_9174_out0;
wire v$G$AB_9175_out0;
wire v$G$AB_9176_out0;
wire v$G$AB_9177_out0;
wire v$G$AB_9178_out0;
wire v$G$AB_9179_out0;
wire v$G$AB_9180_out0;
wire v$G$AB_9181_out0;
wire v$G$AB_9182_out0;
wire v$G$AB_9183_out0;
wire v$G$AB_9184_out0;
wire v$G$AB_9185_out0;
wire v$G$AB_9186_out0;
wire v$G$AB_9187_out0;
wire v$G$AB_9188_out0;
wire v$G$AB_9189_out0;
wire v$G$AB_9190_out0;
wire v$G$AB_9191_out0;
wire v$G$AB_9192_out0;
wire v$G$AB_9193_out0;
wire v$G$AB_9194_out0;
wire v$G$AB_9195_out0;
wire v$G$AB_9196_out0;
wire v$G$AB_9197_out0;
wire v$G$AB_9198_out0;
wire v$G$AB_9199_out0;
wire v$G$AB_9200_out0;
wire v$G$AB_9201_out0;
wire v$G$AB_9202_out0;
wire v$G$AB_9203_out0;
wire v$G$AB_9204_out0;
wire v$G$AB_9205_out0;
wire v$G$AB_9206_out0;
wire v$G$AB_9207_out0;
wire v$G$AB_9208_out0;
wire v$G$AB_9209_out0;
wire v$G$AB_9210_out0;
wire v$G$AB_9211_out0;
wire v$G$AB_9212_out0;
wire v$G$AB_9213_out0;
wire v$G$AB_9214_out0;
wire v$G$AB_9215_out0;
wire v$G$AB_9216_out0;
wire v$G$AB_9217_out0;
wire v$G$AB_9218_out0;
wire v$G$AB_9219_out0;
wire v$G$AB_9220_out0;
wire v$G$AB_9221_out0;
wire v$G$AB_9222_out0;
wire v$G$AB_9223_out0;
wire v$G$AB_9224_out0;
wire v$G$AB_9225_out0;
wire v$G$AB_9226_out0;
wire v$G$AB_9227_out0;
wire v$G$AB_9228_out0;
wire v$G$AB_9229_out0;
wire v$G$AB_9230_out0;
wire v$G$AB_9231_out0;
wire v$G$AB_9232_out0;
wire v$G$AB_9233_out0;
wire v$G$AB_9234_out0;
wire v$G$AB_9235_out0;
wire v$G$AB_9236_out0;
wire v$G$AB_9237_out0;
wire v$G$AB_9238_out0;
wire v$G$AB_9239_out0;
wire v$G$AB_9240_out0;
wire v$G$AB_9241_out0;
wire v$G$AB_9242_out0;
wire v$G$AB_9243_out0;
wire v$G$AB_9244_out0;
wire v$G$AB_9245_out0;
wire v$G$AB_9246_out0;
wire v$G$AB_9247_out0;
wire v$G$AB_9248_out0;
wire v$G$AB_9249_out0;
wire v$G$AB_9250_out0;
wire v$G$AB_9251_out0;
wire v$G$AB_9252_out0;
wire v$G$AB_9253_out0;
wire v$G$AB_9254_out0;
wire v$G$AB_9255_out0;
wire v$G$AB_9256_out0;
wire v$G$AB_9257_out0;
wire v$G$AB_9258_out0;
wire v$G$AB_9259_out0;
wire v$G$AB_9260_out0;
wire v$G$AB_9261_out0;
wire v$G$AB_9262_out0;
wire v$G$AB_9263_out0;
wire v$G$AB_9264_out0;
wire v$G$AB_9265_out0;
wire v$G$AB_9266_out0;
wire v$G$AB_9267_out0;
wire v$G$AB_9268_out0;
wire v$G$AB_9269_out0;
wire v$G$AB_9270_out0;
wire v$G$AB_9271_out0;
wire v$G$AB_9272_out0;
wire v$G$AB_9273_out0;
wire v$G$AB_9274_out0;
wire v$G$AB_9275_out0;
wire v$G$AB_9276_out0;
wire v$G$AB_9277_out0;
wire v$G$AB_9278_out0;
wire v$G$AB_9279_out0;
wire v$G$AB_9280_out0;
wire v$G$AB_9281_out0;
wire v$G$AB_9282_out0;
wire v$G$AB_9283_out0;
wire v$G$AB_9284_out0;
wire v$G$AB_9285_out0;
wire v$G$AB_9286_out0;
wire v$G$AB_9287_out0;
wire v$G$AB_9288_out0;
wire v$G$AB_9289_out0;
wire v$G$AB_9290_out0;
wire v$G$AB_9291_out0;
wire v$G$AB_9292_out0;
wire v$G$AB_9293_out0;
wire v$G$AB_9294_out0;
wire v$G$AB_9295_out0;
wire v$G$AB_9296_out0;
wire v$G$AB_9297_out0;
wire v$G$AB_9298_out0;
wire v$G$AB_9299_out0;
wire v$G$AB_9300_out0;
wire v$G$AB_9301_out0;
wire v$G$AB_9302_out0;
wire v$G$AB_9303_out0;
wire v$G$AB_9304_out0;
wire v$G$AB_9305_out0;
wire v$G$AB_9306_out0;
wire v$G$AB_9307_out0;
wire v$G$AB_9308_out0;
wire v$G$AB_9309_out0;
wire v$G$AB_9310_out0;
wire v$G$AB_9311_out0;
wire v$G$AB_9312_out0;
wire v$G$AB_9313_out0;
wire v$G$AB_9314_out0;
wire v$G$AB_9315_out0;
wire v$G$AB_9316_out0;
wire v$G$AB_9317_out0;
wire v$G$AB_9318_out0;
wire v$G$AB_9319_out0;
wire v$G$AB_9320_out0;
wire v$G$AB_9321_out0;
wire v$G$AB_9322_out0;
wire v$G$AB_9323_out0;
wire v$G$AB_9324_out0;
wire v$G$AB_9325_out0;
wire v$G$AB_9326_out0;
wire v$G$AB_9327_out0;
wire v$G$AB_9328_out0;
wire v$G$AB_9329_out0;
wire v$G$AB_9330_out0;
wire v$G$AB_9331_out0;
wire v$G$AB_9332_out0;
wire v$G$AB_9333_out0;
wire v$G$AB_9334_out0;
wire v$G$AB_9335_out0;
wire v$G$AB_9336_out0;
wire v$G$AB_9337_out0;
wire v$G$AB_9338_out0;
wire v$G$AB_9339_out0;
wire v$G$AB_9340_out0;
wire v$G$AD_17086_out0;
wire v$G$AD_17087_out0;
wire v$G$AD_17088_out0;
wire v$G$AD_17089_out0;
wire v$G$AD_17090_out0;
wire v$G$AD_17091_out0;
wire v$G$AD_17092_out0;
wire v$G$AD_17093_out0;
wire v$G$AD_17094_out0;
wire v$G$AD_17095_out0;
wire v$G$AD_17096_out0;
wire v$G$AD_17097_out0;
wire v$G$AD_17098_out0;
wire v$G$AD_17099_out0;
wire v$G$AD_17100_out0;
wire v$G$AD_17101_out0;
wire v$G$AD_17102_out0;
wire v$G$AD_17103_out0;
wire v$G$AD_17104_out0;
wire v$G$AD_17105_out0;
wire v$G$AD_17106_out0;
wire v$G$AD_17107_out0;
wire v$G$AD_17108_out0;
wire v$G$AD_17109_out0;
wire v$G$AD_17110_out0;
wire v$G$AD_17111_out0;
wire v$G$AD_17112_out0;
wire v$G$AD_17113_out0;
wire v$G$AD_17114_out0;
wire v$G$AD_17115_out0;
wire v$G$AD_17116_out0;
wire v$G$AD_17117_out0;
wire v$G$AD_17118_out0;
wire v$G$AD_17119_out0;
wire v$G$AD_17120_out0;
wire v$G$AD_17121_out0;
wire v$G$AD_17122_out0;
wire v$G$AD_17123_out0;
wire v$G$AD_17124_out0;
wire v$G$AD_17125_out0;
wire v$G$AD_17126_out0;
wire v$G$AD_17127_out0;
wire v$G$AD_17128_out0;
wire v$G$AD_17129_out0;
wire v$G$AD_17130_out0;
wire v$G$AD_17131_out0;
wire v$G$AD_17132_out0;
wire v$G$AD_17133_out0;
wire v$G$AD_17134_out0;
wire v$G$AD_17135_out0;
wire v$G$AD_17136_out0;
wire v$G$AD_17137_out0;
wire v$G$AD_17138_out0;
wire v$G$AD_17139_out0;
wire v$G$AD_17140_out0;
wire v$G$AD_17141_out0;
wire v$G$AD_17142_out0;
wire v$G$AD_17143_out0;
wire v$G$AD_17144_out0;
wire v$G$AD_17145_out0;
wire v$G$AD_17146_out0;
wire v$G$AD_17147_out0;
wire v$G$AD_17148_out0;
wire v$G$AD_17149_out0;
wire v$G$AD_17150_out0;
wire v$G$AD_17151_out0;
wire v$G$AD_17152_out0;
wire v$G$AD_17153_out0;
wire v$G$AD_17154_out0;
wire v$G$AD_17155_out0;
wire v$G$AD_17156_out0;
wire v$G$AD_17157_out0;
wire v$G$AD_17158_out0;
wire v$G$AD_17159_out0;
wire v$G$AD_17160_out0;
wire v$G$AD_17161_out0;
wire v$G$AD_17162_out0;
wire v$G$AD_17163_out0;
wire v$G$AD_17164_out0;
wire v$G$AD_17165_out0;
wire v$G$AD_17166_out0;
wire v$G$AD_17167_out0;
wire v$G$AD_17168_out0;
wire v$G$AD_17169_out0;
wire v$G$AD_17170_out0;
wire v$G$AD_17171_out0;
wire v$G$AD_17172_out0;
wire v$G$AD_17173_out0;
wire v$G$AD_17174_out0;
wire v$G$AD_17175_out0;
wire v$G$AD_17176_out0;
wire v$G$AD_17177_out0;
wire v$G$AD_17178_out0;
wire v$G$AD_17179_out0;
wire v$G$AD_17180_out0;
wire v$G$AD_17181_out0;
wire v$G$AD_17182_out0;
wire v$G$AD_17183_out0;
wire v$G$AD_17184_out0;
wire v$G$AD_17185_out0;
wire v$G$AD_17186_out0;
wire v$G$AD_17187_out0;
wire v$G$AD_17188_out0;
wire v$G$AD_17189_out0;
wire v$G$AD_17190_out0;
wire v$G$AD_17191_out0;
wire v$G$AD_17192_out0;
wire v$G$AD_17193_out0;
wire v$G$AD_17194_out0;
wire v$G$AD_17195_out0;
wire v$G$AD_17196_out0;
wire v$G$AD_17197_out0;
wire v$G$AD_17198_out0;
wire v$G$AD_17199_out0;
wire v$G$AD_17200_out0;
wire v$G$AD_17201_out0;
wire v$G$AD_17202_out0;
wire v$G$AD_17203_out0;
wire v$G$AD_17204_out0;
wire v$G$AD_17205_out0;
wire v$G$AD_17206_out0;
wire v$G$AD_17207_out0;
wire v$G$AD_17208_out0;
wire v$G$AD_17209_out0;
wire v$G$AD_17210_out0;
wire v$G$AD_17211_out0;
wire v$G$AD_17212_out0;
wire v$G$AD_17213_out0;
wire v$G$AD_17214_out0;
wire v$G$AD_17215_out0;
wire v$G$AD_17216_out0;
wire v$G$AD_17217_out0;
wire v$G$AD_17218_out0;
wire v$G$AD_17219_out0;
wire v$G$AD_17220_out0;
wire v$G$AD_17221_out0;
wire v$G$AD_17222_out0;
wire v$G$AD_17223_out0;
wire v$G$AD_17224_out0;
wire v$G$AD_17225_out0;
wire v$G$AD_17226_out0;
wire v$G$AD_17227_out0;
wire v$G$AD_17228_out0;
wire v$G$AD_17229_out0;
wire v$G$AD_17230_out0;
wire v$G$AD_17231_out0;
wire v$G$AD_17232_out0;
wire v$G$AD_17233_out0;
wire v$G$AD_17234_out0;
wire v$G$AD_17235_out0;
wire v$G$AD_17236_out0;
wire v$G$AD_17237_out0;
wire v$G$AD_17238_out0;
wire v$G$AD_17239_out0;
wire v$G$AD_17240_out0;
wire v$G$AD_17241_out0;
wire v$G$AD_17242_out0;
wire v$G$AD_17243_out0;
wire v$G$AD_17244_out0;
wire v$G$AD_17245_out0;
wire v$G$AD_17246_out0;
wire v$G$AD_17247_out0;
wire v$G$AD_17248_out0;
wire v$G$AD_17249_out0;
wire v$G$AD_17250_out0;
wire v$G$AD_17251_out0;
wire v$G$AD_17252_out0;
wire v$G$AD_17253_out0;
wire v$G$AD_17254_out0;
wire v$G$AD_17255_out0;
wire v$G$AD_17256_out0;
wire v$G$AD_17257_out0;
wire v$G$AD_17258_out0;
wire v$G$AD_17259_out0;
wire v$G$AD_17260_out0;
wire v$G$AD_17261_out0;
wire v$G$AD_17262_out0;
wire v$G$AD_17263_out0;
wire v$G$AD_17264_out0;
wire v$G$AD_17265_out0;
wire v$G$AD_17266_out0;
wire v$G$AD_17267_out0;
wire v$G$AD_17268_out0;
wire v$G$AD_17269_out0;
wire v$G$AD_17270_out0;
wire v$G$AD_17271_out0;
wire v$G$AD_17272_out0;
wire v$G$AD_17273_out0;
wire v$G$AD_17274_out0;
wire v$G$AD_17275_out0;
wire v$G$AD_17276_out0;
wire v$G$AD_17277_out0;
wire v$G$AD_17278_out0;
wire v$G$AD_17279_out0;
wire v$G$AD_17280_out0;
wire v$G$AD_17281_out0;
wire v$G$AD_17282_out0;
wire v$G$AD_17283_out0;
wire v$G$AD_17284_out0;
wire v$G$AD_17285_out0;
wire v$G$AD_17286_out0;
wire v$G$AD_17287_out0;
wire v$G$AD_17288_out0;
wire v$G$AD_17289_out0;
wire v$G$AD_17290_out0;
wire v$G$CD_1000_out0;
wire v$G$CD_1001_out0;
wire v$G$CD_1002_out0;
wire v$G$CD_1003_out0;
wire v$G$CD_1004_out0;
wire v$G$CD_1005_out0;
wire v$G$CD_1006_out0;
wire v$G$CD_1007_out0;
wire v$G$CD_1008_out0;
wire v$G$CD_1009_out0;
wire v$G$CD_1010_out0;
wire v$G$CD_1011_out0;
wire v$G$CD_1012_out0;
wire v$G$CD_1013_out0;
wire v$G$CD_1014_out0;
wire v$G$CD_1015_out0;
wire v$G$CD_1016_out0;
wire v$G$CD_1017_out0;
wire v$G$CD_1018_out0;
wire v$G$CD_1019_out0;
wire v$G$CD_1020_out0;
wire v$G$CD_1021_out0;
wire v$G$CD_1022_out0;
wire v$G$CD_1023_out0;
wire v$G$CD_1024_out0;
wire v$G$CD_1025_out0;
wire v$G$CD_1026_out0;
wire v$G$CD_1027_out0;
wire v$G$CD_1028_out0;
wire v$G$CD_1029_out0;
wire v$G$CD_1030_out0;
wire v$G$CD_1031_out0;
wire v$G$CD_1032_out0;
wire v$G$CD_1033_out0;
wire v$G$CD_1034_out0;
wire v$G$CD_1035_out0;
wire v$G$CD_1036_out0;
wire v$G$CD_1037_out0;
wire v$G$CD_1038_out0;
wire v$G$CD_1039_out0;
wire v$G$CD_1040_out0;
wire v$G$CD_1041_out0;
wire v$G$CD_1042_out0;
wire v$G$CD_1043_out0;
wire v$G$CD_1044_out0;
wire v$G$CD_1045_out0;
wire v$G$CD_1046_out0;
wire v$G$CD_1047_out0;
wire v$G$CD_1048_out0;
wire v$G$CD_1049_out0;
wire v$G$CD_1050_out0;
wire v$G$CD_1051_out0;
wire v$G$CD_1052_out0;
wire v$G$CD_1053_out0;
wire v$G$CD_1054_out0;
wire v$G$CD_1055_out0;
wire v$G$CD_1056_out0;
wire v$G$CD_1057_out0;
wire v$G$CD_1058_out0;
wire v$G$CD_1059_out0;
wire v$G$CD_1060_out0;
wire v$G$CD_1061_out0;
wire v$G$CD_1062_out0;
wire v$G$CD_1063_out0;
wire v$G$CD_1064_out0;
wire v$G$CD_1065_out0;
wire v$G$CD_1066_out0;
wire v$G$CD_1067_out0;
wire v$G$CD_1068_out0;
wire v$G$CD_1069_out0;
wire v$G$CD_1070_out0;
wire v$G$CD_1071_out0;
wire v$G$CD_1072_out0;
wire v$G$CD_1073_out0;
wire v$G$CD_1074_out0;
wire v$G$CD_1075_out0;
wire v$G$CD_1076_out0;
wire v$G$CD_1077_out0;
wire v$G$CD_1078_out0;
wire v$G$CD_1079_out0;
wire v$G$CD_1080_out0;
wire v$G$CD_1081_out0;
wire v$G$CD_1082_out0;
wire v$G$CD_1083_out0;
wire v$G$CD_1084_out0;
wire v$G$CD_1085_out0;
wire v$G$CD_1086_out0;
wire v$G$CD_1087_out0;
wire v$G$CD_1088_out0;
wire v$G$CD_1089_out0;
wire v$G$CD_1090_out0;
wire v$G$CD_1091_out0;
wire v$G$CD_1092_out0;
wire v$G$CD_1093_out0;
wire v$G$CD_1094_out0;
wire v$G$CD_1095_out0;
wire v$G$CD_1096_out0;
wire v$G$CD_1097_out0;
wire v$G$CD_1098_out0;
wire v$G$CD_1099_out0;
wire v$G$CD_1100_out0;
wire v$G$CD_1101_out0;
wire v$G$CD_1102_out0;
wire v$G$CD_1103_out0;
wire v$G$CD_1104_out0;
wire v$G$CD_1105_out0;
wire v$G$CD_1106_out0;
wire v$G$CD_1107_out0;
wire v$G$CD_1108_out0;
wire v$G$CD_1109_out0;
wire v$G$CD_1110_out0;
wire v$G$CD_1111_out0;
wire v$G$CD_1112_out0;
wire v$G$CD_1113_out0;
wire v$G$CD_1114_out0;
wire v$G$CD_1115_out0;
wire v$G$CD_1116_out0;
wire v$G$CD_1117_out0;
wire v$G$CD_1118_out0;
wire v$G$CD_914_out0;
wire v$G$CD_915_out0;
wire v$G$CD_916_out0;
wire v$G$CD_917_out0;
wire v$G$CD_918_out0;
wire v$G$CD_919_out0;
wire v$G$CD_920_out0;
wire v$G$CD_921_out0;
wire v$G$CD_922_out0;
wire v$G$CD_923_out0;
wire v$G$CD_924_out0;
wire v$G$CD_925_out0;
wire v$G$CD_926_out0;
wire v$G$CD_927_out0;
wire v$G$CD_928_out0;
wire v$G$CD_929_out0;
wire v$G$CD_930_out0;
wire v$G$CD_931_out0;
wire v$G$CD_932_out0;
wire v$G$CD_933_out0;
wire v$G$CD_934_out0;
wire v$G$CD_935_out0;
wire v$G$CD_936_out0;
wire v$G$CD_937_out0;
wire v$G$CD_938_out0;
wire v$G$CD_939_out0;
wire v$G$CD_940_out0;
wire v$G$CD_941_out0;
wire v$G$CD_942_out0;
wire v$G$CD_943_out0;
wire v$G$CD_944_out0;
wire v$G$CD_945_out0;
wire v$G$CD_946_out0;
wire v$G$CD_947_out0;
wire v$G$CD_948_out0;
wire v$G$CD_949_out0;
wire v$G$CD_950_out0;
wire v$G$CD_951_out0;
wire v$G$CD_952_out0;
wire v$G$CD_953_out0;
wire v$G$CD_954_out0;
wire v$G$CD_955_out0;
wire v$G$CD_956_out0;
wire v$G$CD_957_out0;
wire v$G$CD_958_out0;
wire v$G$CD_959_out0;
wire v$G$CD_960_out0;
wire v$G$CD_961_out0;
wire v$G$CD_962_out0;
wire v$G$CD_963_out0;
wire v$G$CD_964_out0;
wire v$G$CD_965_out0;
wire v$G$CD_966_out0;
wire v$G$CD_967_out0;
wire v$G$CD_968_out0;
wire v$G$CD_969_out0;
wire v$G$CD_970_out0;
wire v$G$CD_971_out0;
wire v$G$CD_972_out0;
wire v$G$CD_973_out0;
wire v$G$CD_974_out0;
wire v$G$CD_975_out0;
wire v$G$CD_976_out0;
wire v$G$CD_977_out0;
wire v$G$CD_978_out0;
wire v$G$CD_979_out0;
wire v$G$CD_980_out0;
wire v$G$CD_981_out0;
wire v$G$CD_982_out0;
wire v$G$CD_983_out0;
wire v$G$CD_984_out0;
wire v$G$CD_985_out0;
wire v$G$CD_986_out0;
wire v$G$CD_987_out0;
wire v$G$CD_988_out0;
wire v$G$CD_989_out0;
wire v$G$CD_990_out0;
wire v$G$CD_991_out0;
wire v$G$CD_992_out0;
wire v$G$CD_993_out0;
wire v$G$CD_994_out0;
wire v$G$CD_995_out0;
wire v$G$CD_996_out0;
wire v$G$CD_997_out0;
wire v$G$CD_998_out0;
wire v$G$CD_999_out0;
wire v$G0_15942_out0;
wire v$G0_15943_out0;
wire v$G0_15944_out0;
wire v$G0_15945_out0;
wire v$G0_15946_out0;
wire v$G10_10271_out0;
wire v$G10_10272_out0;
wire v$G10_1182_out0;
wire v$G10_1183_out0;
wire v$G10_13314_out0;
wire v$G10_13315_out0;
wire v$G10_1380_out0;
wire v$G10_1381_out0;
wire v$G10_1382_out0;
wire v$G10_1383_out0;
wire v$G10_1384_out0;
wire v$G10_1385_out0;
wire v$G10_1386_out0;
wire v$G10_1387_out0;
wire v$G10_1388_out0;
wire v$G10_1389_out0;
wire v$G10_1390_out0;
wire v$G10_1391_out0;
wire v$G10_1392_out0;
wire v$G10_1393_out0;
wire v$G10_1394_out0;
wire v$G10_1395_out0;
wire v$G10_1396_out0;
wire v$G10_1397_out0;
wire v$G10_1398_out0;
wire v$G10_1399_out0;
wire v$G10_1400_out0;
wire v$G10_1401_out0;
wire v$G10_1402_out0;
wire v$G10_1403_out0;
wire v$G10_1404_out0;
wire v$G10_1405_out0;
wire v$G10_1406_out0;
wire v$G10_1407_out0;
wire v$G10_1408_out0;
wire v$G10_1409_out0;
wire v$G10_1410_out0;
wire v$G10_1411_out0;
wire v$G10_1412_out0;
wire v$G10_1413_out0;
wire v$G10_1414_out0;
wire v$G10_1415_out0;
wire v$G10_1416_out0;
wire v$G10_1417_out0;
wire v$G10_1418_out0;
wire v$G10_1419_out0;
wire v$G10_1420_out0;
wire v$G10_1421_out0;
wire v$G10_1422_out0;
wire v$G10_1423_out0;
wire v$G10_1424_out0;
wire v$G10_1425_out0;
wire v$G10_1426_out0;
wire v$G10_1427_out0;
wire v$G10_14566_out0;
wire v$G10_14567_out0;
wire v$G10_14588_out0;
wire v$G10_14589_out0;
wire v$G10_14893_out0;
wire v$G10_14894_out0;
wire v$G10_16091_out0;
wire v$G10_16092_out0;
wire v$G10_16500_out0;
wire v$G10_16501_out0;
wire v$G10_18186_out0;
wire v$G10_18187_out0;
wire v$G10_1833_out0;
wire v$G10_1834_out0;
wire v$G10_1835_out0;
wire v$G10_1836_out0;
wire v$G10_1837_out0;
wire v$G10_18485_out0;
wire v$G10_18486_out0;
wire v$G10_1998_out0;
wire v$G10_1999_out0;
wire v$G10_2906_out0;
wire v$G10_2907_out0;
wire v$G10_3803_out0;
wire v$G10_3804_out0;
wire v$G10_6689_out0;
wire v$G10_6690_out0;
wire v$G11_11063_out0;
wire v$G11_11064_out0;
wire v$G11_11065_out0;
wire v$G11_11066_out0;
wire v$G11_11067_out0;
wire v$G11_11845_out0;
wire v$G11_11846_out0;
wire v$G11_13406_out0;
wire v$G11_13407_out0;
wire v$G11_14584_out0;
wire v$G11_14585_out0;
wire v$G11_15637_out0;
wire v$G11_15638_out0;
wire v$G11_15639_out0;
wire v$G11_15640_out0;
wire v$G11_15641_out0;
wire v$G11_15642_out0;
wire v$G11_15643_out0;
wire v$G11_15644_out0;
wire v$G11_15645_out0;
wire v$G11_15646_out0;
wire v$G11_15647_out0;
wire v$G11_15648_out0;
wire v$G11_15649_out0;
wire v$G11_15650_out0;
wire v$G11_15651_out0;
wire v$G11_15652_out0;
wire v$G11_15653_out0;
wire v$G11_15654_out0;
wire v$G11_15655_out0;
wire v$G11_15656_out0;
wire v$G11_15657_out0;
wire v$G11_15658_out0;
wire v$G11_15659_out0;
wire v$G11_15660_out0;
wire v$G11_1619_out0;
wire v$G11_1620_out0;
wire v$G11_18016_out0;
wire v$G11_18017_out0;
wire v$G11_2287_out0;
wire v$G11_2288_out0;
wire v$G11_2978_out0;
wire v$G11_2979_out0;
wire v$G11_3012_out0;
wire v$G11_3013_out0;
wire v$G11_3251_out0;
wire v$G11_3252_out0;
wire v$G11_4865_out0;
wire v$G11_4866_out0;
wire v$G11_8202_out0;
wire v$G11_8203_out0;
wire v$G11_8230_out0;
wire v$G11_8231_out0;
wire v$G11_8263_out0;
wire v$G11_8264_out0;
wire v$G11_8842_out0;
wire v$G11_8843_out0;
wire v$G11_8844_out0;
wire v$G11_8845_out0;
wire v$G11_8846_out0;
wire v$G11_8847_out0;
wire v$G11_8848_out0;
wire v$G11_8849_out0;
wire v$G11_8850_out0;
wire v$G11_8851_out0;
wire v$G11_8852_out0;
wire v$G11_8853_out0;
wire v$G11_8854_out0;
wire v$G11_8855_out0;
wire v$G11_8856_out0;
wire v$G11_8857_out0;
wire v$G11_8858_out0;
wire v$G11_8859_out0;
wire v$G11_8860_out0;
wire v$G11_8861_out0;
wire v$G11_8862_out0;
wire v$G11_8863_out0;
wire v$G11_8864_out0;
wire v$G11_8865_out0;
wire v$G11_8866_out0;
wire v$G11_8867_out0;
wire v$G11_8868_out0;
wire v$G11_8869_out0;
wire v$G11_8870_out0;
wire v$G11_8871_out0;
wire v$G11_8872_out0;
wire v$G11_8873_out0;
wire v$G11_8874_out0;
wire v$G11_8875_out0;
wire v$G11_8876_out0;
wire v$G11_8877_out0;
wire v$G11_8878_out0;
wire v$G11_8879_out0;
wire v$G11_8880_out0;
wire v$G11_8881_out0;
wire v$G11_8882_out0;
wire v$G11_8883_out0;
wire v$G11_8884_out0;
wire v$G11_8885_out0;
wire v$G11_8886_out0;
wire v$G11_8887_out0;
wire v$G11_8888_out0;
wire v$G11_8889_out0;
wire v$G11_9603_out0;
wire v$G11_9604_out0;
wire v$G12_11896_out0;
wire v$G12_11897_out0;
wire v$G12_11978_out0;
wire v$G12_11979_out0;
wire v$G12_13795_out0;
wire v$G12_13796_out0;
wire v$G12_14705_out0;
wire v$G12_14706_out0;
wire v$G12_16252_out0;
wire v$G12_16253_out0;
wire v$G12_16468_out0;
wire v$G12_16469_out0;
wire v$G12_16470_out0;
wire v$G12_16471_out0;
wire v$G12_16472_out0;
wire v$G12_16473_out0;
wire v$G12_16474_out0;
wire v$G12_16475_out0;
wire v$G12_16476_out0;
wire v$G12_16477_out0;
wire v$G12_16478_out0;
wire v$G12_16479_out0;
wire v$G12_16480_out0;
wire v$G12_16481_out0;
wire v$G12_16482_out0;
wire v$G12_16483_out0;
wire v$G12_16484_out0;
wire v$G12_16485_out0;
wire v$G12_16486_out0;
wire v$G12_16487_out0;
wire v$G12_16488_out0;
wire v$G12_16489_out0;
wire v$G12_16490_out0;
wire v$G12_16491_out0;
wire v$G12_1820_out0;
wire v$G12_1821_out0;
wire v$G12_2215_out0;
wire v$G12_2216_out0;
wire v$G12_3615_out0;
wire v$G12_3616_out0;
wire v$G12_4833_out0;
wire v$G12_4834_out0;
wire v$G12_6167_out0;
wire v$G12_6168_out0;
wire v$G12_7042_out0;
wire v$G12_7043_out0;
wire v$G12_7044_out0;
wire v$G12_7045_out0;
wire v$G12_7046_out0;
wire v$G12_9942_out0;
wire v$G12_9943_out0;
wire v$G13_10230_out0;
wire v$G13_10231_out0;
wire v$G13_12160_out0;
wire v$G13_12161_out0;
wire v$G13_13444_out0;
wire v$G13_13445_out0;
wire v$G13_14852_out0;
wire v$G13_14853_out0;
wire v$G13_15105_out0;
wire v$G13_15106_out0;
wire v$G13_16532_out0;
wire v$G13_16533_out0;
wire v$G13_1689_out0;
wire v$G13_1690_out0;
wire v$G13_198_out0;
wire v$G13_199_out0;
wire v$G13_2828_out0;
wire v$G13_2829_out0;
wire v$G13_2830_out0;
wire v$G13_2831_out0;
wire v$G13_2832_out0;
wire v$G13_4351_out0;
wire v$G13_4352_out0;
wire v$G13_4399_out0;
wire v$G13_4400_out0;
wire v$G13_4401_out0;
wire v$G13_4402_out0;
wire v$G13_4403_out0;
wire v$G13_4404_out0;
wire v$G13_4405_out0;
wire v$G13_4406_out0;
wire v$G13_4407_out0;
wire v$G13_4408_out0;
wire v$G13_4409_out0;
wire v$G13_4410_out0;
wire v$G13_4411_out0;
wire v$G13_4412_out0;
wire v$G13_4413_out0;
wire v$G13_4414_out0;
wire v$G13_4415_out0;
wire v$G13_4416_out0;
wire v$G13_4417_out0;
wire v$G13_4418_out0;
wire v$G13_4419_out0;
wire v$G13_4420_out0;
wire v$G13_4421_out0;
wire v$G13_4422_out0;
wire v$G13_7894_out0;
wire v$G13_7895_out0;
wire v$G14_12046_out0;
wire v$G14_12047_out0;
wire v$G14_12643_out0;
wire v$G14_12644_out0;
wire v$G14_12645_out0;
wire v$G14_12646_out0;
wire v$G14_14681_out0;
wire v$G14_14682_out0;
wire v$G14_15291_out0;
wire v$G14_15292_out0;
wire v$G14_15815_out0;
wire v$G14_15816_out0;
wire v$G14_1673_out0;
wire v$G14_1674_out0;
wire v$G14_17038_out0;
wire v$G14_17039_out0;
wire v$G14_17976_out0;
wire v$G14_17977_out0;
wire v$G14_17978_out0;
wire v$G14_17979_out0;
wire v$G14_17980_out0;
wire v$G14_18435_out0;
wire v$G14_18436_out0;
wire v$G14_5129_out0;
wire v$G14_5130_out0;
wire v$G14_5384_out0;
wire v$G14_5385_out0;
wire v$G14_6127_out0;
wire v$G14_6128_out0;
wire v$G14_6428_out0;
wire v$G14_6429_out0;
wire v$G15_11030_out0;
wire v$G15_11031_out0;
wire v$G15_11032_out0;
wire v$G15_11033_out0;
wire v$G15_11034_out0;
wire v$G15_13391_out0;
wire v$G15_13392_out0;
wire v$G15_13420_out0;
wire v$G15_13421_out0;
wire v$G15_13603_out0;
wire v$G15_13604_out0;
wire v$G15_13643_out0;
wire v$G15_13644_out0;
wire v$G15_13645_out0;
wire v$G15_13646_out0;
wire v$G15_13647_out0;
wire v$G15_13648_out0;
wire v$G15_13649_out0;
wire v$G15_13650_out0;
wire v$G15_13651_out0;
wire v$G15_13652_out0;
wire v$G15_13653_out0;
wire v$G15_13654_out0;
wire v$G15_13655_out0;
wire v$G15_13656_out0;
wire v$G15_13657_out0;
wire v$G15_13658_out0;
wire v$G15_13659_out0;
wire v$G15_13660_out0;
wire v$G15_13661_out0;
wire v$G15_13662_out0;
wire v$G15_13663_out0;
wire v$G15_13664_out0;
wire v$G15_13665_out0;
wire v$G15_13666_out0;
wire v$G15_14582_out0;
wire v$G15_14583_out0;
wire v$G15_17828_out0;
wire v$G15_17829_out0;
wire v$G15_18535_out0;
wire v$G15_18536_out0;
wire v$G15_1868_out0;
wire v$G15_1869_out0;
wire v$G15_2283_out0;
wire v$G15_2677_out0;
wire v$G15_2678_out0;
wire v$G15_4205_out0;
wire v$G15_4206_out0;
wire v$G15_5478_out0;
wire v$G15_5479_out0;
wire v$G16_11965_out0;
wire v$G16_11966_out0;
wire v$G16_1314_out0;
wire v$G16_1315_out0;
wire v$G16_16448_out0;
wire v$G16_16449_out0;
wire v$G16_16450_out0;
wire v$G16_16451_out0;
wire v$G16_16452_out0;
wire v$G16_16862_out0;
wire v$G16_16863_out0;
wire v$G16_16864_out0;
wire v$G16_16865_out0;
wire v$G16_16866_out0;
wire v$G16_16867_out0;
wire v$G16_16868_out0;
wire v$G16_16869_out0;
wire v$G16_16870_out0;
wire v$G16_16871_out0;
wire v$G16_16872_out0;
wire v$G16_16873_out0;
wire v$G16_16874_out0;
wire v$G16_16875_out0;
wire v$G16_16876_out0;
wire v$G16_16877_out0;
wire v$G16_16878_out0;
wire v$G16_16879_out0;
wire v$G16_16880_out0;
wire v$G16_16881_out0;
wire v$G16_16882_out0;
wire v$G16_16883_out0;
wire v$G16_16884_out0;
wire v$G16_16885_out0;
wire v$G16_16978_out0;
wire v$G16_16979_out0;
wire v$G16_16990_out0;
wire v$G16_16991_out0;
wire v$G16_18781_out0;
wire v$G16_18782_out0;
wire v$G16_3022_out0;
wire v$G16_3023_out0;
wire v$G16_3520_out0;
wire v$G16_3521_out0;
wire v$G16_3839_out0;
wire v$G16_4469_out0;
wire v$G16_4470_out0;
wire v$G16_6391_out0;
wire v$G16_6392_out0;
wire v$G16_6407_out0;
wire v$G16_6408_out0;
wire v$G17_11683_out0;
wire v$G17_11684_out0;
wire v$G17_12139_out0;
wire v$G17_12140_out0;
wire v$G17_13831_out0;
wire v$G17_13832_out0;
wire v$G17_14794_out0;
wire v$G17_14795_out0;
wire v$G17_362_out0;
wire v$G17_363_out0;
wire v$G17_5460_out0;
wire v$G17_5461_out0;
wire v$G17_5476_out0;
wire v$G17_5477_out0;
wire v$G17_5521_out0;
wire v$G17_8178_out0;
wire v$G17_8179_out0;
wire v$G17_8180_out0;
wire v$G17_8181_out0;
wire v$G17_8182_out0;
wire v$G17_8183_out0;
wire v$G17_8184_out0;
wire v$G17_8185_out0;
wire v$G17_8186_out0;
wire v$G17_8187_out0;
wire v$G17_8188_out0;
wire v$G17_8189_out0;
wire v$G17_8190_out0;
wire v$G17_8191_out0;
wire v$G17_8192_out0;
wire v$G17_8193_out0;
wire v$G17_8194_out0;
wire v$G17_8195_out0;
wire v$G17_8196_out0;
wire v$G17_8197_out0;
wire v$G17_8198_out0;
wire v$G17_8199_out0;
wire v$G17_8200_out0;
wire v$G17_8201_out0;
wire v$G17_8830_out0;
wire v$G17_8831_out0;
wire v$G17_8894_out0;
wire v$G17_8895_out0;
wire v$G17_9346_out0;
wire v$G17_9347_out0;
wire v$G17_9348_out0;
wire v$G17_9349_out0;
wire v$G17_9350_out0;
wire v$G18_10254_out0;
wire v$G18_10255_out0;
wire v$G18_11028_out0;
wire v$G18_11029_out0;
wire v$G18_12938_out0;
wire v$G18_12939_out0;
wire v$G18_12940_out0;
wire v$G18_12941_out0;
wire v$G18_12942_out0;
wire v$G18_13513_out0;
wire v$G18_13514_out0;
wire v$G18_13600_out0;
wire v$G18_13601_out0;
wire v$G18_18097_out0;
wire v$G18_18098_out0;
wire v$G18_2988_out0;
wire v$G18_2989_out0;
wire v$G18_3399_out0;
wire v$G18_3400_out0;
wire v$G18_4973_out0;
wire v$G18_4974_out0;
wire v$G18_4975_out0;
wire v$G18_4976_out0;
wire v$G18_4977_out0;
wire v$G18_4978_out0;
wire v$G18_4979_out0;
wire v$G18_4980_out0;
wire v$G18_4981_out0;
wire v$G18_4982_out0;
wire v$G18_4983_out0;
wire v$G18_4984_out0;
wire v$G18_4985_out0;
wire v$G18_4986_out0;
wire v$G18_4987_out0;
wire v$G18_4988_out0;
wire v$G18_4989_out0;
wire v$G18_4990_out0;
wire v$G18_4991_out0;
wire v$G18_4992_out0;
wire v$G18_4993_out0;
wire v$G18_4994_out0;
wire v$G18_4995_out0;
wire v$G18_4996_out0;
wire v$G18_7510_out0;
wire v$G18_8420_out0;
wire v$G18_8421_out0;
wire v$G19_10246_out0;
wire v$G19_10247_out0;
wire v$G19_10248_out0;
wire v$G19_10249_out0;
wire v$G19_13997_out0;
wire v$G19_13998_out0;
wire v$G19_15874_out0;
wire v$G19_15875_out0;
wire v$G19_15948_out0;
wire v$G19_15949_out0;
wire v$G19_16043_out0;
wire v$G19_16044_out0;
wire v$G19_16696_out0;
wire v$G19_16697_out0;
wire v$G19_1881_out0;
wire v$G19_1882_out0;
wire v$G19_1883_out0;
wire v$G19_1884_out0;
wire v$G19_1885_out0;
wire v$G19_2412_out0;
wire v$G19_2413_out0;
wire v$G19_2826_out0;
wire v$G19_2827_out0;
wire v$G19_336_out0;
wire v$G19_337_out0;
wire v$G19_8261_out0;
wire v$G19_8262_out0;
wire v$G1_10317_out0;
wire v$G1_10318_out0;
wire v$G1_1195_out0;
wire v$G1_1196_out0;
wire v$G1_12124_out0;
wire v$G1_12125_out0;
wire v$G1_12223_out0;
wire v$G1_12335_out0;
wire v$G1_12336_out0;
wire v$G1_12337_out0;
wire v$G1_12338_out0;
wire v$G1_12339_out0;
wire v$G1_12340_out0;
wire v$G1_12341_out0;
wire v$G1_12342_out0;
wire v$G1_12343_out0;
wire v$G1_12344_out0;
wire v$G1_12345_out0;
wire v$G1_12346_out0;
wire v$G1_12347_out0;
wire v$G1_12348_out0;
wire v$G1_12349_out0;
wire v$G1_12350_out0;
wire v$G1_12351_out0;
wire v$G1_12352_out0;
wire v$G1_12353_out0;
wire v$G1_12354_out0;
wire v$G1_12355_out0;
wire v$G1_12356_out0;
wire v$G1_12357_out0;
wire v$G1_12358_out0;
wire v$G1_12359_out0;
wire v$G1_12360_out0;
wire v$G1_12361_out0;
wire v$G1_12362_out0;
wire v$G1_12363_out0;
wire v$G1_12364_out0;
wire v$G1_12365_out0;
wire v$G1_12366_out0;
wire v$G1_12367_out0;
wire v$G1_12368_out0;
wire v$G1_12369_out0;
wire v$G1_12370_out0;
wire v$G1_12371_out0;
wire v$G1_12372_out0;
wire v$G1_12373_out0;
wire v$G1_12374_out0;
wire v$G1_12375_out0;
wire v$G1_12376_out0;
wire v$G1_12377_out0;
wire v$G1_12378_out0;
wire v$G1_12379_out0;
wire v$G1_12380_out0;
wire v$G1_12381_out0;
wire v$G1_12382_out0;
wire v$G1_12383_out0;
wire v$G1_12384_out0;
wire v$G1_12385_out0;
wire v$G1_12386_out0;
wire v$G1_12387_out0;
wire v$G1_12388_out0;
wire v$G1_12389_out0;
wire v$G1_12390_out0;
wire v$G1_12391_out0;
wire v$G1_12392_out0;
wire v$G1_12393_out0;
wire v$G1_12394_out0;
wire v$G1_12395_out0;
wire v$G1_12396_out0;
wire v$G1_12397_out0;
wire v$G1_12398_out0;
wire v$G1_12399_out0;
wire v$G1_12400_out0;
wire v$G1_12401_out0;
wire v$G1_12402_out0;
wire v$G1_12403_out0;
wire v$G1_12404_out0;
wire v$G1_12405_out0;
wire v$G1_12406_out0;
wire v$G1_12407_out0;
wire v$G1_12408_out0;
wire v$G1_12409_out0;
wire v$G1_12410_out0;
wire v$G1_12411_out0;
wire v$G1_12412_out0;
wire v$G1_12413_out0;
wire v$G1_12414_out0;
wire v$G1_12415_out0;
wire v$G1_12416_out0;
wire v$G1_12417_out0;
wire v$G1_12418_out0;
wire v$G1_12419_out0;
wire v$G1_12420_out0;
wire v$G1_12421_out0;
wire v$G1_12422_out0;
wire v$G1_12423_out0;
wire v$G1_12424_out0;
wire v$G1_12425_out0;
wire v$G1_12426_out0;
wire v$G1_12427_out0;
wire v$G1_12428_out0;
wire v$G1_12429_out0;
wire v$G1_12430_out0;
wire v$G1_12431_out0;
wire v$G1_12432_out0;
wire v$G1_12433_out0;
wire v$G1_12434_out0;
wire v$G1_12435_out0;
wire v$G1_12436_out0;
wire v$G1_12437_out0;
wire v$G1_12438_out0;
wire v$G1_12439_out0;
wire v$G1_12440_out0;
wire v$G1_12441_out0;
wire v$G1_12442_out0;
wire v$G1_12443_out0;
wire v$G1_12444_out0;
wire v$G1_12445_out0;
wire v$G1_12446_out0;
wire v$G1_12447_out0;
wire v$G1_12448_out0;
wire v$G1_12449_out0;
wire v$G1_12450_out0;
wire v$G1_12451_out0;
wire v$G1_12452_out0;
wire v$G1_12453_out0;
wire v$G1_12454_out0;
wire v$G1_1249_out0;
wire v$G1_1250_out0;
wire v$G1_12982_out0;
wire v$G1_12983_out0;
wire v$G1_12984_out0;
wire v$G1_12985_out0;
wire v$G1_12986_out0;
wire v$G1_13147_out0;
wire v$G1_13148_out0;
wire v$G1_13188_out0;
wire v$G1_13189_out0;
wire v$G1_13190_out0;
wire v$G1_13191_out0;
wire v$G1_13546_out0;
wire v$G1_13547_out0;
wire v$G1_14410_out0;
wire v$G1_14473_out0;
wire v$G1_14474_out0;
wire v$G1_14591_out0;
wire v$G1_14592_out0;
wire v$G1_14593_out0;
wire v$G1_14594_out0;
wire v$G1_14595_out0;
wire v$G1_14596_out0;
wire v$G1_14597_out0;
wire v$G1_14598_out0;
wire v$G1_15142_out0;
wire v$G1_15143_out0;
wire v$G1_15293_out0;
wire v$G1_15294_out0;
wire v$G1_15586_out0;
wire v$G1_15587_out0;
wire v$G1_15782_out0;
wire v$G1_15783_out0;
wire v$G1_1592_out0;
wire v$G1_1593_out0;
wire v$G1_16029_out0;
wire v$G1_16030_out0;
wire v$G1_16031_out0;
wire v$G1_16032_out0;
wire v$G1_16033_out0;
wire v$G1_16034_out0;
wire v$G1_16035_out0;
wire v$G1_16036_out0;
wire v$G1_16141_out0;
wire v$G1_16142_out0;
wire v$G1_16143_out0;
wire v$G1_16144_out0;
wire v$G1_16145_out0;
wire v$G1_16146_out0;
wire v$G1_16147_out0;
wire v$G1_16148_out0;
wire v$G1_16401_out0;
wire v$G1_16402_out0;
wire v$G1_16496_out0;
wire v$G1_16497_out0;
wire v$G1_166_out0;
wire v$G1_167_out0;
wire v$G1_17016_out0;
wire v$G1_17017_out0;
wire v$G1_17446_out0;
wire v$G1_17447_out0;
wire v$G1_17448_out0;
wire v$G1_17449_out0;
wire v$G1_17887_out0;
wire v$G1_17888_out0;
wire v$G1_18647_out0;
wire v$G1_18648_out0;
wire v$G1_1915_out0;
wire v$G1_1916_out0;
wire v$G1_33_out0;
wire v$G1_34_out0;
wire v$G1_4213_out0;
wire v$G1_4214_out0;
wire v$G1_5053_out0;
wire v$G1_5054_out0;
wire v$G1_5055_out0;
wire v$G1_5056_out0;
wire v$G1_5057_out0;
wire v$G1_5421_out0;
wire v$G1_5422_out0;
wire v$G1_5522_out0;
wire v$G1_5523_out0;
wire v$G1_5524_out0;
wire v$G1_5525_out0;
wire v$G1_5526_out0;
wire v$G1_5527_out0;
wire v$G1_5528_out0;
wire v$G1_5529_out0;
wire v$G1_5530_out0;
wire v$G1_5531_out0;
wire v$G1_5532_out0;
wire v$G1_5533_out0;
wire v$G1_5534_out0;
wire v$G1_5535_out0;
wire v$G1_5536_out0;
wire v$G1_5537_out0;
wire v$G1_5538_out0;
wire v$G1_5539_out0;
wire v$G1_5540_out0;
wire v$G1_5541_out0;
wire v$G1_5542_out0;
wire v$G1_5543_out0;
wire v$G1_5544_out0;
wire v$G1_5545_out0;
wire v$G1_5546_out0;
wire v$G1_5547_out0;
wire v$G1_5548_out0;
wire v$G1_5549_out0;
wire v$G1_5550_out0;
wire v$G1_5551_out0;
wire v$G1_5552_out0;
wire v$G1_5553_out0;
wire v$G1_5554_out0;
wire v$G1_5555_out0;
wire v$G1_5556_out0;
wire v$G1_5557_out0;
wire v$G1_5558_out0;
wire v$G1_5559_out0;
wire v$G1_5560_out0;
wire v$G1_5561_out0;
wire v$G1_5562_out0;
wire v$G1_5563_out0;
wire v$G1_5564_out0;
wire v$G1_5565_out0;
wire v$G1_5566_out0;
wire v$G1_5567_out0;
wire v$G1_5568_out0;
wire v$G1_5569_out0;
wire v$G1_5570_out0;
wire v$G1_5571_out0;
wire v$G1_5572_out0;
wire v$G1_5573_out0;
wire v$G1_5574_out0;
wire v$G1_5575_out0;
wire v$G1_5576_out0;
wire v$G1_5577_out0;
wire v$G1_5578_out0;
wire v$G1_5579_out0;
wire v$G1_5580_out0;
wire v$G1_5581_out0;
wire v$G1_5582_out0;
wire v$G1_5583_out0;
wire v$G1_5584_out0;
wire v$G1_5585_out0;
wire v$G1_5586_out0;
wire v$G1_5587_out0;
wire v$G1_5588_out0;
wire v$G1_5589_out0;
wire v$G1_5590_out0;
wire v$G1_5591_out0;
wire v$G1_5592_out0;
wire v$G1_5593_out0;
wire v$G1_5594_out0;
wire v$G1_5595_out0;
wire v$G1_5596_out0;
wire v$G1_5597_out0;
wire v$G1_5598_out0;
wire v$G1_5599_out0;
wire v$G1_5600_out0;
wire v$G1_5601_out0;
wire v$G1_5602_out0;
wire v$G1_5603_out0;
wire v$G1_5604_out0;
wire v$G1_5605_out0;
wire v$G1_5606_out0;
wire v$G1_5607_out0;
wire v$G1_5608_out0;
wire v$G1_5609_out0;
wire v$G1_5610_out0;
wire v$G1_5611_out0;
wire v$G1_5612_out0;
wire v$G1_5613_out0;
wire v$G1_5614_out0;
wire v$G1_5615_out0;
wire v$G1_5616_out0;
wire v$G1_5617_out0;
wire v$G1_5618_out0;
wire v$G1_5619_out0;
wire v$G1_5620_out0;
wire v$G1_5621_out0;
wire v$G1_5622_out0;
wire v$G1_5623_out0;
wire v$G1_5624_out0;
wire v$G1_5625_out0;
wire v$G1_5626_out0;
wire v$G1_5627_out0;
wire v$G1_5628_out0;
wire v$G1_5629_out0;
wire v$G1_5630_out0;
wire v$G1_5631_out0;
wire v$G1_5632_out0;
wire v$G1_5633_out0;
wire v$G1_5634_out0;
wire v$G1_5635_out0;
wire v$G1_5636_out0;
wire v$G1_5637_out0;
wire v$G1_5638_out0;
wire v$G1_5639_out0;
wire v$G1_5640_out0;
wire v$G1_5641_out0;
wire v$G1_5642_out0;
wire v$G1_5643_out0;
wire v$G1_5644_out0;
wire v$G1_5645_out0;
wire v$G1_5646_out0;
wire v$G1_5647_out0;
wire v$G1_5648_out0;
wire v$G1_5649_out0;
wire v$G1_5650_out0;
wire v$G1_5651_out0;
wire v$G1_5652_out0;
wire v$G1_5653_out0;
wire v$G1_5654_out0;
wire v$G1_5655_out0;
wire v$G1_5656_out0;
wire v$G1_5657_out0;
wire v$G1_5658_out0;
wire v$G1_5659_out0;
wire v$G1_5660_out0;
wire v$G1_5661_out0;
wire v$G1_5662_out0;
wire v$G1_5663_out0;
wire v$G1_5664_out0;
wire v$G1_5665_out0;
wire v$G1_5666_out0;
wire v$G1_5667_out0;
wire v$G1_5668_out0;
wire v$G1_5669_out0;
wire v$G1_5670_out0;
wire v$G1_5671_out0;
wire v$G1_5672_out0;
wire v$G1_5673_out0;
wire v$G1_5674_out0;
wire v$G1_5675_out0;
wire v$G1_5676_out0;
wire v$G1_5677_out0;
wire v$G1_5678_out0;
wire v$G1_5679_out0;
wire v$G1_5680_out0;
wire v$G1_5681_out0;
wire v$G1_5682_out0;
wire v$G1_5683_out0;
wire v$G1_5684_out0;
wire v$G1_5685_out0;
wire v$G1_5686_out0;
wire v$G1_5687_out0;
wire v$G1_5688_out0;
wire v$G1_5689_out0;
wire v$G1_5690_out0;
wire v$G1_5691_out0;
wire v$G1_5692_out0;
wire v$G1_5693_out0;
wire v$G1_5694_out0;
wire v$G1_5695_out0;
wire v$G1_5696_out0;
wire v$G1_5697_out0;
wire v$G1_5698_out0;
wire v$G1_5699_out0;
wire v$G1_5700_out0;
wire v$G1_5701_out0;
wire v$G1_5702_out0;
wire v$G1_5703_out0;
wire v$G1_5704_out0;
wire v$G1_5705_out0;
wire v$G1_5706_out0;
wire v$G1_5707_out0;
wire v$G1_5708_out0;
wire v$G1_5709_out0;
wire v$G1_5710_out0;
wire v$G1_5711_out0;
wire v$G1_5712_out0;
wire v$G1_5713_out0;
wire v$G1_5714_out0;
wire v$G1_5715_out0;
wire v$G1_5716_out0;
wire v$G1_5717_out0;
wire v$G1_5718_out0;
wire v$G1_5719_out0;
wire v$G1_5720_out0;
wire v$G1_5721_out0;
wire v$G1_5722_out0;
wire v$G1_5723_out0;
wire v$G1_5724_out0;
wire v$G1_5725_out0;
wire v$G1_5726_out0;
wire v$G1_7223_out0;
wire v$G1_7224_out0;
wire v$G1_7325_out0;
wire v$G1_7326_out0;
wire v$G1_7333_out0;
wire v$G1_8792_out0;
wire v$G1_8793_out0;
wire v$G1_8794_out0;
wire v$G1_8795_out0;
wire v$G1_9386_out0;
wire v$G1_9387_out0;
wire v$G1_9388_out0;
wire v$G1_9389_out0;
wire v$G1_9390_out0;
wire v$G1_9391_out0;
wire v$G1_9392_out0;
wire v$G1_9393_out0;
wire v$G20_11710_out0;
wire v$G20_11711_out0;
wire v$G20_12209_out0;
wire v$G20_12210_out0;
wire v$G20_12292_out0;
wire v$G20_12293_out0;
wire v$G20_12740_out0;
wire v$G20_12741_out0;
wire v$G20_15936_out0;
wire v$G20_15937_out0;
wire v$G20_18281_out0;
wire v$G20_18282_out0;
wire v$G20_2594_out0;
wire v$G20_2595_out0;
wire v$G20_5451_out0;
wire v$G20_5452_out0;
wire v$G20_7402_out0;
wire v$G20_7403_out0;
wire v$G20_8225_out0;
wire v$G20_8226_out0;
wire v$G20_8227_out0;
wire v$G20_8228_out0;
wire v$G20_8229_out0;
wire v$G20_9882_out0;
wire v$G20_9883_out0;
wire v$G20_9884_out0;
wire v$G20_9885_out0;
wire v$G20_9886_out0;
wire v$G20_9887_out0;
wire v$G20_9888_out0;
wire v$G20_9889_out0;
wire v$G20_9890_out0;
wire v$G20_9891_out0;
wire v$G20_9892_out0;
wire v$G20_9893_out0;
wire v$G20_9894_out0;
wire v$G20_9895_out0;
wire v$G20_9896_out0;
wire v$G20_9897_out0;
wire v$G20_9898_out0;
wire v$G20_9899_out0;
wire v$G20_9900_out0;
wire v$G20_9901_out0;
wire v$G20_9902_out0;
wire v$G20_9903_out0;
wire v$G20_9904_out0;
wire v$G20_9905_out0;
wire v$G21_11874_out0;
wire v$G21_11875_out0;
wire v$G21_14017_out0;
wire v$G21_14018_out0;
wire v$G21_14019_out0;
wire v$G21_14020_out0;
wire v$G21_14021_out0;
wire v$G21_14245_out0;
wire v$G21_14246_out0;
wire v$G21_14710_out0;
wire v$G21_14711_out0;
wire v$G21_15312_out0;
wire v$G21_15313_out0;
wire v$G21_15822_out0;
wire v$G21_15823_out0;
wire v$G21_17674_out0;
wire v$G21_17675_out0;
wire v$G21_18680_out0;
wire v$G21_18681_out0;
wire v$G21_3522_out0;
wire v$G21_3523_out0;
wire v$G21_3524_out0;
wire v$G21_3525_out0;
wire v$G21_3526_out0;
wire v$G21_3527_out0;
wire v$G21_3528_out0;
wire v$G21_3529_out0;
wire v$G21_3530_out0;
wire v$G21_3531_out0;
wire v$G21_3532_out0;
wire v$G21_3533_out0;
wire v$G21_3534_out0;
wire v$G21_3535_out0;
wire v$G21_3536_out0;
wire v$G21_3537_out0;
wire v$G21_3538_out0;
wire v$G21_3539_out0;
wire v$G21_3540_out0;
wire v$G21_3541_out0;
wire v$G21_3542_out0;
wire v$G21_3543_out0;
wire v$G21_3544_out0;
wire v$G21_3545_out0;
wire v$G21_7036_out0;
wire v$G21_7037_out0;
wire v$G21_7484_out0;
wire v$G21_7485_out0;
wire v$G22_12510_out0;
wire v$G22_12511_out0;
wire v$G22_12512_out0;
wire v$G22_12513_out0;
wire v$G22_12514_out0;
wire v$G22_13327_out0;
wire v$G22_13328_out0;
wire v$G22_13329_out0;
wire v$G22_13330_out0;
wire v$G22_13331_out0;
wire v$G22_13332_out0;
wire v$G22_13333_out0;
wire v$G22_13334_out0;
wire v$G22_13335_out0;
wire v$G22_13336_out0;
wire v$G22_13337_out0;
wire v$G22_13338_out0;
wire v$G22_13339_out0;
wire v$G22_13340_out0;
wire v$G22_13341_out0;
wire v$G22_13342_out0;
wire v$G22_13343_out0;
wire v$G22_13344_out0;
wire v$G22_13345_out0;
wire v$G22_13346_out0;
wire v$G22_13347_out0;
wire v$G22_13348_out0;
wire v$G22_13349_out0;
wire v$G22_13350_out0;
wire v$G22_15342_out0;
wire v$G22_15343_out0;
wire v$G22_15631_out0;
wire v$G22_15632_out0;
wire v$G22_15852_out0;
wire v$G22_15853_out0;
wire v$G22_4313_out0;
wire v$G22_4314_out0;
wire v$G22_4882_out0;
wire v$G22_4883_out0;
wire v$G22_5462_out0;
wire v$G22_5463_out0;
wire v$G22_7267_out0;
wire v$G22_7268_out0;
wire v$G23_12175_out0;
wire v$G23_12176_out0;
wire v$G23_12177_out0;
wire v$G23_12178_out0;
wire v$G23_12179_out0;
wire v$G23_12180_out0;
wire v$G23_12181_out0;
wire v$G23_12182_out0;
wire v$G23_12183_out0;
wire v$G23_12184_out0;
wire v$G23_12185_out0;
wire v$G23_12186_out0;
wire v$G23_12187_out0;
wire v$G23_12188_out0;
wire v$G23_12189_out0;
wire v$G23_12190_out0;
wire v$G23_12191_out0;
wire v$G23_12192_out0;
wire v$G23_12193_out0;
wire v$G23_12194_out0;
wire v$G23_12195_out0;
wire v$G23_12196_out0;
wire v$G23_12197_out0;
wire v$G23_12198_out0;
wire v$G23_14080_out0;
wire v$G23_14081_out0;
wire v$G23_14317_out0;
wire v$G23_14318_out0;
wire v$G23_14319_out0;
wire v$G23_14320_out0;
wire v$G23_14321_out0;
wire v$G23_15947_out0;
wire v$G23_16770_out0;
wire v$G23_16771_out0;
wire v$G23_17687_out0;
wire v$G23_17688_out0;
wire v$G23_18654_out0;
wire v$G23_18655_out0;
wire v$G23_2277_out0;
wire v$G23_2278_out0;
wire v$G23_4385_out0;
wire v$G23_4386_out0;
wire v$G23_6992_out0;
wire v$G23_6993_out0;
wire v$G23_9360_out0;
wire v$G23_9361_out0;
wire v$G23_9601_out0;
wire v$G23_9602_out0;
wire v$G24_10343_out0;
wire v$G24_10344_out0;
wire v$G24_12087_out0;
wire v$G24_12088_out0;
wire v$G24_13860_out0;
wire v$G24_13861_out0;
wire v$G24_15684_out0;
wire v$G24_15685_out0;
wire v$G24_15686_out0;
wire v$G24_15687_out0;
wire v$G24_15688_out0;
wire v$G24_15689_out0;
wire v$G24_15690_out0;
wire v$G24_15691_out0;
wire v$G24_15692_out0;
wire v$G24_15693_out0;
wire v$G24_15694_out0;
wire v$G24_15695_out0;
wire v$G24_15696_out0;
wire v$G24_15697_out0;
wire v$G24_15698_out0;
wire v$G24_15699_out0;
wire v$G24_15700_out0;
wire v$G24_15701_out0;
wire v$G24_15702_out0;
wire v$G24_15703_out0;
wire v$G24_15704_out0;
wire v$G24_15705_out0;
wire v$G24_15706_out0;
wire v$G24_15707_out0;
wire v$G24_17018_out0;
wire v$G24_17019_out0;
wire v$G24_17931_out0;
wire v$G24_17932_out0;
wire v$G24_18388_out0;
wire v$G24_18389_out0;
wire v$G24_240_out0;
wire v$G24_3401_out0;
wire v$G24_3402_out0;
wire v$G24_672_out0;
wire v$G24_673_out0;
wire v$G24_7896_out0;
wire v$G24_7897_out0;
wire v$G24_9618_out0;
wire v$G24_9619_out0;
wire v$G25_10273_out0;
wire v$G25_10934_out0;
wire v$G25_10935_out0;
wire v$G25_10936_out0;
wire v$G25_10937_out0;
wire v$G25_10938_out0;
wire v$G25_10939_out0;
wire v$G25_10940_out0;
wire v$G25_10941_out0;
wire v$G25_10942_out0;
wire v$G25_10943_out0;
wire v$G25_10944_out0;
wire v$G25_10945_out0;
wire v$G25_10946_out0;
wire v$G25_10947_out0;
wire v$G25_10948_out0;
wire v$G25_10949_out0;
wire v$G25_10950_out0;
wire v$G25_10951_out0;
wire v$G25_10952_out0;
wire v$G25_10953_out0;
wire v$G25_10954_out0;
wire v$G25_10955_out0;
wire v$G25_10956_out0;
wire v$G25_10957_out0;
wire v$G25_12754_out0;
wire v$G25_12755_out0;
wire v$G25_13011_out0;
wire v$G25_13012_out0;
wire v$G25_1309_out0;
wire v$G25_1310_out0;
wire v$G25_14030_out0;
wire v$G25_14031_out0;
wire v$G25_14578_out0;
wire v$G25_14579_out0;
wire v$G25_14659_out0;
wire v$G25_14660_out0;
wire v$G25_16104_out0;
wire v$G25_16105_out0;
wire v$G25_18095_out0;
wire v$G25_18096_out0;
wire v$G25_2464_out0;
wire v$G25_2465_out0;
wire v$G25_3549_out0;
wire v$G25_3550_out0;
wire v$G26_10319_out0;
wire v$G26_10320_out0;
wire v$G26_11368_out0;
wire v$G26_11369_out0;
wire v$G26_11370_out0;
wire v$G26_11371_out0;
wire v$G26_12654_out0;
wire v$G26_12655_out0;
wire v$G26_13177_out0;
wire v$G26_13178_out0;
wire v$G26_13641_out0;
wire v$G26_13642_out0;
wire v$G26_14899_out0;
wire v$G26_14900_out0;
wire v$G26_16019_out0;
wire v$G26_16020_out0;
wire v$G26_16025_out0;
wire v$G26_16026_out0;
wire v$G26_18115_out0;
wire v$G26_4097_out0;
wire v$G26_4098_out0;
wire v$G26_5127_out0;
wire v$G27_10235_out0;
wire v$G27_10236_out0;
wire v$G27_10726_out0;
wire v$G27_11706_out0;
wire v$G27_11707_out0;
wire v$G27_11708_out0;
wire v$G27_11709_out0;
wire v$G27_16528_out0;
wire v$G27_16529_out0;
wire v$G27_18489_out0;
wire v$G27_18490_out0;
wire v$G27_2512_out0;
wire v$G27_2513_out0;
wire v$G27_260_out0;
wire v$G27_261_out0;
wire v$G27_3882_out0;
wire v$G27_4776_out0;
wire v$G27_4777_out0;
wire v$G27_4778_out0;
wire v$G27_4779_out0;
wire v$G27_4780_out0;
wire v$G27_4781_out0;
wire v$G27_4782_out0;
wire v$G27_4783_out0;
wire v$G27_4784_out0;
wire v$G27_4785_out0;
wire v$G27_4786_out0;
wire v$G27_4787_out0;
wire v$G27_4788_out0;
wire v$G27_4789_out0;
wire v$G27_4790_out0;
wire v$G27_4791_out0;
wire v$G27_4792_out0;
wire v$G27_4793_out0;
wire v$G27_4794_out0;
wire v$G27_4795_out0;
wire v$G27_4796_out0;
wire v$G27_4797_out0;
wire v$G27_4798_out0;
wire v$G27_4799_out0;
wire v$G28_10803_out0;
wire v$G28_10804_out0;
wire v$G28_11939_out0;
wire v$G28_11940_out0;
wire v$G28_13015_out0;
wire v$G28_13016_out0;
wire v$G28_13017_out0;
wire v$G28_13018_out0;
wire v$G28_13019_out0;
wire v$G28_13020_out0;
wire v$G28_13021_out0;
wire v$G28_13022_out0;
wire v$G28_13023_out0;
wire v$G28_13024_out0;
wire v$G28_13025_out0;
wire v$G28_13026_out0;
wire v$G28_13027_out0;
wire v$G28_13028_out0;
wire v$G28_13029_out0;
wire v$G28_13030_out0;
wire v$G28_13031_out0;
wire v$G28_13032_out0;
wire v$G28_13033_out0;
wire v$G28_13034_out0;
wire v$G28_13035_out0;
wire v$G28_13036_out0;
wire v$G28_13037_out0;
wire v$G28_13038_out0;
wire v$G28_13787_out0;
wire v$G28_14668_out0;
wire v$G28_14669_out0;
wire v$G28_15384_out0;
wire v$G28_15385_out0;
wire v$G28_15633_out0;
wire v$G28_15634_out0;
wire v$G28_18550_out0;
wire v$G28_18551_out0;
wire v$G28_3167_out0;
wire v$G28_3168_out0;
wire v$G28_3765_out0;
wire v$G28_3766_out0;
wire v$G28_8690_out0;
wire v$G29_10298_out0;
wire v$G29_10299_out0;
wire v$G29_10300_out0;
wire v$G29_10301_out0;
wire v$G29_10829_out0;
wire v$G29_13993_out0;
wire v$G29_13994_out0;
wire v$G29_15774_out0;
wire v$G29_15775_out0;
wire v$G29_3624_out0;
wire v$G29_3625_out0;
wire v$G29_5485_out0;
wire v$G29_5486_out0;
wire v$G29_681_out0;
wire v$G29_682_out0;
wire v$G29_7465_out0;
wire v$G29_7466_out0;
wire v$G29_7851_out0;
wire v$G29_7852_out0;
wire v$G2_10400_out0;
wire v$G2_10401_out0;
wire v$G2_10402_out0;
wire v$G2_10403_out0;
wire v$G2_11697_out0;
wire v$G2_11902_out0;
wire v$G2_11903_out0;
wire v$G2_11904_out0;
wire v$G2_11905_out0;
wire v$G2_1288_out0;
wire v$G2_1289_out0;
wire v$G2_12904_out0;
wire v$G2_12905_out0;
wire v$G2_12906_out0;
wire v$G2_12907_out0;
wire v$G2_12908_out0;
wire v$G2_12909_out0;
wire v$G2_12910_out0;
wire v$G2_12911_out0;
wire v$G2_13693_out0;
wire v$G2_13694_out0;
wire v$G2_14499_out0;
wire v$G2_14500_out0;
wire v$G2_15033_out0;
wire v$G2_15034_out0;
wire v$G2_15035_out0;
wire v$G2_15036_out0;
wire v$G2_15037_out0;
wire v$G2_15038_out0;
wire v$G2_15039_out0;
wire v$G2_15040_out0;
wire v$G2_15041_out0;
wire v$G2_15042_out0;
wire v$G2_15043_out0;
wire v$G2_15044_out0;
wire v$G2_15542_out0;
wire v$G2_15543_out0;
wire v$G2_15761_out0;
wire v$G2_15762_out0;
wire v$G2_15863_out0;
wire v$G2_15864_out0;
wire v$G2_15960_out0;
wire v$G2_15961_out0;
wire v$G2_15962_out0;
wire v$G2_15963_out0;
wire v$G2_15964_out0;
wire v$G2_16502_out0;
wire v$G2_16503_out0;
wire v$G2_17064_out0;
wire v$G2_17065_out0;
wire v$G2_17411_out0;
wire v$G2_17412_out0;
wire v$G2_17413_out0;
wire v$G2_17414_out0;
wire v$G2_17415_out0;
wire v$G2_17416_out0;
wire v$G2_17417_out0;
wire v$G2_17418_out0;
wire v$G2_17663_out0;
wire v$G2_17664_out0;
wire v$G2_18239_out0;
wire v$G2_18240_out0;
wire v$G2_18241_out0;
wire v$G2_18242_out0;
wire v$G2_18429_out0;
wire v$G2_18430_out0;
wire v$G2_18697_out0;
wire v$G2_18698_out0;
wire v$G2_1894_out0;
wire v$G2_1895_out0;
wire v$G2_2425_out0;
wire v$G2_2426_out0;
wire v$G2_3724_out0;
wire v$G2_3725_out0;
wire v$G2_4089_out0;
wire v$G2_4090_out0;
wire v$G2_5047_out0;
wire v$G2_5048_out0;
wire v$G2_5253_out0;
wire v$G2_5254_out0;
wire v$G2_5261_out0;
wire v$G2_5262_out0;
wire v$G2_5263_out0;
wire v$G2_5264_out0;
wire v$G2_5265_out0;
wire v$G2_5266_out0;
wire v$G2_5267_out0;
wire v$G2_5268_out0;
wire v$G2_5269_out0;
wire v$G2_5270_out0;
wire v$G2_5271_out0;
wire v$G2_5272_out0;
wire v$G2_5273_out0;
wire v$G2_5274_out0;
wire v$G2_5275_out0;
wire v$G2_5276_out0;
wire v$G2_5277_out0;
wire v$G2_5278_out0;
wire v$G2_5279_out0;
wire v$G2_5280_out0;
wire v$G2_5281_out0;
wire v$G2_5282_out0;
wire v$G2_5283_out0;
wire v$G2_5284_out0;
wire v$G2_5285_out0;
wire v$G2_5286_out0;
wire v$G2_5287_out0;
wire v$G2_5288_out0;
wire v$G2_5289_out0;
wire v$G2_5290_out0;
wire v$G2_5291_out0;
wire v$G2_5292_out0;
wire v$G2_5293_out0;
wire v$G2_5294_out0;
wire v$G2_5295_out0;
wire v$G2_5296_out0;
wire v$G2_5297_out0;
wire v$G2_5298_out0;
wire v$G2_5299_out0;
wire v$G2_5300_out0;
wire v$G2_5301_out0;
wire v$G2_5302_out0;
wire v$G2_5303_out0;
wire v$G2_5304_out0;
wire v$G2_5305_out0;
wire v$G2_5306_out0;
wire v$G2_5307_out0;
wire v$G2_5308_out0;
wire v$G2_5309_out0;
wire v$G2_5310_out0;
wire v$G2_5311_out0;
wire v$G2_5312_out0;
wire v$G2_5313_out0;
wire v$G2_5314_out0;
wire v$G2_5315_out0;
wire v$G2_5316_out0;
wire v$G2_5317_out0;
wire v$G2_5318_out0;
wire v$G2_5319_out0;
wire v$G2_5320_out0;
wire v$G2_5321_out0;
wire v$G2_5322_out0;
wire v$G2_5323_out0;
wire v$G2_5324_out0;
wire v$G2_5325_out0;
wire v$G2_5326_out0;
wire v$G2_5327_out0;
wire v$G2_5328_out0;
wire v$G2_5329_out0;
wire v$G2_5330_out0;
wire v$G2_5331_out0;
wire v$G2_5332_out0;
wire v$G2_5333_out0;
wire v$G2_5334_out0;
wire v$G2_5335_out0;
wire v$G2_5336_out0;
wire v$G2_5337_out0;
wire v$G2_5338_out0;
wire v$G2_5339_out0;
wire v$G2_5340_out0;
wire v$G2_5341_out0;
wire v$G2_5342_out0;
wire v$G2_5343_out0;
wire v$G2_5344_out0;
wire v$G2_5345_out0;
wire v$G2_5346_out0;
wire v$G2_5347_out0;
wire v$G2_5348_out0;
wire v$G2_5349_out0;
wire v$G2_5350_out0;
wire v$G2_5351_out0;
wire v$G2_5352_out0;
wire v$G2_5353_out0;
wire v$G2_5354_out0;
wire v$G2_5355_out0;
wire v$G2_5356_out0;
wire v$G2_5357_out0;
wire v$G2_5358_out0;
wire v$G2_5359_out0;
wire v$G2_5360_out0;
wire v$G2_5361_out0;
wire v$G2_5362_out0;
wire v$G2_5363_out0;
wire v$G2_5364_out0;
wire v$G2_5365_out0;
wire v$G2_5366_out0;
wire v$G2_5367_out0;
wire v$G2_5368_out0;
wire v$G2_5369_out0;
wire v$G2_5370_out0;
wire v$G2_5371_out0;
wire v$G2_5372_out0;
wire v$G2_5373_out0;
wire v$G2_5374_out0;
wire v$G2_5375_out0;
wire v$G2_5376_out0;
wire v$G2_5377_out0;
wire v$G2_5378_out0;
wire v$G2_5379_out0;
wire v$G2_5380_out0;
wire v$G2_5429_out0;
wire v$G2_5430_out0;
wire v$G2_65_out0;
wire v$G2_66_out0;
wire v$G2_7562_out0;
wire v$G2_7574_out0;
wire v$G2_7575_out0;
wire v$G2_7576_out0;
wire v$G2_7577_out0;
wire v$G2_7578_out0;
wire v$G2_7777_out0;
wire v$G2_7778_out0;
wire v$G2_8130_out0;
wire v$G2_8334_out0;
wire v$G2_8335_out0;
wire v$G2_9078_out0;
wire v$G2_9079_out0;
wire v$G30_15903_out0;
wire v$G30_15904_out0;
wire v$G30_1717_out0;
wire v$G30_1718_out0;
wire v$G30_1769_out0;
wire v$G30_1770_out0;
wire v$G30_1771_out0;
wire v$G30_1772_out0;
wire v$G30_1773_out0;
wire v$G30_1774_out0;
wire v$G30_1775_out0;
wire v$G30_1776_out0;
wire v$G30_1777_out0;
wire v$G30_1778_out0;
wire v$G30_1779_out0;
wire v$G30_1780_out0;
wire v$G30_1781_out0;
wire v$G30_1782_out0;
wire v$G30_1783_out0;
wire v$G30_1784_out0;
wire v$G30_1785_out0;
wire v$G30_1786_out0;
wire v$G30_1787_out0;
wire v$G30_1788_out0;
wire v$G30_1789_out0;
wire v$G30_1790_out0;
wire v$G30_1791_out0;
wire v$G30_1792_out0;
wire v$G30_18605_out0;
wire v$G30_18606_out0;
wire v$G30_2466_out0;
wire v$G30_2467_out0;
wire v$G30_3764_out0;
wire v$G30_4923_out0;
wire v$G30_4924_out0;
wire v$G31_10793_out0;
wire v$G31_10794_out0;
wire v$G31_15506_out0;
wire v$G31_15507_out0;
wire v$G31_15508_out0;
wire v$G31_15509_out0;
wire v$G31_15510_out0;
wire v$G31_15511_out0;
wire v$G31_15512_out0;
wire v$G31_15513_out0;
wire v$G31_15514_out0;
wire v$G31_15515_out0;
wire v$G31_15516_out0;
wire v$G31_15517_out0;
wire v$G31_15518_out0;
wire v$G31_15519_out0;
wire v$G31_15520_out0;
wire v$G31_15521_out0;
wire v$G31_15522_out0;
wire v$G31_15523_out0;
wire v$G31_15524_out0;
wire v$G31_15525_out0;
wire v$G31_15526_out0;
wire v$G31_15527_out0;
wire v$G31_15528_out0;
wire v$G31_15529_out0;
wire v$G31_1822_out0;
wire v$G31_1823_out0;
wire v$G31_18635_out0;
wire v$G31_18636_out0;
wire v$G31_2344_out0;
wire v$G31_9632_out0;
wire v$G31_9633_out0;
wire v$G32_11884_out0;
wire v$G32_11885_out0;
wire v$G32_14201_out0;
wire v$G32_14202_out0;
wire v$G32_16333_out0;
wire v$G32_16334_out0;
wire v$G32_16335_out0;
wire v$G32_16412_out0;
wire v$G32_16413_out0;
wire v$G32_1826_out0;
wire v$G32_1827_out0;
wire v$G32_392_out0;
wire v$G32_393_out0;
wire v$G32_394_out0;
wire v$G32_395_out0;
wire v$G32_396_out0;
wire v$G32_397_out0;
wire v$G32_398_out0;
wire v$G32_399_out0;
wire v$G32_400_out0;
wire v$G32_401_out0;
wire v$G32_402_out0;
wire v$G32_403_out0;
wire v$G32_404_out0;
wire v$G32_405_out0;
wire v$G32_406_out0;
wire v$G32_407_out0;
wire v$G32_408_out0;
wire v$G32_409_out0;
wire v$G32_410_out0;
wire v$G32_411_out0;
wire v$G32_412_out0;
wire v$G32_413_out0;
wire v$G32_414_out0;
wire v$G32_415_out0;
wire v$G32_9114_out0;
wire v$G32_9115_out0;
wire v$G33_10750_out0;
wire v$G33_10751_out0;
wire v$G33_1233_out0;
wire v$G33_1234_out0;
wire v$G33_13099_out0;
wire v$G33_13100_out0;
wire v$G33_13101_out0;
wire v$G33_13102_out0;
wire v$G33_13103_out0;
wire v$G33_13104_out0;
wire v$G33_13105_out0;
wire v$G33_13106_out0;
wire v$G33_13107_out0;
wire v$G33_13108_out0;
wire v$G33_13109_out0;
wire v$G33_13110_out0;
wire v$G33_13111_out0;
wire v$G33_13112_out0;
wire v$G33_13113_out0;
wire v$G33_13114_out0;
wire v$G33_13115_out0;
wire v$G33_13116_out0;
wire v$G33_13117_out0;
wire v$G33_13118_out0;
wire v$G33_13119_out0;
wire v$G33_13120_out0;
wire v$G33_13121_out0;
wire v$G33_13122_out0;
wire v$G33_18616_out0;
wire v$G33_18617_out0;
wire v$G33_324_out0;
wire v$G33_5131_out0;
wire v$G33_5132_out0;
wire v$G34_1570_out0;
wire v$G34_1571_out0;
wire v$G34_17292_out0;
wire v$G34_17293_out0;
wire v$G34_17294_out0;
wire v$G34_17295_out0;
wire v$G34_17296_out0;
wire v$G34_17297_out0;
wire v$G34_17298_out0;
wire v$G34_17299_out0;
wire v$G34_17300_out0;
wire v$G34_17301_out0;
wire v$G34_17302_out0;
wire v$G34_17303_out0;
wire v$G34_17304_out0;
wire v$G34_17305_out0;
wire v$G34_17306_out0;
wire v$G34_17307_out0;
wire v$G34_17308_out0;
wire v$G34_17309_out0;
wire v$G34_17310_out0;
wire v$G34_17311_out0;
wire v$G34_17312_out0;
wire v$G34_17313_out0;
wire v$G34_17314_out0;
wire v$G34_17315_out0;
wire v$G34_4880_out0;
wire v$G34_4881_out0;
wire v$G34_4917_out0;
wire v$G34_4918_out0;
wire v$G35_10321_out0;
wire v$G35_10322_out0;
wire v$G35_1145_out0;
wire v$G35_1146_out0;
wire v$G35_12635_out0;
wire v$G35_12636_out0;
wire v$G35_14523_out0;
wire v$G35_14524_out0;
wire v$G35_14525_out0;
wire v$G35_14526_out0;
wire v$G35_14527_out0;
wire v$G35_14528_out0;
wire v$G35_14529_out0;
wire v$G35_14530_out0;
wire v$G35_14531_out0;
wire v$G35_14532_out0;
wire v$G35_14533_out0;
wire v$G35_14534_out0;
wire v$G35_14535_out0;
wire v$G35_14536_out0;
wire v$G35_14537_out0;
wire v$G35_14538_out0;
wire v$G35_14539_out0;
wire v$G35_14540_out0;
wire v$G35_14541_out0;
wire v$G35_14542_out0;
wire v$G35_14543_out0;
wire v$G35_14544_out0;
wire v$G35_14545_out0;
wire v$G35_14546_out0;
wire v$G35_18495_out0;
wire v$G35_18496_out0;
wire v$G35_4315_out0;
wire v$G35_4316_out0;
wire v$G36_10864_out0;
wire v$G36_10865_out0;
wire v$G36_14103_out0;
wire v$G36_14104_out0;
wire v$G36_16700_out0;
wire v$G36_17349_out0;
wire v$G36_17350_out0;
wire v$G36_5906_out0;
wire v$G36_5907_out0;
wire v$G36_5908_out0;
wire v$G36_5909_out0;
wire v$G36_5910_out0;
wire v$G36_5911_out0;
wire v$G36_5912_out0;
wire v$G36_5913_out0;
wire v$G36_5914_out0;
wire v$G36_5915_out0;
wire v$G36_5916_out0;
wire v$G36_5917_out0;
wire v$G36_5918_out0;
wire v$G36_5919_out0;
wire v$G36_5920_out0;
wire v$G36_5921_out0;
wire v$G36_5922_out0;
wire v$G36_5923_out0;
wire v$G36_5924_out0;
wire v$G36_5925_out0;
wire v$G36_5926_out0;
wire v$G36_5927_out0;
wire v$G36_5928_out0;
wire v$G36_5929_out0;
wire v$G36_8050_out0;
wire v$G36_8051_out0;
wire v$G37_1360_out0;
wire v$G37_1361_out0;
wire v$G37_14088_out0;
wire v$G37_14089_out0;
wire v$G37_1517_out0;
wire v$G37_1518_out0;
wire v$G37_1519_out0;
wire v$G37_1520_out0;
wire v$G37_18464_out0;
wire v$G37_18465_out0;
wire v$G37_685_out0;
wire v$G37_686_out0;
wire v$G38_10252_out0;
wire v$G38_10253_out0;
wire v$G38_7291_out0;
wire v$G38_7292_out0;
wire v$G38_7293_out0;
wire v$G38_7294_out0;
wire v$G38_7295_out0;
wire v$G38_7296_out0;
wire v$G38_7297_out0;
wire v$G38_7298_out0;
wire v$G38_7299_out0;
wire v$G38_7300_out0;
wire v$G38_7301_out0;
wire v$G38_7302_out0;
wire v$G38_7303_out0;
wire v$G38_7304_out0;
wire v$G38_7305_out0;
wire v$G38_7306_out0;
wire v$G38_7307_out0;
wire v$G38_7308_out0;
wire v$G38_7309_out0;
wire v$G38_7310_out0;
wire v$G38_7311_out0;
wire v$G38_7312_out0;
wire v$G38_7313_out0;
wire v$G38_7314_out0;
wire v$G39_16890_out0;
wire v$G39_16891_out0;
wire v$G39_17358_out0;
wire v$G39_17359_out0;
wire v$G39_17360_out0;
wire v$G39_17361_out0;
wire v$G39_6045_out0;
wire v$G39_6046_out0;
wire v$G3_0_out0;
wire v$G3_10233_out0;
wire v$G3_10234_out0;
wire v$G3_10988_out0;
wire v$G3_10989_out0;
wire v$G3_11104_out0;
wire v$G3_11105_out0;
wire v$G3_11106_out0;
wire v$G3_11107_out0;
wire v$G3_11108_out0;
wire v$G3_12662_out0;
wire v$G3_12663_out0;
wire v$G3_12664_out0;
wire v$G3_12665_out0;
wire v$G3_12666_out0;
wire v$G3_12667_out0;
wire v$G3_12668_out0;
wire v$G3_12669_out0;
wire v$G3_12670_out0;
wire v$G3_12671_out0;
wire v$G3_12672_out0;
wire v$G3_12673_out0;
wire v$G3_12674_out0;
wire v$G3_12675_out0;
wire v$G3_12676_out0;
wire v$G3_12677_out0;
wire v$G3_12678_out0;
wire v$G3_12679_out0;
wire v$G3_12680_out0;
wire v$G3_12681_out0;
wire v$G3_12682_out0;
wire v$G3_12683_out0;
wire v$G3_12684_out0;
wire v$G3_12685_out0;
wire v$G3_12686_out0;
wire v$G3_12687_out0;
wire v$G3_12688_out0;
wire v$G3_12689_out0;
wire v$G3_12690_out0;
wire v$G3_12691_out0;
wire v$G3_12692_out0;
wire v$G3_12693_out0;
wire v$G3_12694_out0;
wire v$G3_12695_out0;
wire v$G3_12696_out0;
wire v$G3_12697_out0;
wire v$G3_12698_out0;
wire v$G3_12699_out0;
wire v$G3_12700_out0;
wire v$G3_12701_out0;
wire v$G3_12702_out0;
wire v$G3_12703_out0;
wire v$G3_12704_out0;
wire v$G3_12705_out0;
wire v$G3_12706_out0;
wire v$G3_12707_out0;
wire v$G3_12708_out0;
wire v$G3_12709_out0;
wire v$G3_12948_out0;
wire v$G3_12949_out0;
wire v$G3_13061_out0;
wire v$G3_13062_out0;
wire v$G3_13063_out0;
wire v$G3_13064_out0;
wire v$G3_14181_out0;
wire v$G3_14182_out0;
wire v$G3_15837_out0;
wire v$G3_15838_out0;
wire v$G3_16009_out0;
wire v$G3_16010_out0;
wire v$G3_16089_out0;
wire v$G3_17452_out0;
wire v$G3_17453_out0;
wire v$G3_17690_out0;
wire v$G3_17691_out0;
wire v$G3_17692_out0;
wire v$G3_17693_out0;
wire v$G3_17694_out0;
wire v$G3_18414_out0;
wire v$G3_18415_out0;
wire v$G3_1_out0;
wire v$G3_20_out0;
wire v$G3_21_out0;
wire v$G3_2441_out0;
wire v$G3_2442_out0;
wire v$G3_2605_out0;
wire v$G3_2606_out0;
wire v$G3_2607_out0;
wire v$G3_2608_out0;
wire v$G3_2609_out0;
wire v$G3_2610_out0;
wire v$G3_2611_out0;
wire v$G3_2612_out0;
wire v$G3_2671_out0;
wire v$G3_2672_out0;
wire v$G3_2977_out0;
wire v$G3_3941_out0;
wire v$G3_3942_out0;
wire v$G3_3950_out0;
wire v$G3_3951_out0;
wire v$G3_4104_out0;
wire v$G3_4105_out0;
wire v$G3_4724_out0;
wire v$G3_4725_out0;
wire v$G3_5001_out0;
wire v$G3_7486_out0;
wire v$G3_7487_out0;
wire v$G3_7488_out0;
wire v$G3_7489_out0;
wire v$G3_7518_out0;
wire v$G3_7519_out0;
wire v$G3_7598_out0;
wire v$G3_7599_out0;
wire v$G3_8040_out0;
wire v$G3_8041_out0;
wire v$G3_8814_out0;
wire v$G3_8815_out0;
wire v$G3_8816_out0;
wire v$G3_8817_out0;
wire v$G3_8818_out0;
wire v$G3_8819_out0;
wire v$G3_8820_out0;
wire v$G3_8821_out0;
wire v$G3_8822_out0;
wire v$G3_8823_out0;
wire v$G3_9357_out0;
wire v$G3_9434_out0;
wire v$G3_9435_out0;
wire v$G3_9940_out0;
wire v$G3_9941_out0;
wire v$G40_13360_out0;
wire v$G40_13361_out0;
wire v$G40_13362_out0;
wire v$G40_13363_out0;
wire v$G40_13364_out0;
wire v$G40_13365_out0;
wire v$G40_13366_out0;
wire v$G40_13367_out0;
wire v$G40_13368_out0;
wire v$G40_13369_out0;
wire v$G40_13370_out0;
wire v$G40_13371_out0;
wire v$G40_13372_out0;
wire v$G40_13373_out0;
wire v$G40_13374_out0;
wire v$G40_13375_out0;
wire v$G40_13376_out0;
wire v$G40_13377_out0;
wire v$G40_13378_out0;
wire v$G40_13379_out0;
wire v$G40_13380_out0;
wire v$G40_13381_out0;
wire v$G40_13382_out0;
wire v$G40_13383_out0;
wire v$G40_13678_out0;
wire v$G40_13679_out0;
wire v$G40_15130_out0;
wire v$G40_15131_out0;
wire v$G41_10872_out0;
wire v$G41_10873_out0;
wire v$G41_10874_out0;
wire v$G41_10875_out0;
wire v$G41_10876_out0;
wire v$G41_10877_out0;
wire v$G41_10878_out0;
wire v$G41_10879_out0;
wire v$G41_10880_out0;
wire v$G41_10881_out0;
wire v$G41_10882_out0;
wire v$G41_10883_out0;
wire v$G41_10884_out0;
wire v$G41_10885_out0;
wire v$G41_10886_out0;
wire v$G41_10887_out0;
wire v$G41_10888_out0;
wire v$G41_10889_out0;
wire v$G41_10890_out0;
wire v$G41_10891_out0;
wire v$G41_10892_out0;
wire v$G41_10893_out0;
wire v$G41_10894_out0;
wire v$G41_10895_out0;
wire v$G41_18479_out0;
wire v$G41_18480_out0;
wire v$G42_18475_out0;
wire v$G42_18476_out0;
wire v$G42_9578_out0;
wire v$G42_9579_out0;
wire v$G43_390_out0;
wire v$G43_391_out0;
wire v$G43_7051_out0;
wire v$G43_7052_out0;
wire v$G44_8251_out0;
wire v$G45_15360_out0;
wire v$G45_16900_out0;
wire v$G45_16901_out0;
wire v$G46_10902_out0;
wire v$G46_10903_out0;
wire v$G46_16116_out0;
wire v$G46_16117_out0;
wire v$G47_1531_out0;
wire v$G47_1532_out0;
wire v$G47_5419_out0;
wire v$G47_5420_out0;
wire v$G48_18516_out0;
wire v$G48_18517_out0;
wire v$G48_2281_out0;
wire v$G48_2282_out0;
wire v$G48_4876_out0;
wire v$G48_4877_out0;
wire v$G49_10451_out0;
wire v$G49_10452_out0;
wire v$G49_11052_out0;
wire v$G49_11053_out0;
wire v$G49_5244_out0;
wire v$G49_5245_out0;
wire v$G4_11111_out0;
wire v$G4_11112_out0;
wire v$G4_11113_out0;
wire v$G4_11114_out0;
wire v$G4_11115_out0;
wire v$G4_11116_out0;
wire v$G4_11117_out0;
wire v$G4_11118_out0;
wire v$G4_11119_out0;
wire v$G4_11120_out0;
wire v$G4_11121_out0;
wire v$G4_11122_out0;
wire v$G4_11123_out0;
wire v$G4_11124_out0;
wire v$G4_11125_out0;
wire v$G4_11126_out0;
wire v$G4_11127_out0;
wire v$G4_11128_out0;
wire v$G4_11129_out0;
wire v$G4_11130_out0;
wire v$G4_11131_out0;
wire v$G4_11132_out0;
wire v$G4_11133_out0;
wire v$G4_11134_out0;
wire v$G4_11135_out0;
wire v$G4_11136_out0;
wire v$G4_11137_out0;
wire v$G4_11138_out0;
wire v$G4_11139_out0;
wire v$G4_11140_out0;
wire v$G4_11141_out0;
wire v$G4_11142_out0;
wire v$G4_11143_out0;
wire v$G4_11144_out0;
wire v$G4_11145_out0;
wire v$G4_11146_out0;
wire v$G4_11147_out0;
wire v$G4_11148_out0;
wire v$G4_11149_out0;
wire v$G4_11150_out0;
wire v$G4_11151_out0;
wire v$G4_11152_out0;
wire v$G4_11153_out0;
wire v$G4_11154_out0;
wire v$G4_11155_out0;
wire v$G4_11156_out0;
wire v$G4_11157_out0;
wire v$G4_11158_out0;
wire v$G4_11159_out0;
wire v$G4_11160_out0;
wire v$G4_11161_out0;
wire v$G4_11162_out0;
wire v$G4_11163_out0;
wire v$G4_11164_out0;
wire v$G4_11165_out0;
wire v$G4_11166_out0;
wire v$G4_11167_out0;
wire v$G4_11168_out0;
wire v$G4_11169_out0;
wire v$G4_11170_out0;
wire v$G4_11171_out0;
wire v$G4_11172_out0;
wire v$G4_11173_out0;
wire v$G4_11174_out0;
wire v$G4_11175_out0;
wire v$G4_11176_out0;
wire v$G4_11177_out0;
wire v$G4_11178_out0;
wire v$G4_11179_out0;
wire v$G4_11180_out0;
wire v$G4_11181_out0;
wire v$G4_11182_out0;
wire v$G4_11183_out0;
wire v$G4_11184_out0;
wire v$G4_11185_out0;
wire v$G4_11186_out0;
wire v$G4_11187_out0;
wire v$G4_11188_out0;
wire v$G4_11189_out0;
wire v$G4_11190_out0;
wire v$G4_11191_out0;
wire v$G4_11192_out0;
wire v$G4_11193_out0;
wire v$G4_11194_out0;
wire v$G4_11195_out0;
wire v$G4_11196_out0;
wire v$G4_11197_out0;
wire v$G4_11198_out0;
wire v$G4_11199_out0;
wire v$G4_11200_out0;
wire v$G4_11201_out0;
wire v$G4_11202_out0;
wire v$G4_11203_out0;
wire v$G4_11204_out0;
wire v$G4_11205_out0;
wire v$G4_11206_out0;
wire v$G4_11207_out0;
wire v$G4_11208_out0;
wire v$G4_11209_out0;
wire v$G4_11210_out0;
wire v$G4_11211_out0;
wire v$G4_11212_out0;
wire v$G4_11213_out0;
wire v$G4_11214_out0;
wire v$G4_11215_out0;
wire v$G4_11216_out0;
wire v$G4_11217_out0;
wire v$G4_11218_out0;
wire v$G4_11219_out0;
wire v$G4_11220_out0;
wire v$G4_11221_out0;
wire v$G4_11222_out0;
wire v$G4_11223_out0;
wire v$G4_11224_out0;
wire v$G4_11225_out0;
wire v$G4_11226_out0;
wire v$G4_11227_out0;
wire v$G4_11228_out0;
wire v$G4_11229_out0;
wire v$G4_11230_out0;
wire v$G4_11231_out0;
wire v$G4_11232_out0;
wire v$G4_11233_out0;
wire v$G4_11234_out0;
wire v$G4_11235_out0;
wire v$G4_11236_out0;
wire v$G4_11237_out0;
wire v$G4_11238_out0;
wire v$G4_11239_out0;
wire v$G4_11240_out0;
wire v$G4_11241_out0;
wire v$G4_11242_out0;
wire v$G4_11243_out0;
wire v$G4_11244_out0;
wire v$G4_11245_out0;
wire v$G4_11246_out0;
wire v$G4_11247_out0;
wire v$G4_11248_out0;
wire v$G4_11249_out0;
wire v$G4_11250_out0;
wire v$G4_11251_out0;
wire v$G4_11252_out0;
wire v$G4_11253_out0;
wire v$G4_11254_out0;
wire v$G4_11255_out0;
wire v$G4_11256_out0;
wire v$G4_11257_out0;
wire v$G4_11258_out0;
wire v$G4_11259_out0;
wire v$G4_11260_out0;
wire v$G4_11261_out0;
wire v$G4_11262_out0;
wire v$G4_11263_out0;
wire v$G4_11264_out0;
wire v$G4_11265_out0;
wire v$G4_11266_out0;
wire v$G4_11267_out0;
wire v$G4_11268_out0;
wire v$G4_11269_out0;
wire v$G4_11270_out0;
wire v$G4_11271_out0;
wire v$G4_11272_out0;
wire v$G4_11273_out0;
wire v$G4_11274_out0;
wire v$G4_11275_out0;
wire v$G4_11276_out0;
wire v$G4_11277_out0;
wire v$G4_11278_out0;
wire v$G4_11279_out0;
wire v$G4_11280_out0;
wire v$G4_11281_out0;
wire v$G4_11282_out0;
wire v$G4_11283_out0;
wire v$G4_11284_out0;
wire v$G4_11285_out0;
wire v$G4_11286_out0;
wire v$G4_11287_out0;
wire v$G4_11288_out0;
wire v$G4_11289_out0;
wire v$G4_11290_out0;
wire v$G4_11291_out0;
wire v$G4_11292_out0;
wire v$G4_11293_out0;
wire v$G4_11294_out0;
wire v$G4_11295_out0;
wire v$G4_11296_out0;
wire v$G4_11297_out0;
wire v$G4_11298_out0;
wire v$G4_11299_out0;
wire v$G4_11300_out0;
wire v$G4_11301_out0;
wire v$G4_11302_out0;
wire v$G4_11303_out0;
wire v$G4_11304_out0;
wire v$G4_11305_out0;
wire v$G4_11306_out0;
wire v$G4_11307_out0;
wire v$G4_11308_out0;
wire v$G4_11309_out0;
wire v$G4_11310_out0;
wire v$G4_11311_out0;
wire v$G4_11312_out0;
wire v$G4_11313_out0;
wire v$G4_11314_out0;
wire v$G4_11315_out0;
wire v$G4_11833_out0;
wire v$G4_11834_out0;
wire v$G4_11835_out0;
wire v$G4_11836_out0;
wire v$G4_11837_out0;
wire v$G4_11838_out0;
wire v$G4_11839_out0;
wire v$G4_11840_out0;
wire v$G4_11841_out0;
wire v$G4_11842_out0;
wire v$G4_11870_out0;
wire v$G4_11871_out0;
wire v$G4_11988_out0;
wire v$G4_11989_out0;
wire v$G4_13187_out0;
wire v$G4_1329_out0;
wire v$G4_1330_out0;
wire v$G4_13999_out0;
wire v$G4_14000_out0;
wire v$G4_14214_out0;
wire v$G4_14215_out0;
wire v$G4_14501_out0;
wire v$G4_14502_out0;
wire v$G4_14683_out0;
wire v$G4_14684_out0;
wire v$G4_15127_out0;
wire v$G4_15128_out0;
wire v$G4_15340_out0;
wire v$G4_15341_out0;
wire v$G4_15457_out0;
wire v$G4_15458_out0;
wire v$G4_15544_out0;
wire v$G4_15545_out0;
wire v$G4_15824_out0;
wire v$G4_15825_out0;
wire v$G4_17523_out0;
wire v$G4_17524_out0;
wire v$G4_17525_out0;
wire v$G4_17526_out0;
wire v$G4_17527_out0;
wire v$G4_17528_out0;
wire v$G4_17529_out0;
wire v$G4_17530_out0;
wire v$G4_17531_out0;
wire v$G4_17532_out0;
wire v$G4_17533_out0;
wire v$G4_17534_out0;
wire v$G4_17535_out0;
wire v$G4_17536_out0;
wire v$G4_17537_out0;
wire v$G4_17538_out0;
wire v$G4_17539_out0;
wire v$G4_17540_out0;
wire v$G4_17541_out0;
wire v$G4_17542_out0;
wire v$G4_17543_out0;
wire v$G4_17544_out0;
wire v$G4_17545_out0;
wire v$G4_17546_out0;
wire v$G4_17547_out0;
wire v$G4_17548_out0;
wire v$G4_17549_out0;
wire v$G4_17550_out0;
wire v$G4_17551_out0;
wire v$G4_17552_out0;
wire v$G4_17553_out0;
wire v$G4_17554_out0;
wire v$G4_17555_out0;
wire v$G4_17556_out0;
wire v$G4_17557_out0;
wire v$G4_17558_out0;
wire v$G4_17559_out0;
wire v$G4_17560_out0;
wire v$G4_17561_out0;
wire v$G4_17562_out0;
wire v$G4_17563_out0;
wire v$G4_17564_out0;
wire v$G4_17565_out0;
wire v$G4_17566_out0;
wire v$G4_17567_out0;
wire v$G4_17568_out0;
wire v$G4_17569_out0;
wire v$G4_17570_out0;
wire v$G4_17586_out0;
wire v$G4_17587_out0;
wire v$G4_18277_out0;
wire v$G4_18278_out0;
wire v$G4_2889_out0;
wire v$G4_2890_out0;
wire v$G4_4029_out0;
wire v$G4_4030_out0;
wire v$G4_4031_out0;
wire v$G4_4032_out0;
wire v$G4_4033_out0;
wire v$G4_4034_out0;
wire v$G4_4035_out0;
wire v$G4_4036_out0;
wire v$G4_4900_out0;
wire v$G4_4901_out0;
wire v$G4_5735_out0;
wire v$G4_5736_out0;
wire v$G4_5737_out0;
wire v$G4_5738_out0;
wire v$G4_5739_out0;
wire v$G4_6053_out0;
wire v$G4_6054_out0;
wire v$G4_6055_out0;
wire v$G4_6056_out0;
wire v$G4_6057_out0;
wire v$G4_6058_out0;
wire v$G4_6059_out0;
wire v$G4_6060_out0;
wire v$G4_6417_out0;
wire v$G4_7548_out0;
wire v$G4_7549_out0;
wire v$G4_7739_out0;
wire v$G4_7740_out0;
wire v$G50_13210_out0;
wire v$G50_13211_out0;
wire v$G50_13303_out0;
wire v$G50_16361_out0;
wire v$G50_16362_out0;
wire v$G50_17323_out0;
wire v$G50_17324_out0;
wire v$G51_14015_out0;
wire v$G51_14016_out0;
wire v$G51_18762_out0;
wire v$G51_2863_out0;
wire v$G51_2864_out0;
wire v$G51_3464_out0;
wire v$G51_3465_out0;
wire v$G52_15938_out0;
wire v$G52_15939_out0;
wire v$G52_2971_out0;
wire v$G52_2972_out0;
wire v$G52_7887_out0;
wire v$G53_12714_out0;
wire v$G53_12715_out0;
wire v$G53_15830_out0;
wire v$G53_15831_out0;
wire v$G53_17493_out0;
wire v$G54_13285_out0;
wire v$G54_14197_out0;
wire v$G54_14198_out0;
wire v$G54_1901_out0;
wire v$G54_1902_out0;
wire v$G54_8133_out0;
wire v$G54_8134_out0;
wire v$G55_13697_out0;
wire v$G55_16658_out0;
wire v$G55_16659_out0;
wire v$G55_18199_out0;
wire v$G55_18200_out0;
wire v$G55_5049_out0;
wire v$G55_5050_out0;
wire v$G56_17676_out0;
wire v$G56_3143_out0;
wire v$G56_3144_out0;
wire v$G56_648_out0;
wire v$G56_649_out0;
wire v$G57_11652_out0;
wire v$G57_11653_out0;
wire v$G57_13452_out0;
wire v$G57_13453_out0;
wire v$G57_17955_out0;
wire v$G57_8978_out0;
wire v$G57_8979_out0;
wire v$G58_168_out0;
wire v$G58_169_out0;
wire v$G58_2518_out0;
wire v$G58_2519_out0;
wire v$G58_7047_out0;
wire v$G58_7048_out0;
wire v$G59_15123_out0;
wire v$G59_15124_out0;
wire v$G59_2571_out0;
wire v$G59_3843_out0;
wire v$G59_3844_out0;
wire v$G5_10676_out0;
wire v$G5_10677_out0;
wire v$G5_10678_out0;
wire v$G5_10679_out0;
wire v$G5_10680_out0;
wire v$G5_10690_out0;
wire v$G5_10691_out0;
wire v$G5_1123_out0;
wire v$G5_1124_out0;
wire v$G5_1125_out0;
wire v$G5_1126_out0;
wire v$G5_1127_out0;
wire v$G5_1128_out0;
wire v$G5_1129_out0;
wire v$G5_1130_out0;
wire v$G5_1131_out0;
wire v$G5_1132_out0;
wire v$G5_12747_out0;
wire v$G5_12748_out0;
wire v$G5_13549_out0;
wire v$G5_13550_out0;
wire v$G5_14649_out0;
wire v$G5_14650_out0;
wire v$G5_14653_out0;
wire v$G5_14654_out0;
wire v$G5_15232_out0;
wire v$G5_15233_out0;
wire v$G5_15791_out0;
wire v$G5_15792_out0;
wire v$G5_16118_out0;
wire v$G5_16119_out0;
wire v$G5_16154_out0;
wire v$G5_16155_out0;
wire v$G5_16556_out0;
wire v$G5_16557_out0;
wire v$G5_17507_out0;
wire v$G5_17508_out0;
wire v$G5_17509_out0;
wire v$G5_17510_out0;
wire v$G5_17511_out0;
wire v$G5_17512_out0;
wire v$G5_17513_out0;
wire v$G5_17514_out0;
wire v$G5_17879_out0;
wire v$G5_17880_out0;
wire v$G5_2235_out0;
wire v$G5_2236_out0;
wire v$G5_2668_out0;
wire v$G5_4519_out0;
wire v$G5_4520_out0;
wire v$G5_4521_out0;
wire v$G5_4522_out0;
wire v$G5_4523_out0;
wire v$G5_4524_out0;
wire v$G5_4525_out0;
wire v$G5_4526_out0;
wire v$G5_4527_out0;
wire v$G5_4528_out0;
wire v$G5_4529_out0;
wire v$G5_4530_out0;
wire v$G5_4531_out0;
wire v$G5_4532_out0;
wire v$G5_4533_out0;
wire v$G5_4534_out0;
wire v$G5_4535_out0;
wire v$G5_4536_out0;
wire v$G5_4537_out0;
wire v$G5_4538_out0;
wire v$G5_4539_out0;
wire v$G5_4540_out0;
wire v$G5_4541_out0;
wire v$G5_4542_out0;
wire v$G5_4543_out0;
wire v$G5_4544_out0;
wire v$G5_4545_out0;
wire v$G5_4546_out0;
wire v$G5_4547_out0;
wire v$G5_4548_out0;
wire v$G5_4549_out0;
wire v$G5_4550_out0;
wire v$G5_4551_out0;
wire v$G5_4552_out0;
wire v$G5_4553_out0;
wire v$G5_4554_out0;
wire v$G5_4555_out0;
wire v$G5_4556_out0;
wire v$G5_4557_out0;
wire v$G5_4558_out0;
wire v$G5_4559_out0;
wire v$G5_4560_out0;
wire v$G5_4561_out0;
wire v$G5_4562_out0;
wire v$G5_4563_out0;
wire v$G5_4564_out0;
wire v$G5_4565_out0;
wire v$G5_4566_out0;
wire v$G5_4567_out0;
wire v$G5_4568_out0;
wire v$G5_4569_out0;
wire v$G5_4570_out0;
wire v$G5_4571_out0;
wire v$G5_4572_out0;
wire v$G5_4573_out0;
wire v$G5_4574_out0;
wire v$G5_4575_out0;
wire v$G5_4576_out0;
wire v$G5_4577_out0;
wire v$G5_4578_out0;
wire v$G5_4579_out0;
wire v$G5_4580_out0;
wire v$G5_4581_out0;
wire v$G5_4582_out0;
wire v$G5_4583_out0;
wire v$G5_4584_out0;
wire v$G5_4585_out0;
wire v$G5_4586_out0;
wire v$G5_4587_out0;
wire v$G5_4588_out0;
wire v$G5_4589_out0;
wire v$G5_4590_out0;
wire v$G5_4591_out0;
wire v$G5_4592_out0;
wire v$G5_4593_out0;
wire v$G5_4594_out0;
wire v$G5_4595_out0;
wire v$G5_4596_out0;
wire v$G5_4597_out0;
wire v$G5_4598_out0;
wire v$G5_4599_out0;
wire v$G5_4600_out0;
wire v$G5_4601_out0;
wire v$G5_4602_out0;
wire v$G5_4603_out0;
wire v$G5_4604_out0;
wire v$G5_4605_out0;
wire v$G5_4606_out0;
wire v$G5_4607_out0;
wire v$G5_4608_out0;
wire v$G5_4609_out0;
wire v$G5_4610_out0;
wire v$G5_4611_out0;
wire v$G5_4612_out0;
wire v$G5_4613_out0;
wire v$G5_4614_out0;
wire v$G5_4615_out0;
wire v$G5_4616_out0;
wire v$G5_4617_out0;
wire v$G5_4618_out0;
wire v$G5_4619_out0;
wire v$G5_4620_out0;
wire v$G5_4621_out0;
wire v$G5_4622_out0;
wire v$G5_4623_out0;
wire v$G5_4624_out0;
wire v$G5_4625_out0;
wire v$G5_4626_out0;
wire v$G5_4627_out0;
wire v$G5_4628_out0;
wire v$G5_4629_out0;
wire v$G5_4630_out0;
wire v$G5_4631_out0;
wire v$G5_4632_out0;
wire v$G5_4633_out0;
wire v$G5_4634_out0;
wire v$G5_4635_out0;
wire v$G5_4636_out0;
wire v$G5_4637_out0;
wire v$G5_4638_out0;
wire v$G5_4639_out0;
wire v$G5_4640_out0;
wire v$G5_4641_out0;
wire v$G5_4642_out0;
wire v$G5_4643_out0;
wire v$G5_4644_out0;
wire v$G5_4645_out0;
wire v$G5_4646_out0;
wire v$G5_4647_out0;
wire v$G5_4648_out0;
wire v$G5_4649_out0;
wire v$G5_4650_out0;
wire v$G5_4651_out0;
wire v$G5_4652_out0;
wire v$G5_4653_out0;
wire v$G5_4654_out0;
wire v$G5_4655_out0;
wire v$G5_4656_out0;
wire v$G5_4657_out0;
wire v$G5_4658_out0;
wire v$G5_4659_out0;
wire v$G5_4660_out0;
wire v$G5_4661_out0;
wire v$G5_4662_out0;
wire v$G5_4663_out0;
wire v$G5_4664_out0;
wire v$G5_4665_out0;
wire v$G5_4666_out0;
wire v$G5_4667_out0;
wire v$G5_4668_out0;
wire v$G5_4669_out0;
wire v$G5_4670_out0;
wire v$G5_4671_out0;
wire v$G5_4672_out0;
wire v$G5_4673_out0;
wire v$G5_4674_out0;
wire v$G5_4675_out0;
wire v$G5_4676_out0;
wire v$G5_4677_out0;
wire v$G5_4678_out0;
wire v$G5_4679_out0;
wire v$G5_4680_out0;
wire v$G5_4681_out0;
wire v$G5_4682_out0;
wire v$G5_4683_out0;
wire v$G5_4684_out0;
wire v$G5_4685_out0;
wire v$G5_4686_out0;
wire v$G5_4687_out0;
wire v$G5_4688_out0;
wire v$G5_4689_out0;
wire v$G5_4690_out0;
wire v$G5_4691_out0;
wire v$G5_4692_out0;
wire v$G5_4693_out0;
wire v$G5_4694_out0;
wire v$G5_4695_out0;
wire v$G5_4696_out0;
wire v$G5_4697_out0;
wire v$G5_4698_out0;
wire v$G5_4699_out0;
wire v$G5_4700_out0;
wire v$G5_4701_out0;
wire v$G5_4702_out0;
wire v$G5_4703_out0;
wire v$G5_4704_out0;
wire v$G5_4705_out0;
wire v$G5_4706_out0;
wire v$G5_4707_out0;
wire v$G5_4708_out0;
wire v$G5_4709_out0;
wire v$G5_4710_out0;
wire v$G5_4711_out0;
wire v$G5_4712_out0;
wire v$G5_4713_out0;
wire v$G5_4714_out0;
wire v$G5_4715_out0;
wire v$G5_4716_out0;
wire v$G5_4717_out0;
wire v$G5_4718_out0;
wire v$G5_4719_out0;
wire v$G5_4720_out0;
wire v$G5_4721_out0;
wire v$G5_4722_out0;
wire v$G5_4723_out0;
wire v$G5_5797_out0;
wire v$G5_5831_out0;
wire v$G5_5832_out0;
wire v$G5_5833_out0;
wire v$G5_5834_out0;
wire v$G5_5835_out0;
wire v$G5_5836_out0;
wire v$G5_5837_out0;
wire v$G5_5838_out0;
wire v$G5_5839_out0;
wire v$G5_5840_out0;
wire v$G5_5841_out0;
wire v$G5_5842_out0;
wire v$G5_5843_out0;
wire v$G5_5844_out0;
wire v$G5_5845_out0;
wire v$G5_5846_out0;
wire v$G5_5847_out0;
wire v$G5_5848_out0;
wire v$G5_5849_out0;
wire v$G5_5850_out0;
wire v$G5_5851_out0;
wire v$G5_5852_out0;
wire v$G5_5853_out0;
wire v$G5_5854_out0;
wire v$G5_5855_out0;
wire v$G5_5856_out0;
wire v$G5_5857_out0;
wire v$G5_5858_out0;
wire v$G5_5859_out0;
wire v$G5_5860_out0;
wire v$G5_5861_out0;
wire v$G5_5862_out0;
wire v$G5_5863_out0;
wire v$G5_5864_out0;
wire v$G5_5865_out0;
wire v$G5_5866_out0;
wire v$G5_5867_out0;
wire v$G5_5868_out0;
wire v$G5_5869_out0;
wire v$G5_5870_out0;
wire v$G5_5871_out0;
wire v$G5_5872_out0;
wire v$G5_5873_out0;
wire v$G5_5874_out0;
wire v$G5_5875_out0;
wire v$G5_5876_out0;
wire v$G5_5877_out0;
wire v$G5_5878_out0;
wire v$G5_6198_out0;
wire v$G5_6199_out0;
wire v$G5_6934_out0;
wire v$G5_6935_out0;
wire v$G5_6936_out0;
wire v$G5_6937_out0;
wire v$G5_6938_out0;
wire v$G5_6939_out0;
wire v$G5_6940_out0;
wire v$G5_6941_out0;
wire v$G5_6942_out0;
wire v$G5_6943_out0;
wire v$G5_6944_out0;
wire v$G5_6945_out0;
wire v$G5_6946_out0;
wire v$G5_6947_out0;
wire v$G5_6948_out0;
wire v$G5_6949_out0;
wire v$G5_6950_out0;
wire v$G5_6951_out0;
wire v$G5_6952_out0;
wire v$G5_6953_out0;
wire v$G5_6954_out0;
wire v$G5_6955_out0;
wire v$G5_6956_out0;
wire v$G5_6957_out0;
wire v$G5_7583_out0;
wire v$G5_7584_out0;
wire v$G5_8448_out0;
wire v$G5_8449_out0;
wire v$G60_18758_out0;
wire v$G60_18759_out0;
wire v$G60_9467_out0;
wire v$G60_9468_out0;
wire v$G61_11603_out0;
wire v$G61_11604_out0;
wire v$G61_16446_out0;
wire v$G61_16447_out0;
wire v$G61_8281_out0;
wire v$G61_8282_out0;
wire v$G62_11755_out0;
wire v$G62_11756_out0;
wire v$G62_11967_out0;
wire v$G62_14987_out0;
wire v$G62_14988_out0;
wire v$G63_10019_out0;
wire v$G63_10020_out0;
wire v$G63_13677_out0;
wire v$G63_16810_out0;
wire v$G63_16811_out0;
wire v$G64_15260_out0;
wire v$G64_15261_out0;
wire v$G64_6395_out0;
wire v$G64_6396_out0;
wire v$G64_6432_out0;
wire v$G64_7783_out0;
wire v$G64_7784_out0;
wire v$G65_14120_out0;
wire v$G65_14121_out0;
wire v$G65_18211_out0;
wire v$G65_18212_out0;
wire v$G65_2460_out0;
wire v$G65_2461_out0;
wire v$G65_8809_out0;
wire v$G66_15270_out0;
wire v$G66_15271_out0;
wire v$G66_16844_out0;
wire v$G66_16845_out0;
wire v$G66_8673_out0;
wire v$G66_8674_out0;
wire v$G66_8931_out0;
wire v$G67_11059_out0;
wire v$G67_11060_out0;
wire v$G67_13755_out0;
wire v$G67_14107_out0;
wire v$G67_14108_out0;
wire v$G68_14822_out0;
wire v$G68_15184_out0;
wire v$G68_15185_out0;
wire v$G68_18108_out0;
wire v$G68_18109_out0;
wire v$G69_1206_out0;
wire v$G69_1207_out0;
wire v$G69_15812_out0;
wire v$G69_8210_out0;
wire v$G69_8211_out0;
wire v$G6_11934_out0;
wire v$G6_11935_out0;
wire v$G6_12126_out0;
wire v$G6_12127_out0;
wire v$G6_13009_out0;
wire v$G6_13010_out0;
wire v$G6_13627_out0;
wire v$G6_13628_out0;
wire v$G6_15559_out0;
wire v$G6_15560_out0;
wire v$G6_15561_out0;
wire v$G6_15562_out0;
wire v$G6_15563_out0;
wire v$G6_15564_out0;
wire v$G6_15565_out0;
wire v$G6_15566_out0;
wire v$G6_15567_out0;
wire v$G6_15568_out0;
wire v$G6_15569_out0;
wire v$G6_15570_out0;
wire v$G6_15571_out0;
wire v$G6_15572_out0;
wire v$G6_15573_out0;
wire v$G6_15574_out0;
wire v$G6_15575_out0;
wire v$G6_15576_out0;
wire v$G6_15577_out0;
wire v$G6_15578_out0;
wire v$G6_15579_out0;
wire v$G6_15580_out0;
wire v$G6_16353_out0;
wire v$G6_16354_out0;
wire v$G6_16355_out0;
wire v$G6_16356_out0;
wire v$G6_16357_out0;
wire v$G6_16809_out0;
wire v$G6_17398_out0;
wire v$G6_2247_out0;
wire v$G6_2248_out0;
wire v$G6_269_out0;
wire v$G6_270_out0;
wire v$G6_3163_out0;
wire v$G6_3164_out0;
wire v$G6_3357_out0;
wire v$G6_3358_out0;
wire v$G6_3503_out0;
wire v$G6_3555_out0;
wire v$G6_3556_out0;
wire v$G6_3557_out0;
wire v$G6_3558_out0;
wire v$G6_3559_out0;
wire v$G6_3560_out0;
wire v$G6_3561_out0;
wire v$G6_3562_out0;
wire v$G6_3563_out0;
wire v$G6_3564_out0;
wire v$G6_3565_out0;
wire v$G6_3566_out0;
wire v$G6_3567_out0;
wire v$G6_3568_out0;
wire v$G6_3569_out0;
wire v$G6_3570_out0;
wire v$G6_3571_out0;
wire v$G6_3572_out0;
wire v$G6_3573_out0;
wire v$G6_3574_out0;
wire v$G6_3575_out0;
wire v$G6_3576_out0;
wire v$G6_3577_out0;
wire v$G6_3578_out0;
wire v$G6_3579_out0;
wire v$G6_3580_out0;
wire v$G6_3581_out0;
wire v$G6_3582_out0;
wire v$G6_3583_out0;
wire v$G6_3584_out0;
wire v$G6_3585_out0;
wire v$G6_3586_out0;
wire v$G6_3587_out0;
wire v$G6_3588_out0;
wire v$G6_3589_out0;
wire v$G6_3590_out0;
wire v$G6_3591_out0;
wire v$G6_3592_out0;
wire v$G6_3593_out0;
wire v$G6_3594_out0;
wire v$G6_3595_out0;
wire v$G6_3596_out0;
wire v$G6_3597_out0;
wire v$G6_3598_out0;
wire v$G6_3599_out0;
wire v$G6_3600_out0;
wire v$G6_3601_out0;
wire v$G6_3602_out0;
wire v$G6_433_out0;
wire v$G6_434_out0;
wire v$G6_435_out0;
wire v$G6_436_out0;
wire v$G6_437_out0;
wire v$G6_438_out0;
wire v$G6_439_out0;
wire v$G6_440_out0;
wire v$G6_441_out0;
wire v$G6_442_out0;
wire v$G6_443_out0;
wire v$G6_444_out0;
wire v$G6_445_out0;
wire v$G6_446_out0;
wire v$G6_447_out0;
wire v$G6_448_out0;
wire v$G6_449_out0;
wire v$G6_450_out0;
wire v$G6_451_out0;
wire v$G6_452_out0;
wire v$G6_453_out0;
wire v$G6_454_out0;
wire v$G6_455_out0;
wire v$G6_456_out0;
wire v$G6_457_out0;
wire v$G6_458_out0;
wire v$G6_459_out0;
wire v$G6_460_out0;
wire v$G6_461_out0;
wire v$G6_462_out0;
wire v$G6_463_out0;
wire v$G6_464_out0;
wire v$G6_465_out0;
wire v$G6_466_out0;
wire v$G6_467_out0;
wire v$G6_468_out0;
wire v$G6_469_out0;
wire v$G6_470_out0;
wire v$G6_471_out0;
wire v$G6_472_out0;
wire v$G6_473_out0;
wire v$G6_474_out0;
wire v$G6_475_out0;
wire v$G6_476_out0;
wire v$G6_477_out0;
wire v$G6_478_out0;
wire v$G6_479_out0;
wire v$G6_480_out0;
wire v$G6_481_out0;
wire v$G6_482_out0;
wire v$G6_483_out0;
wire v$G6_484_out0;
wire v$G6_485_out0;
wire v$G6_486_out0;
wire v$G6_487_out0;
wire v$G6_488_out0;
wire v$G6_489_out0;
wire v$G6_490_out0;
wire v$G6_491_out0;
wire v$G6_492_out0;
wire v$G6_493_out0;
wire v$G6_494_out0;
wire v$G6_495_out0;
wire v$G6_496_out0;
wire v$G6_497_out0;
wire v$G6_498_out0;
wire v$G6_499_out0;
wire v$G6_500_out0;
wire v$G6_501_out0;
wire v$G6_502_out0;
wire v$G6_503_out0;
wire v$G6_504_out0;
wire v$G6_505_out0;
wire v$G6_506_out0;
wire v$G6_507_out0;
wire v$G6_508_out0;
wire v$G6_509_out0;
wire v$G6_510_out0;
wire v$G6_511_out0;
wire v$G6_512_out0;
wire v$G6_513_out0;
wire v$G6_514_out0;
wire v$G6_515_out0;
wire v$G6_516_out0;
wire v$G6_517_out0;
wire v$G6_518_out0;
wire v$G6_519_out0;
wire v$G6_520_out0;
wire v$G6_521_out0;
wire v$G6_522_out0;
wire v$G6_523_out0;
wire v$G6_524_out0;
wire v$G6_525_out0;
wire v$G6_526_out0;
wire v$G6_527_out0;
wire v$G6_528_out0;
wire v$G6_529_out0;
wire v$G6_530_out0;
wire v$G6_531_out0;
wire v$G6_532_out0;
wire v$G6_533_out0;
wire v$G6_534_out0;
wire v$G6_535_out0;
wire v$G6_536_out0;
wire v$G6_537_out0;
wire v$G6_538_out0;
wire v$G6_539_out0;
wire v$G6_540_out0;
wire v$G6_541_out0;
wire v$G6_542_out0;
wire v$G6_543_out0;
wire v$G6_544_out0;
wire v$G6_545_out0;
wire v$G6_5464_out0;
wire v$G6_5465_out0;
wire v$G6_546_out0;
wire v$G6_547_out0;
wire v$G6_548_out0;
wire v$G6_549_out0;
wire v$G6_550_out0;
wire v$G6_551_out0;
wire v$G6_552_out0;
wire v$G6_553_out0;
wire v$G6_554_out0;
wire v$G6_555_out0;
wire v$G6_556_out0;
wire v$G6_557_out0;
wire v$G6_558_out0;
wire v$G6_559_out0;
wire v$G6_560_out0;
wire v$G6_561_out0;
wire v$G6_562_out0;
wire v$G6_563_out0;
wire v$G6_564_out0;
wire v$G6_565_out0;
wire v$G6_566_out0;
wire v$G6_567_out0;
wire v$G6_568_out0;
wire v$G6_569_out0;
wire v$G6_570_out0;
wire v$G6_571_out0;
wire v$G6_572_out0;
wire v$G6_573_out0;
wire v$G6_574_out0;
wire v$G6_575_out0;
wire v$G6_576_out0;
wire v$G6_577_out0;
wire v$G6_578_out0;
wire v$G6_579_out0;
wire v$G6_580_out0;
wire v$G6_581_out0;
wire v$G6_582_out0;
wire v$G6_583_out0;
wire v$G6_584_out0;
wire v$G6_585_out0;
wire v$G6_586_out0;
wire v$G6_587_out0;
wire v$G6_588_out0;
wire v$G6_589_out0;
wire v$G6_590_out0;
wire v$G6_591_out0;
wire v$G6_592_out0;
wire v$G6_593_out0;
wire v$G6_5944_out0;
wire v$G6_5945_out0;
wire v$G6_594_out0;
wire v$G6_595_out0;
wire v$G6_596_out0;
wire v$G6_597_out0;
wire v$G6_598_out0;
wire v$G6_599_out0;
wire v$G6_600_out0;
wire v$G6_601_out0;
wire v$G6_602_out0;
wire v$G6_603_out0;
wire v$G6_604_out0;
wire v$G6_605_out0;
wire v$G6_606_out0;
wire v$G6_607_out0;
wire v$G6_608_out0;
wire v$G6_609_out0;
wire v$G6_610_out0;
wire v$G6_611_out0;
wire v$G6_612_out0;
wire v$G6_613_out0;
wire v$G6_614_out0;
wire v$G6_615_out0;
wire v$G6_6163_out0;
wire v$G6_6164_out0;
wire v$G6_6169_out0;
wire v$G6_616_out0;
wire v$G6_6170_out0;
wire v$G6_6171_out0;
wire v$G6_6172_out0;
wire v$G6_6173_out0;
wire v$G6_6174_out0;
wire v$G6_6175_out0;
wire v$G6_6176_out0;
wire v$G6_6177_out0;
wire v$G6_6178_out0;
wire v$G6_6179_out0;
wire v$G6_617_out0;
wire v$G6_6180_out0;
wire v$G6_618_out0;
wire v$G6_619_out0;
wire v$G6_620_out0;
wire v$G6_621_out0;
wire v$G6_622_out0;
wire v$G6_623_out0;
wire v$G6_624_out0;
wire v$G6_625_out0;
wire v$G6_626_out0;
wire v$G6_627_out0;
wire v$G6_628_out0;
wire v$G6_629_out0;
wire v$G6_630_out0;
wire v$G6_631_out0;
wire v$G6_632_out0;
wire v$G6_633_out0;
wire v$G6_634_out0;
wire v$G6_635_out0;
wire v$G6_636_out0;
wire v$G6_637_out0;
wire v$G6_6549_out0;
wire v$G6_6550_out0;
wire v$G6_6551_out0;
wire v$G6_6552_out0;
wire v$G6_6553_out0;
wire v$G6_6554_out0;
wire v$G6_6555_out0;
wire v$G6_6556_out0;
wire v$G6_6557_out0;
wire v$G6_6558_out0;
wire v$G6_6559_out0;
wire v$G6_6560_out0;
wire v$G6_6561_out0;
wire v$G6_6562_out0;
wire v$G6_6563_out0;
wire v$G6_6564_out0;
wire v$G6_6565_out0;
wire v$G6_6566_out0;
wire v$G6_6567_out0;
wire v$G6_6568_out0;
wire v$G6_6569_out0;
wire v$G6_6570_out0;
wire v$G6_6571_out0;
wire v$G6_6572_out0;
wire v$G6_668_out0;
wire v$G6_669_out0;
wire v$G6_7480_out0;
wire v$G6_7481_out0;
wire v$G6_7939_out0;
wire v$G6_7940_out0;
wire v$G6_9076_out0;
wire v$G6_9077_out0;
wire v$G70_10280_out0;
wire v$G70_10281_out0;
wire v$G70_14028_out0;
wire v$G71_15274_out0;
wire v$G71_15275_out0;
wire v$G72_5901_out0;
wire v$G74_15740_out0;
wire v$G77_18210_out0;
wire v$G78_7096_out0;
wire v$G79_12737_out0;
wire v$G7_10967_out0;
wire v$G7_10968_out0;
wire v$G7_11796_out0;
wire v$G7_11797_out0;
wire v$G7_12203_out0;
wire v$G7_12204_out0;
wire v$G7_12647_out0;
wire v$G7_12648_out0;
wire v$G7_13431_out0;
wire v$G7_13432_out0;
wire v$G7_13559_out0;
wire v$G7_13560_out0;
wire v$G7_14122_out0;
wire v$G7_14123_out0;
wire v$G7_14124_out0;
wire v$G7_14125_out0;
wire v$G7_14126_out0;
wire v$G7_14127_out0;
wire v$G7_14128_out0;
wire v$G7_14129_out0;
wire v$G7_14130_out0;
wire v$G7_14131_out0;
wire v$G7_14132_out0;
wire v$G7_14133_out0;
wire v$G7_14311_out0;
wire v$G7_14312_out0;
wire v$G7_14673_out0;
wire v$G7_14674_out0;
wire v$G7_14806_out0;
wire v$G7_1498_out0;
wire v$G7_1499_out0;
wire v$G7_1691_out0;
wire v$G7_1692_out0;
wire v$G7_1693_out0;
wire v$G7_1694_out0;
wire v$G7_1695_out0;
wire v$G7_17665_out0;
wire v$G7_18131_out0;
wire v$G7_18132_out0;
wire v$G7_18133_out0;
wire v$G7_18134_out0;
wire v$G7_18135_out0;
wire v$G7_18136_out0;
wire v$G7_18137_out0;
wire v$G7_18138_out0;
wire v$G7_18139_out0;
wire v$G7_18140_out0;
wire v$G7_18141_out0;
wire v$G7_18142_out0;
wire v$G7_18143_out0;
wire v$G7_18144_out0;
wire v$G7_18145_out0;
wire v$G7_18146_out0;
wire v$G7_18147_out0;
wire v$G7_18148_out0;
wire v$G7_18149_out0;
wire v$G7_18150_out0;
wire v$G7_18151_out0;
wire v$G7_18152_out0;
wire v$G7_18153_out0;
wire v$G7_18154_out0;
wire v$G7_18155_out0;
wire v$G7_18156_out0;
wire v$G7_18157_out0;
wire v$G7_18158_out0;
wire v$G7_18159_out0;
wire v$G7_18160_out0;
wire v$G7_18161_out0;
wire v$G7_18162_out0;
wire v$G7_18163_out0;
wire v$G7_18164_out0;
wire v$G7_18165_out0;
wire v$G7_18166_out0;
wire v$G7_18167_out0;
wire v$G7_18168_out0;
wire v$G7_18169_out0;
wire v$G7_18170_out0;
wire v$G7_18171_out0;
wire v$G7_18172_out0;
wire v$G7_18173_out0;
wire v$G7_18174_out0;
wire v$G7_18175_out0;
wire v$G7_18176_out0;
wire v$G7_18177_out0;
wire v$G7_18178_out0;
wire v$G7_1831_out0;
wire v$G7_1832_out0;
wire v$G7_18641_out0;
wire v$G7_18642_out0;
wire v$G7_2237_out0;
wire v$G7_2238_out0;
wire v$G7_2239_out0;
wire v$G7_2240_out0;
wire v$G7_3159_out0;
wire v$G7_3160_out0;
wire v$G7_7726_out0;
wire v$G7_7727_out0;
wire v$G7_7846_out0;
wire v$G7_7847_out0;
wire v$G7_9635_out0;
wire v$G7_9636_out0;
wire v$G7_9637_out0;
wire v$G7_9638_out0;
wire v$G7_9639_out0;
wire v$G7_9640_out0;
wire v$G7_9641_out0;
wire v$G7_9642_out0;
wire v$G7_9643_out0;
wire v$G7_9644_out0;
wire v$G7_9645_out0;
wire v$G7_9646_out0;
wire v$G7_9647_out0;
wire v$G7_9648_out0;
wire v$G7_9649_out0;
wire v$G7_9650_out0;
wire v$G7_9651_out0;
wire v$G7_9652_out0;
wire v$G7_9653_out0;
wire v$G7_9654_out0;
wire v$G7_9655_out0;
wire v$G7_9656_out0;
wire v$G7_9657_out0;
wire v$G7_9658_out0;
wire v$G7_9659_out0;
wire v$G7_9660_out0;
wire v$G7_9661_out0;
wire v$G7_9662_out0;
wire v$G7_9663_out0;
wire v$G7_9664_out0;
wire v$G7_9665_out0;
wire v$G7_9666_out0;
wire v$G7_9667_out0;
wire v$G7_9668_out0;
wire v$G7_9669_out0;
wire v$G7_9670_out0;
wire v$G7_9671_out0;
wire v$G7_9672_out0;
wire v$G7_9673_out0;
wire v$G7_9674_out0;
wire v$G7_9675_out0;
wire v$G7_9676_out0;
wire v$G7_9677_out0;
wire v$G7_9678_out0;
wire v$G7_9679_out0;
wire v$G7_9680_out0;
wire v$G7_9681_out0;
wire v$G7_9682_out0;
wire v$G7_9683_out0;
wire v$G7_9684_out0;
wire v$G7_9685_out0;
wire v$G7_9686_out0;
wire v$G7_9687_out0;
wire v$G7_9688_out0;
wire v$G7_9689_out0;
wire v$G7_9690_out0;
wire v$G7_9691_out0;
wire v$G7_9692_out0;
wire v$G7_9693_out0;
wire v$G7_9694_out0;
wire v$G7_9695_out0;
wire v$G7_9696_out0;
wire v$G7_9697_out0;
wire v$G7_9698_out0;
wire v$G7_9699_out0;
wire v$G7_9700_out0;
wire v$G7_9701_out0;
wire v$G7_9702_out0;
wire v$G7_9703_out0;
wire v$G7_9704_out0;
wire v$G7_9705_out0;
wire v$G7_9706_out0;
wire v$G7_9707_out0;
wire v$G7_9708_out0;
wire v$G7_9709_out0;
wire v$G7_9710_out0;
wire v$G7_9711_out0;
wire v$G7_9712_out0;
wire v$G7_9713_out0;
wire v$G7_9714_out0;
wire v$G7_9715_out0;
wire v$G7_9716_out0;
wire v$G7_9717_out0;
wire v$G7_9718_out0;
wire v$G7_9719_out0;
wire v$G7_9720_out0;
wire v$G7_9721_out0;
wire v$G7_9722_out0;
wire v$G7_9723_out0;
wire v$G7_9724_out0;
wire v$G7_9725_out0;
wire v$G7_9726_out0;
wire v$G7_9727_out0;
wire v$G7_9728_out0;
wire v$G7_9729_out0;
wire v$G7_9730_out0;
wire v$G7_9731_out0;
wire v$G7_9732_out0;
wire v$G7_9733_out0;
wire v$G7_9734_out0;
wire v$G7_9735_out0;
wire v$G7_9736_out0;
wire v$G7_9737_out0;
wire v$G7_9738_out0;
wire v$G7_9739_out0;
wire v$G7_9740_out0;
wire v$G7_9741_out0;
wire v$G7_9742_out0;
wire v$G7_9743_out0;
wire v$G7_9744_out0;
wire v$G7_9745_out0;
wire v$G7_9746_out0;
wire v$G7_9747_out0;
wire v$G7_9748_out0;
wire v$G7_9749_out0;
wire v$G7_9750_out0;
wire v$G7_9751_out0;
wire v$G7_9752_out0;
wire v$G7_9753_out0;
wire v$G7_9754_out0;
wire v$G7_9755_out0;
wire v$G7_9756_out0;
wire v$G7_9757_out0;
wire v$G7_9758_out0;
wire v$G7_9759_out0;
wire v$G7_9760_out0;
wire v$G7_9761_out0;
wire v$G7_9762_out0;
wire v$G7_9763_out0;
wire v$G7_9764_out0;
wire v$G7_9765_out0;
wire v$G7_9766_out0;
wire v$G7_9767_out0;
wire v$G7_9768_out0;
wire v$G7_9769_out0;
wire v$G7_9770_out0;
wire v$G7_9771_out0;
wire v$G7_9772_out0;
wire v$G7_9773_out0;
wire v$G7_9774_out0;
wire v$G7_9775_out0;
wire v$G7_9776_out0;
wire v$G7_9777_out0;
wire v$G7_9778_out0;
wire v$G7_9779_out0;
wire v$G7_9780_out0;
wire v$G7_9781_out0;
wire v$G7_9782_out0;
wire v$G7_9783_out0;
wire v$G7_9784_out0;
wire v$G7_9785_out0;
wire v$G7_9786_out0;
wire v$G7_9787_out0;
wire v$G7_9788_out0;
wire v$G7_9789_out0;
wire v$G7_9790_out0;
wire v$G7_9791_out0;
wire v$G7_9792_out0;
wire v$G7_9793_out0;
wire v$G7_9794_out0;
wire v$G7_9795_out0;
wire v$G7_9796_out0;
wire v$G7_9797_out0;
wire v$G7_9798_out0;
wire v$G7_9799_out0;
wire v$G7_9800_out0;
wire v$G7_9801_out0;
wire v$G7_9802_out0;
wire v$G7_9803_out0;
wire v$G7_9804_out0;
wire v$G7_9805_out0;
wire v$G7_9806_out0;
wire v$G7_9807_out0;
wire v$G7_9808_out0;
wire v$G7_9809_out0;
wire v$G7_9810_out0;
wire v$G7_9811_out0;
wire v$G7_9812_out0;
wire v$G7_9813_out0;
wire v$G7_9814_out0;
wire v$G7_9815_out0;
wire v$G7_9816_out0;
wire v$G7_9817_out0;
wire v$G7_9818_out0;
wire v$G7_9819_out0;
wire v$G7_9820_out0;
wire v$G7_9821_out0;
wire v$G7_9822_out0;
wire v$G7_9823_out0;
wire v$G7_9824_out0;
wire v$G7_9825_out0;
wire v$G7_9826_out0;
wire v$G7_9827_out0;
wire v$G7_9828_out0;
wire v$G7_9829_out0;
wire v$G7_9830_out0;
wire v$G7_9831_out0;
wire v$G7_9832_out0;
wire v$G7_9833_out0;
wire v$G7_9834_out0;
wire v$G7_9835_out0;
wire v$G7_9836_out0;
wire v$G7_9837_out0;
wire v$G7_9838_out0;
wire v$G7_9839_out0;
wire v$G7_9851_out0;
wire v$G7_9852_out0;
wire v$G7_9853_out0;
wire v$G7_9854_out0;
wire v$G7_9855_out0;
wire v$G7_9856_out0;
wire v$G7_9857_out0;
wire v$G7_9858_out0;
wire v$G7_9859_out0;
wire v$G7_9860_out0;
wire v$G7_9875_out0;
wire v$G7_9938_out0;
wire v$G7_9939_out0;
wire v$G83_428_out0;
wire v$G84_1235_out0;
wire v$G85_6200_out0;
wire v$G86_13527_out0;
wire v$G87_5144_out0;
wire v$G88_7401_out0;
wire v$G89_17772_out0;
wire v$G8_11068_out0;
wire v$G8_11069_out0;
wire v$G8_11395_out0;
wire v$G8_11396_out0;
wire v$G8_11397_out0;
wire v$G8_11398_out0;
wire v$G8_11399_out0;
wire v$G8_11400_out0;
wire v$G8_11401_out0;
wire v$G8_11402_out0;
wire v$G8_11403_out0;
wire v$G8_11404_out0;
wire v$G8_11405_out0;
wire v$G8_11406_out0;
wire v$G8_11407_out0;
wire v$G8_11408_out0;
wire v$G8_11409_out0;
wire v$G8_11410_out0;
wire v$G8_11411_out0;
wire v$G8_11412_out0;
wire v$G8_11413_out0;
wire v$G8_11414_out0;
wire v$G8_11415_out0;
wire v$G8_11416_out0;
wire v$G8_11417_out0;
wire v$G8_11418_out0;
wire v$G8_11419_out0;
wire v$G8_11420_out0;
wire v$G8_11421_out0;
wire v$G8_11422_out0;
wire v$G8_11423_out0;
wire v$G8_11424_out0;
wire v$G8_11425_out0;
wire v$G8_11426_out0;
wire v$G8_11427_out0;
wire v$G8_11428_out0;
wire v$G8_11429_out0;
wire v$G8_11430_out0;
wire v$G8_11431_out0;
wire v$G8_11432_out0;
wire v$G8_11433_out0;
wire v$G8_11434_out0;
wire v$G8_11435_out0;
wire v$G8_11436_out0;
wire v$G8_11437_out0;
wire v$G8_11438_out0;
wire v$G8_11439_out0;
wire v$G8_11440_out0;
wire v$G8_11441_out0;
wire v$G8_11442_out0;
wire v$G8_11443_out0;
wire v$G8_11444_out0;
wire v$G8_11445_out0;
wire v$G8_11446_out0;
wire v$G8_11447_out0;
wire v$G8_11448_out0;
wire v$G8_11449_out0;
wire v$G8_11450_out0;
wire v$G8_11451_out0;
wire v$G8_11452_out0;
wire v$G8_11453_out0;
wire v$G8_11454_out0;
wire v$G8_11455_out0;
wire v$G8_11456_out0;
wire v$G8_11457_out0;
wire v$G8_11458_out0;
wire v$G8_11459_out0;
wire v$G8_11460_out0;
wire v$G8_11461_out0;
wire v$G8_11462_out0;
wire v$G8_11463_out0;
wire v$G8_11464_out0;
wire v$G8_11465_out0;
wire v$G8_11466_out0;
wire v$G8_11467_out0;
wire v$G8_11468_out0;
wire v$G8_11469_out0;
wire v$G8_11470_out0;
wire v$G8_11471_out0;
wire v$G8_11472_out0;
wire v$G8_11473_out0;
wire v$G8_11474_out0;
wire v$G8_11475_out0;
wire v$G8_11476_out0;
wire v$G8_11477_out0;
wire v$G8_11478_out0;
wire v$G8_11479_out0;
wire v$G8_11480_out0;
wire v$G8_11481_out0;
wire v$G8_11482_out0;
wire v$G8_11483_out0;
wire v$G8_11484_out0;
wire v$G8_11485_out0;
wire v$G8_11486_out0;
wire v$G8_11487_out0;
wire v$G8_11488_out0;
wire v$G8_11489_out0;
wire v$G8_11490_out0;
wire v$G8_11491_out0;
wire v$G8_11492_out0;
wire v$G8_11493_out0;
wire v$G8_11494_out0;
wire v$G8_11495_out0;
wire v$G8_11496_out0;
wire v$G8_11497_out0;
wire v$G8_11498_out0;
wire v$G8_11499_out0;
wire v$G8_11500_out0;
wire v$G8_11501_out0;
wire v$G8_11502_out0;
wire v$G8_11503_out0;
wire v$G8_11504_out0;
wire v$G8_11505_out0;
wire v$G8_11506_out0;
wire v$G8_11507_out0;
wire v$G8_11508_out0;
wire v$G8_11509_out0;
wire v$G8_11510_out0;
wire v$G8_11511_out0;
wire v$G8_11512_out0;
wire v$G8_11513_out0;
wire v$G8_11514_out0;
wire v$G8_11515_out0;
wire v$G8_11516_out0;
wire v$G8_11517_out0;
wire v$G8_11518_out0;
wire v$G8_11519_out0;
wire v$G8_11520_out0;
wire v$G8_11521_out0;
wire v$G8_11522_out0;
wire v$G8_11523_out0;
wire v$G8_11524_out0;
wire v$G8_11525_out0;
wire v$G8_11526_out0;
wire v$G8_11527_out0;
wire v$G8_11528_out0;
wire v$G8_11529_out0;
wire v$G8_11530_out0;
wire v$G8_11531_out0;
wire v$G8_11532_out0;
wire v$G8_11533_out0;
wire v$G8_11534_out0;
wire v$G8_11535_out0;
wire v$G8_11536_out0;
wire v$G8_11537_out0;
wire v$G8_11538_out0;
wire v$G8_11539_out0;
wire v$G8_11540_out0;
wire v$G8_11541_out0;
wire v$G8_11542_out0;
wire v$G8_11543_out0;
wire v$G8_11544_out0;
wire v$G8_11545_out0;
wire v$G8_11546_out0;
wire v$G8_11547_out0;
wire v$G8_11548_out0;
wire v$G8_11549_out0;
wire v$G8_11550_out0;
wire v$G8_11551_out0;
wire v$G8_11552_out0;
wire v$G8_11553_out0;
wire v$G8_11554_out0;
wire v$G8_11555_out0;
wire v$G8_11556_out0;
wire v$G8_11557_out0;
wire v$G8_11558_out0;
wire v$G8_11559_out0;
wire v$G8_11560_out0;
wire v$G8_11561_out0;
wire v$G8_11562_out0;
wire v$G8_11563_out0;
wire v$G8_11564_out0;
wire v$G8_11565_out0;
wire v$G8_11566_out0;
wire v$G8_11567_out0;
wire v$G8_11568_out0;
wire v$G8_11569_out0;
wire v$G8_11570_out0;
wire v$G8_11571_out0;
wire v$G8_11572_out0;
wire v$G8_11573_out0;
wire v$G8_11574_out0;
wire v$G8_11575_out0;
wire v$G8_11576_out0;
wire v$G8_11577_out0;
wire v$G8_11578_out0;
wire v$G8_11579_out0;
wire v$G8_11580_out0;
wire v$G8_11581_out0;
wire v$G8_11582_out0;
wire v$G8_11583_out0;
wire v$G8_11584_out0;
wire v$G8_11585_out0;
wire v$G8_11586_out0;
wire v$G8_11587_out0;
wire v$G8_11588_out0;
wire v$G8_11589_out0;
wire v$G8_11590_out0;
wire v$G8_11591_out0;
wire v$G8_11592_out0;
wire v$G8_11593_out0;
wire v$G8_11594_out0;
wire v$G8_11595_out0;
wire v$G8_11596_out0;
wire v$G8_11597_out0;
wire v$G8_11598_out0;
wire v$G8_11599_out0;
wire v$G8_11990_out0;
wire v$G8_11991_out0;
wire v$G8_11992_out0;
wire v$G8_11993_out0;
wire v$G8_11994_out0;
wire v$G8_11995_out0;
wire v$G8_11996_out0;
wire v$G8_11997_out0;
wire v$G8_11998_out0;
wire v$G8_11999_out0;
wire v$G8_12000_out0;
wire v$G8_12001_out0;
wire v$G8_12002_out0;
wire v$G8_12003_out0;
wire v$G8_12004_out0;
wire v$G8_12005_out0;
wire v$G8_12006_out0;
wire v$G8_12007_out0;
wire v$G8_12008_out0;
wire v$G8_12009_out0;
wire v$G8_12010_out0;
wire v$G8_12011_out0;
wire v$G8_12012_out0;
wire v$G8_12013_out0;
wire v$G8_12014_out0;
wire v$G8_12015_out0;
wire v$G8_12016_out0;
wire v$G8_12017_out0;
wire v$G8_12018_out0;
wire v$G8_12019_out0;
wire v$G8_12020_out0;
wire v$G8_12021_out0;
wire v$G8_12022_out0;
wire v$G8_12023_out0;
wire v$G8_12024_out0;
wire v$G8_12025_out0;
wire v$G8_12026_out0;
wire v$G8_12027_out0;
wire v$G8_12028_out0;
wire v$G8_12029_out0;
wire v$G8_12030_out0;
wire v$G8_12031_out0;
wire v$G8_12032_out0;
wire v$G8_12033_out0;
wire v$G8_12034_out0;
wire v$G8_12035_out0;
wire v$G8_12036_out0;
wire v$G8_12037_out0;
wire v$G8_12296_out0;
wire v$G8_12297_out0;
wire v$G8_1247_out0;
wire v$G8_12482_out0;
wire v$G8_12483_out0;
wire v$G8_1248_out0;
wire v$G8_13403_out0;
wire v$G8_13404_out0;
wire v$G8_14256_out0;
wire v$G8_14257_out0;
wire v$G8_14258_out0;
wire v$G8_14259_out0;
wire v$G8_14260_out0;
wire v$G8_14261_out0;
wire v$G8_14262_out0;
wire v$G8_14263_out0;
wire v$G8_14264_out0;
wire v$G8_14265_out0;
wire v$G8_14266_out0;
wire v$G8_14267_out0;
wire v$G8_15479_out0;
wire v$G8_15480_out0;
wire v$G8_15731_out0;
wire v$G8_17897_out0;
wire v$G8_17898_out0;
wire v$G8_18779_out0;
wire v$G8_18780_out0;
wire v$G8_1886_out0;
wire v$G8_1887_out0;
wire v$G8_1888_out0;
wire v$G8_1889_out0;
wire v$G8_1890_out0;
wire v$G8_1891_out0;
wire v$G8_1892_out0;
wire v$G8_1893_out0;
wire v$G8_2243_out0;
wire v$G8_2244_out0;
wire v$G8_2267_out0;
wire v$G8_2268_out0;
wire v$G8_2414_out0;
wire v$G8_2415_out0;
wire v$G8_246_out0;
wire v$G8_247_out0;
wire v$G8_2577_out0;
wire v$G8_2578_out0;
wire v$G8_2579_out0;
wire v$G8_2580_out0;
wire v$G8_2581_out0;
wire v$G8_3726_out0;
wire v$G8_3727_out0;
wire v$G8_3728_out0;
wire v$G8_3729_out0;
wire v$G8_3730_out0;
wire v$G8_3731_out0;
wire v$G8_3732_out0;
wire v$G8_3733_out0;
wire v$G8_3734_out0;
wire v$G8_3735_out0;
wire v$G8_3736_out0;
wire v$G8_3737_out0;
wire v$G8_3738_out0;
wire v$G8_3739_out0;
wire v$G8_3740_out0;
wire v$G8_3741_out0;
wire v$G8_3742_out0;
wire v$G8_3743_out0;
wire v$G8_3744_out0;
wire v$G8_3745_out0;
wire v$G8_3746_out0;
wire v$G8_3747_out0;
wire v$G8_3748_out0;
wire v$G8_3749_out0;
wire v$G8_4819_out0;
wire v$G8_4820_out0;
wire v$G8_6047_out0;
wire v$G8_6048_out0;
wire v$G8_6064_out0;
wire v$G8_6065_out0;
wire v$G8_9083_out0;
wire v$G8_9084_out0;
wire v$G8_9504_out0;
wire v$G8_9505_out0;
wire v$G90_8054_out0;
wire v$G9_1184_out0;
wire v$G9_1185_out0;
wire v$G9_13446_out0;
wire v$G9_13447_out0;
wire v$G9_15125_out0;
wire v$G9_15126_out0;
wire v$G9_15198_out0;
wire v$G9_15199_out0;
wire v$G9_15200_out0;
wire v$G9_15201_out0;
wire v$G9_15202_out0;
wire v$G9_15203_out0;
wire v$G9_15204_out0;
wire v$G9_15205_out0;
wire v$G9_15206_out0;
wire v$G9_15207_out0;
wire v$G9_15208_out0;
wire v$G9_15209_out0;
wire v$G9_15531_out0;
wire v$G9_15532_out0;
wire v$G9_15590_out0;
wire v$G9_15591_out0;
wire v$G9_16037_out0;
wire v$G9_16038_out0;
wire v$G9_16494_out0;
wire v$G9_16495_out0;
wire v$G9_16920_out0;
wire v$G9_16921_out0;
wire v$G9_16963_out0;
wire v$G9_16964_out0;
wire v$G9_17008_out0;
wire v$G9_17009_out0;
wire v$G9_17588_out0;
wire v$G9_17589_out0;
wire v$G9_17590_out0;
wire v$G9_17591_out0;
wire v$G9_17592_out0;
wire v$G9_17593_out0;
wire v$G9_17594_out0;
wire v$G9_17595_out0;
wire v$G9_17596_out0;
wire v$G9_17597_out0;
wire v$G9_17598_out0;
wire v$G9_17599_out0;
wire v$G9_17600_out0;
wire v$G9_17601_out0;
wire v$G9_17602_out0;
wire v$G9_17603_out0;
wire v$G9_17604_out0;
wire v$G9_17605_out0;
wire v$G9_17606_out0;
wire v$G9_17607_out0;
wire v$G9_17608_out0;
wire v$G9_17609_out0;
wire v$G9_17610_out0;
wire v$G9_17611_out0;
wire v$G9_17612_out0;
wire v$G9_17613_out0;
wire v$G9_17614_out0;
wire v$G9_17615_out0;
wire v$G9_17616_out0;
wire v$G9_17617_out0;
wire v$G9_17618_out0;
wire v$G9_17619_out0;
wire v$G9_17620_out0;
wire v$G9_17621_out0;
wire v$G9_17622_out0;
wire v$G9_17623_out0;
wire v$G9_17624_out0;
wire v$G9_17625_out0;
wire v$G9_17626_out0;
wire v$G9_17627_out0;
wire v$G9_17628_out0;
wire v$G9_17629_out0;
wire v$G9_17630_out0;
wire v$G9_17631_out0;
wire v$G9_17632_out0;
wire v$G9_17633_out0;
wire v$G9_17634_out0;
wire v$G9_17635_out0;
wire v$G9_17710_out0;
wire v$G9_17711_out0;
wire v$G9_2527_out0;
wire v$G9_2528_out0;
wire v$G9_3441_out0;
wire v$G9_3442_out0;
wire v$G9_5798_out0;
wire v$G9_5799_out0;
wire v$G9_6226_out0;
wire v$G9_6227_out0;
wire v$G9_6337_out0;
wire v$G9_6338_out0;
wire v$G9_8671_out0;
wire v$G9_8672_out0;
wire v$G9_8925_out0;
wire v$G9_8926_out0;
wire v$G9_8927_out0;
wire v$G9_8928_out0;
wire v$G9_8929_out0;
wire v$GATE1_659_out0;
wire v$GATE1_660_out0;
wire v$GATE1_661_out0;
wire v$GATE1_662_out0;
wire v$GATE1_663_out0;
wire v$GATE2_15756_out0;
wire v$GATE2_15757_out0;
wire v$GATE2_15758_out0;
wire v$GATE2_15759_out0;
wire v$GATE2_15760_out0;
wire v$G_10055_out0;
wire v$G_10056_out0;
wire v$G_10057_out0;
wire v$G_10058_out0;
wire v$G_10059_out0;
wire v$G_10060_out0;
wire v$G_10061_out0;
wire v$G_10062_out0;
wire v$G_10063_out0;
wire v$G_10064_out0;
wire v$G_10065_out0;
wire v$G_10066_out0;
wire v$G_10067_out0;
wire v$G_10068_out0;
wire v$G_10069_out0;
wire v$G_10070_out0;
wire v$G_10071_out0;
wire v$G_10072_out0;
wire v$G_10073_out0;
wire v$G_10074_out0;
wire v$G_10075_out0;
wire v$G_10076_out0;
wire v$G_10077_out0;
wire v$G_10078_out0;
wire v$G_10079_out0;
wire v$G_10080_out0;
wire v$G_10081_out0;
wire v$G_10082_out0;
wire v$G_10083_out0;
wire v$G_10084_out0;
wire v$G_10085_out0;
wire v$G_10086_out0;
wire v$G_10087_out0;
wire v$G_10088_out0;
wire v$G_10089_out0;
wire v$G_10090_out0;
wire v$G_10091_out0;
wire v$G_10092_out0;
wire v$G_10093_out0;
wire v$G_10094_out0;
wire v$G_10095_out0;
wire v$G_10096_out0;
wire v$G_10097_out0;
wire v$G_10098_out0;
wire v$G_10099_out0;
wire v$G_10100_out0;
wire v$G_10101_out0;
wire v$G_10102_out0;
wire v$G_10103_out0;
wire v$G_10104_out0;
wire v$G_10105_out0;
wire v$G_10106_out0;
wire v$G_10107_out0;
wire v$G_10108_out0;
wire v$G_10109_out0;
wire v$G_10110_out0;
wire v$G_10111_out0;
wire v$G_10112_out0;
wire v$G_10113_out0;
wire v$G_10114_out0;
wire v$G_10115_out0;
wire v$G_10116_out0;
wire v$G_10117_out0;
wire v$G_10118_out0;
wire v$G_10119_out0;
wire v$G_10120_out0;
wire v$G_10121_out0;
wire v$G_10122_out0;
wire v$G_10123_out0;
wire v$G_10124_out0;
wire v$G_10125_out0;
wire v$G_10126_out0;
wire v$G_10127_out0;
wire v$G_10128_out0;
wire v$G_10129_out0;
wire v$G_10130_out0;
wire v$G_10131_out0;
wire v$G_10132_out0;
wire v$G_10133_out0;
wire v$G_10134_out0;
wire v$G_10135_out0;
wire v$G_10136_out0;
wire v$G_10137_out0;
wire v$G_10138_out0;
wire v$G_10139_out0;
wire v$G_10140_out0;
wire v$G_10141_out0;
wire v$G_10142_out0;
wire v$G_10143_out0;
wire v$G_10144_out0;
wire v$G_10145_out0;
wire v$G_10146_out0;
wire v$G_10147_out0;
wire v$G_10148_out0;
wire v$G_10149_out0;
wire v$G_10150_out0;
wire v$G_10151_out0;
wire v$G_10152_out0;
wire v$G_10153_out0;
wire v$G_10154_out0;
wire v$G_10155_out0;
wire v$G_10156_out0;
wire v$G_10157_out0;
wire v$G_10158_out0;
wire v$G_10159_out0;
wire v$G_10160_out0;
wire v$G_10161_out0;
wire v$G_10162_out0;
wire v$G_10163_out0;
wire v$G_10164_out0;
wire v$G_10165_out0;
wire v$G_10166_out0;
wire v$G_10167_out0;
wire v$G_10168_out0;
wire v$G_10169_out0;
wire v$G_10170_out0;
wire v$G_10171_out0;
wire v$G_10172_out0;
wire v$G_10173_out0;
wire v$G_10174_out0;
wire v$HALT$PREV$PREV$PREV_7732_out0;
wire v$HALT$PREV$PREV$PREV_7733_out0;
wire v$HALT$PREV$PREV_18074_out0;
wire v$HALT$PREV$PREV_18075_out0;
wire v$HALT$PREV_10386_out0;
wire v$HALT$PREV_10387_out0;
wire v$HALT0_11685_out0;
wire v$HALT0_14137_out0;
wire v$HALT0_361_out0;
wire v$HALT0_5804_out0;
wire v$HALT1_18308_out0;
wire v$HALT1_3104_out0;
wire v$HALT1_4159_out0;
wire v$HALT1_7229_out0;
wire v$HALTED_11827_out0;
wire v$HALTED_11828_out0;
wire v$HALTSEL_14742_out0;
wire v$HALTVALID_13286_out0;
wire v$HALTVALID_7744_out0;
wire v$HALT_12900_out0;
wire v$HALT_12901_out0;
wire v$HALT_1290_out0;
wire v$HALT_16371_out0;
wire v$HALT_17681_out0;
wire v$HALT_17682_out0;
wire v$HALT_2899_out0;
wire v$HALT_2900_out0;
wire v$HALT_7572_out0;
wire v$HALT_7573_out0;
wire v$HIGHER$OUT_3829_out0;
wire v$HIGHER$OUT_3830_out0;
wire v$HIGHER$OUT_3831_out0;
wire v$HIGHER$OUT_3832_out0;
wire v$HIGHER$OUT_3833_out0;
wire v$HIGHER$OUT_3834_out0;
wire v$HIGHER$OUT_3835_out0;
wire v$HIGHER$OUT_3836_out0;
wire v$HIGHER$OUT_7785_out0;
wire v$HIGHER$OUT_7786_out0;
wire v$HIGHER$OUT_7787_out0;
wire v$HIGHER$OUT_7788_out0;
wire v$HIGHER$SAME_15020_out0;
wire v$HIGHER$SAME_15021_out0;
wire v$HIGHER$SAME_15022_out0;
wire v$HIGHER$SAME_15023_out0;
wire v$HIGHER$SAME_15024_out0;
wire v$HIGHER$SAME_15025_out0;
wire v$HIGHER$SAME_15026_out0;
wire v$HIGHER$SAME_15027_out0;
wire v$HIGHER$SAME_9132_out0;
wire v$HIGHER$SAME_9133_out0;
wire v$HIGHER$SAME_9134_out0;
wire v$HIGHER$SAME_9135_out0;
wire v$I0EN_8042_out0;
wire v$I0EN_8043_out0;
wire v$I0P_10308_out0;
wire v$I0P_10309_out0;
wire v$I0P_2438_out0;
wire v$I0P_2439_out0;
wire v$I0P_4347_out0;
wire v$I0P_4348_out0;
wire v$I0REGISTERWRITE_3355_out0;
wire v$I0REGISTERWRITE_3356_out0;
wire v$I0_18506_out0;
wire v$I0_18507_out0;
wire v$I1EN_18402_out0;
wire v$I1EN_18403_out0;
wire v$I1P_14818_out0;
wire v$I1P_14819_out0;
wire v$I1P_2514_out0;
wire v$I1P_2515_out0;
wire v$I1P_6440_out0;
wire v$I1P_6441_out0;
wire v$I1REGISTERWRITE_2931_out0;
wire v$I1REGISTERWRITE_2932_out0;
wire v$I1_4890_out0;
wire v$I1_4891_out0;
wire v$I2EN_15746_out0;
wire v$I2EN_15747_out0;
wire v$I2P_2258_out0;
wire v$I2P_2259_out0;
wire v$I2P_6433_out0;
wire v$I2P_6434_out0;
wire v$I2P_7492_out0;
wire v$I2P_7493_out0;
wire v$I2REGISTERWRITE_11930_out0;
wire v$I2REGISTERWRITE_11931_out0;
wire v$I2_14493_out0;
wire v$I2_14494_out0;
wire v$I3EN_17775_out0;
wire v$I3EN_17776_out0;
wire v$I3P_10827_out0;
wire v$I3P_10828_out0;
wire v$I3P_13619_out0;
wire v$I3P_13620_out0;
wire v$I3P_8969_out0;
wire v$I3P_8970_out0;
wire v$I3REGISTERWRITE_1264_out0;
wire v$I3REGISTERWRITE_1265_out0;
wire v$I3_4823_out0;
wire v$I3_4824_out0;
wire v$IGNORE_11704_out0;
wire v$IGNORE_11705_out0;
wire v$IGNORE_16561_out0;
wire v$IGNORE_16562_out0;
wire v$IGNORE_5408_out0;
wire v$IGNORE_5409_out0;
wire v$IGNORE_8283_out0;
wire v$INCOMINGINTERRUPT_1903_out0;
wire v$INCOMINGINTERRUPT_1904_out0;
wire v$ININTERRUPT_1133_out0;
wire v$ININTERRUPT_1134_out0;
wire v$ININT_15465_out0;
wire v$ININT_15466_out0;
wire v$INITIAL$FETCH$OCCURRED_1537_out0;
wire v$INITIAL$FETCH$OCCURRED_1538_out0;
wire v$INIT_10752_out0;
wire v$INIT_10753_out0;
wire v$INT2_11881_out0;
wire v$INT2_3161_out0;
wire v$INT2_5407_out0;
wire v$INT3_14034_out0;
wire v$INT3_14035_out0;
wire v$INT3_18126_out0;
wire v$INT3_18127_out0;
wire v$INTCAPTURE0_13532_out0;
wire v$INTCAPTURE0_13533_out0;
wire v$INTCLEAR_7775_out0;
wire v$INTCLEAR_7776_out0;
wire v$INTCLR_214_out0;
wire v$INTCLR_215_out0;
wire v$INTCOUNT_7474_out0;
wire v$INTCOUNT_7475_out0;
wire v$INTDISABLE_2684_out0;
wire v$INTDISABLE_2685_out0;
wire v$INTDISABLE_4999_out0;
wire v$INTDISABLE_5000_out0;
wire v$INTENABLE_17402_out0;
wire v$INTENABLE_17403_out0;
wire v$INTENABLE_2939_out0;
wire v$INTENABLE_2940_out0;
wire v$INTERRUPT0_11700_out0;
wire v$INTERRUPT0_11701_out0;
wire v$INTERRUPT0_1805_out0;
wire v$INTERRUPT0_1806_out0;
wire v$INTERRUPT1_17700_out0;
wire v$INTERRUPT1_17701_out0;
wire v$INTERRUPT1_8284_out0;
wire v$INTERRUPT1_8285_out0;
wire v$INTERRUPT2_1663_out0;
wire v$INTERRUPT2_1664_out0;
wire v$INTERRUPT2_3853_out0;
wire v$INTERRUPT2_3854_out0;
wire v$INTERRUPT3_2816_out0;
wire v$INTERRUPT3_2817_out0;
wire v$INTERRUPT3_3508_out0;
wire v$INTERRUPT3_3509_out0;
wire v$INTERRUPTOVERFLOW_15112_out0;
wire v$INTERRUPTOVERFLOW_15113_out0;
wire v$INTERRUPTOVERFLOW_2233_out0;
wire v$INTERRUPTOVERFLOW_2234_out0;
wire v$INTERRUPTSENABLED_9620_out0;
wire v$INTERRUPTSENABLED_9621_out0;
wire v$INTOVERFLOW_16039_out0;
wire v$INTOVERFLOW_16040_out0;
wire v$IR1$15_5758_out0;
wire v$IR1$15_5759_out0;
wire v$IR1$32$BITS_5454_out0;
wire v$IR1$32$BITS_7867_out0;
wire v$IR1$C$L_10053_out0;
wire v$IR1$C$L_10054_out0;
wire v$IR1$IS$FPU$ARITHMETIC_1370_out0;
wire v$IR1$IS$FPU$ARITHMETIC_1371_out0;
wire v$IR1$IS$FPU$LOAD$STORE_8930_out0;
wire v$IR1$IS$LDST_13203_out0;
wire v$IR1$IS$LDST_13204_out0;
wire v$IR1$IS$STORE_4462_out0;
wire v$IR1$IS$STORE_4463_out0;
wire v$IR1$LS_16424_out0;
wire v$IR1$LS_16425_out0;
wire v$IR1$L_5138_out0;
wire v$IR1$L_5139_out0;
wire v$IR1$P_3692_out0;
wire v$IR1$P_3693_out0;
wire v$IR1$S$WB_322_out0;
wire v$IR1$S$WB_323_out0;
wire v$IR1$S_7842_out0;
wire v$IR1$S_7843_out0;
wire v$IR1$U_14776_out0;
wire v$IR1$U_14777_out0;
wire v$IR1$VALID$VIEWER_1613_out0;
wire v$IR1$VALID$VIEWER_1614_out0;
wire v$IR1$VALID_14013_out0;
wire v$IR1$VALID_14014_out0;
wire v$IR1$VALID_17797_out0;
wire v$IR1$VALID_17798_out0;
wire v$IR1$VALID_18427_out0;
wire v$IR1$VALID_18428_out0;
wire v$IR1$VALID_3847_out0;
wire v$IR1$VALID_3848_out0;
wire v$IR1$VALID_5751_out0;
wire v$IR1$VALID_5752_out0;
wire v$IR1$VALID_61_out0;
wire v$IR1$VALID_62_out0;
wire v$IR1$VALID_9455_out0;
wire v$IR1$VALID_9456_out0;
wire v$IR1$W_16548_out0;
wire v$IR1$W_16549_out0;
wire v$IR15_10688_out0;
wire v$IR15_10689_out0;
wire v$IR15_10986_out0;
wire v$IR15_10987_out0;
wire v$IR2$15_7435_out0;
wire v$IR2$15_7436_out0;
wire v$IR2$FPU$32BIT_11800_out0;
wire v$IR2$FPU$32BIT_11801_out0;
wire v$IR2$FPU$LOADA_15268_out0;
wire v$IR2$FPU$LOADA_15269_out0;
wire v$IR2$FPU$LOAD_4231_out0;
wire v$IR2$FPU$LOAD_4232_out0;
wire v$IR2$FPU$L_10744_out0;
wire v$IR2$FPU$L_10745_out0;
wire v$IR2$IS$FPU_11843_out0;
wire v$IR2$IS$FPU_11844_out0;
wire v$IR2$IS$FPU_2929_out0;
wire v$IR2$IS$FPU_2930_out0;
wire v$IR2$IS$FPU_7049_out0;
wire v$IR2$IS$FPU_7050_out0;
wire v$IR2$IS$LDST_4395_out0;
wire v$IR2$IS$LDST_4396_out0;
wire v$IR2$LS_15832_out0;
wire v$IR2$LS_15833_out0;
wire v$IR2$L_12464_out0;
wire v$IR2$L_12465_out0;
wire v$IR2$P_17316_out0;
wire v$IR2$P_17317_out0;
wire v$IR2$REG$IMMEDIATE_6195_out0;
wire v$IR2$REG$IMMEDIATE_6196_out0;
wire v$IR2$S$WB_17436_out0;
wire v$IR2$S$WB_17437_out0;
wire v$IR2$S_1169_out0;
wire v$IR2$S_1170_out0;
wire v$IR2$U_5904_out0;
wire v$IR2$U_5905_out0;
wire v$IR2$VALID$AND$NOT$FLOAD_4878_out0;
wire v$IR2$VALID$AND$NOT$FLOAD_4879_out0;
wire v$IR2$VALID$AND$NOT$FLOAD_7285_out0;
wire v$IR2$VALID$AND$NOT$FLOAD_7286_out0;
wire v$IR2$VALID$VIEWER_5800_out0;
wire v$IR2$VALID$VIEWER_5801_out0;
wire v$IR2$VALID_10666_out0;
wire v$IR2$VALID_10667_out0;
wire v$IR2$VALID_11794_out0;
wire v$IR2$VALID_11795_out0;
wire v$IR2$VALID_13250_out0;
wire v$IR2$VALID_13251_out0;
wire v$IR2$VALID_14823_out0;
wire v$IR2$VALID_14824_out0;
wire v$IR2$VALID_15878_out0;
wire v$IR2$VALID_15879_out0;
wire v$IR2$VALID_18756_out0;
wire v$IR2$VALID_18757_out0;
wire v$IR2$VALID_4217_out0;
wire v$IR2$VALID_4218_out0;
wire v$IR2$VALID_6455_out0;
wire v$IR2$VALID_6456_out0;
wire v$IR2$VALID_7421_out0;
wire v$IR2$VALID_7422_out0;
wire v$IR2$W_15109_out0;
wire v$IR2$W_15110_out0;
wire v$IS$32$BIT$FPU$ADDER_14967_out0;
wire v$IS$32$BIT$FPU$ADDER_14968_out0;
wire v$IS$32$BITS$VIEWER_1236_out0;
wire v$IS$32$BITS_1282_out0;
wire v$IS$32$BITS_14038_out0;
wire v$IS$32$BITS_14039_out0;
wire v$IS$32$BITS_17583_out0;
wire v$IS$32$BITS_17584_out0;
wire v$IS$32$BITS_2992_out0;
wire v$IS$32$BITS_4148_out0;
wire v$IS$32$BITS_4149_out0;
wire v$IS$32$BIT_10862_out0;
wire v$IS$32$BIT_10863_out0;
wire v$IS$32$BIT_11005_out0;
wire v$IS$32$BIT_11006_out0;
wire v$IS$A$LARGER_10444_out0;
wire v$IS$A$LARGER_10445_out0;
wire v$IS$A$LARGER_14661_out0;
wire v$IS$A$LARGER_14662_out0;
wire v$IS$A$LARGER_15988_out0;
wire v$IS$A$LARGER_15989_out0;
wire v$IS$A$LARGER_16832_out0;
wire v$IS$A$LARGER_16833_out0;
wire v$IS$A$LARGER_7072_out0;
wire v$IS$A$LARGER_7073_out0;
wire v$IS$FPU$HAZARD_342_out0;
wire v$IS$FPU$HAZARD_343_out0;
wire v$IS$IR1$FMUL_15296_out0;
wire v$IS$IR1$FMUL_15297_out0;
wire v$IS$IR1$FMUL_2964_out0;
wire v$IS$IR1$FMUL_2965_out0;
wire v$IS$IR2$DATA$PROCESSING_9944_out0;
wire v$IS$IR2$DATA$PROCESSING_9945_out0;
wire v$IS$SUB$MANTISA$ADDER_3169_out0;
wire v$IS$SUB$MANTISA$ADDER_3170_out0;
wire v$IS$SUB$VIEW_227_out0;
wire v$IS$SUB$VIEW_228_out0;
wire v$IS$SUB_13067_out0;
wire v$IS$SUB_13068_out0;
wire v$IS$SUB_15449_out0;
wire v$IS$SUB_15450_out0;
wire v$IS$SUB_4443_out0;
wire v$IS$SUB_4444_out0;
wire v$IS$SUM$0_15623_out0;
wire v$IS$SUM$0_15624_out0;
wire v$IS$SUM$0_15681_out0;
wire v$IS$SUM$0_15682_out0;
wire v$IS$SUM$0_897_out0;
wire v$IS$SUM$0_898_out0;
wire v$ISINTERRUPTED_11856_out0;
wire v$ISINTERRUPTED_11857_out0;
wire v$ISINTERRUPTED_11968_out0;
wire v$ISINTERRUPTED_11969_out0;
wire v$ISMOV_12630_out0;
wire v$ISMOV_12631_out0;
wire v$ISMOV_4078_out0;
wire v$ISMOV_4079_out0;
wire v$ISMOV_6670_out0;
wire v$ISMOV_6671_out0;
wire v$ISMOV_8767_out0;
wire v$ISMOV_8768_out0;
wire v$JEQ_1675_out0;
wire v$JEQ_1676_out0;
wire v$JEQ_18036_out0;
wire v$JEQ_18037_out0;
wire v$JLO_14983_out0;
wire v$JLO_14984_out0;
wire v$JLO_8109_out0;
wire v$JLO_8110_out0;
wire v$JLS_16442_out0;
wire v$JLS_16443_out0;
wire v$JLS_1955_out0;
wire v$JLS_1956_out0;
wire v$JMI_13149_out0;
wire v$JMI_13150_out0;
wire v$JMI_73_out0;
wire v$JMI_74_out0;
wire v$JMP_1667_out0;
wire v$JMP_1668_out0;
wire v$JMP_4337_out0;
wire v$JMP_4338_out0;
wire v$LASTQ_12098_out0;
wire v$LASTQ_12099_out0;
wire v$LASTQ_12100_out0;
wire v$LASTQ_12101_out0;
wire v$LASTQ_12102_out0;
wire v$LASTQ_12103_out0;
wire v$LASTQ_12104_out0;
wire v$LASTQ_12105_out0;
wire v$LASTQ_12106_out0;
wire v$LASTQ_12107_out0;
wire v$LASTQ_12108_out0;
wire v$LASTQ_12109_out0;
wire v$LASTQ_12110_out0;
wire v$LASTQ_12111_out0;
wire v$LASTQ_12112_out0;
wire v$LASTQ_12113_out0;
wire v$LASTQ_12114_out0;
wire v$LASTQ_12115_out0;
wire v$LASTQ_12116_out0;
wire v$LASTQ_12117_out0;
wire v$LASTQ_12118_out0;
wire v$LASTQ_12119_out0;
wire v$LDMAINPC_13634_out0;
wire v$LDMAINPC_13635_out0;
wire v$LDMAIN_13807_out0;
wire v$LDMAIN_13808_out0;
wire v$LDMAIN_3205_out0;
wire v$LDMAIN_3206_out0;
wire v$LDSTRAMMUX_16139_out0;
wire v$LDSTRAMMUX_16140_out0;
wire v$LEFT$SHIFT_12832_out0;
wire v$LEFT$SHIFT_12833_out0;
wire v$LEFT$SHIFT_12834_out0;
wire v$LEFT$SHIFT_12835_out0;
wire v$LEFT$SHIFT_12836_out0;
wire v$LEFT$SHIFT_12837_out0;
wire v$LEFT$SHIFT_12838_out0;
wire v$LEFT$SHIFT_12839_out0;
wire v$LEFT$SHIFT_8798_out0;
wire v$LEFT$SHIFT_8799_out0;
wire v$LEFT$SHIFT_8800_out0;
wire v$LEFT$SHIFT_8801_out0;
wire v$LEFT$SHIFT_8802_out0;
wire v$LEFT$SHIFT_8803_out0;
wire v$LEFT$SHIFT_8804_out0;
wire v$LEFT$SHIFT_8805_out0;
wire v$LEFT$SHIT_3041_out0;
wire v$LEFT$SHIT_3042_out0;
wire v$LEFT$SHIT_3043_out0;
wire v$LEFT$SHIT_3044_out0;
wire v$LEFT$SHIT_3045_out0;
wire v$LEFT$SHIT_3046_out0;
wire v$LEFT$SHIT_3047_out0;
wire v$LEFT$SHIT_3048_out0;
wire v$LEFT$SHIT_3049_out0;
wire v$LEFT$SHIT_3050_out0;
wire v$LEFT$SHIT_3051_out0;
wire v$LEFT$SHIT_3052_out0;
wire v$LEFT$SHIT_3053_out0;
wire v$LEFT$SHIT_3054_out0;
wire v$LEFT$SHIT_3055_out0;
wire v$LEFT$SHIT_3056_out0;
wire v$LEFT$SHIT_3057_out0;
wire v$LEFT$SHIT_3058_out0;
wire v$LEFT$SHIT_3059_out0;
wire v$LEFT$SHIT_3060_out0;
wire v$LEFT$SHIT_3061_out0;
wire v$LEFT$SHIT_3062_out0;
wire v$LEFT$SHIT_3063_out0;
wire v$LEFT$SHIT_3064_out0;
wire v$LEFT$SHIT_3065_out0;
wire v$LEFT$SHIT_3066_out0;
wire v$LEFT$SHIT_3067_out0;
wire v$LEFT$SHIT_3068_out0;
wire v$LEFT$SHIT_3069_out0;
wire v$LEFT$SHIT_3070_out0;
wire v$LEFT$SHIT_3071_out0;
wire v$LEFT$SHIT_3072_out0;
wire v$LEFT$SHIT_3073_out0;
wire v$LEFT$SHIT_3074_out0;
wire v$LEFT$SHIT_3075_out0;
wire v$LEFT$SHIT_3076_out0;
wire v$LEFT$SHIT_3077_out0;
wire v$LEFT$SHIT_3078_out0;
wire v$LEFT$SHIT_3079_out0;
wire v$LEFT$SHIT_3080_out0;
wire v$LEFT$SHIT_3081_out0;
wire v$LEFT$SHIT_3082_out0;
wire v$LEFT$SHIT_3083_out0;
wire v$LEFT$SHIT_3084_out0;
wire v$LEFT$SHIT_3085_out0;
wire v$LEFT$SHIT_3086_out0;
wire v$LEFT$SHIT_3087_out0;
wire v$LEFT$SHIT_3088_out0;
wire v$LEFT$SHIT_3089_out0;
wire v$LEFT$SHIT_3090_out0;
wire v$LEFT$SHIT_3091_out0;
wire v$LEFT$SHIT_3092_out0;
wire v$LEFT$SHIT_3093_out0;
wire v$LEFT$SHIT_3094_out0;
wire v$LEFT$SHIT_3095_out0;
wire v$LEFT$SHIT_3096_out0;
wire v$LEFT$SHIT_3097_out0;
wire v$LEFT$SHIT_3098_out0;
wire v$LEFT$SHIT_3099_out0;
wire v$LEFT$SHIT_3100_out0;
wire v$LEFT$SHIT_3101_out0;
wire v$LEFT$SHIT_3102_out0;
wire v$LEFT$SHIT_3103_out0;
wire v$LOADA_5076_out0;
wire v$LOADA_5077_out0;
wire v$LOADA_5145_out0;
wire v$LOADA_5146_out0;
wire v$LOAD_11702_out0;
wire v$LOAD_11703_out0;
wire v$LOAD_6190_out0;
wire v$LOAD_6191_out0;
wire v$LOWER$OUT_4221_out0;
wire v$LOWER$OUT_4222_out0;
wire v$LOWER$OUT_4223_out0;
wire v$LOWER$OUT_4224_out0;
wire v$LOWER$OUT_4225_out0;
wire v$LOWER$OUT_4226_out0;
wire v$LOWER$OUT_4227_out0;
wire v$LOWER$OUT_4228_out0;
wire v$LOWER$OUT_6422_out0;
wire v$LOWER$OUT_6423_out0;
wire v$LOWER$OUT_6424_out0;
wire v$LOWER$OUT_6425_out0;
wire v$LOWER$PART_6314_out0;
wire v$LOWER$PART_6315_out0;
wire v$LOWER$PART_6316_out0;
wire v$LOWER$PART_6317_out0;
wire v$LOWER$SAME_10181_out0;
wire v$LOWER$SAME_10182_out0;
wire v$LOWER$SAME_10183_out0;
wire v$LOWER$SAME_10184_out0;
wire v$LOWER$SAME_10185_out0;
wire v$LOWER$SAME_10186_out0;
wire v$LOWER$SAME_10187_out0;
wire v$LOWER$SAME_10188_out0;
wire v$LOWER$SAME_3793_out0;
wire v$LOWER$SAME_3794_out0;
wire v$LOWER$SAME_3795_out0;
wire v$LOWER$SAME_3796_out0;
wire v$LSB_7815_out0;
wire v$LSB_7816_out0;
wire v$MANTISA$SAME_2436_out0;
wire v$MANTISA$SAME_2437_out0;
wire v$MEMHALT_17799_out0;
wire v$MEMHALT_17800_out0;
wire v$MI$LDST_17013_out0;
wire v$MI$LDST_17014_out0;
wire v$MI_11878_out0;
wire v$MI_11879_out0;
wire v$MI_12128_out0;
wire v$MI_12129_out0;
wire v$MI_12466_out0;
wire v$MI_12467_out0;
wire v$MI_14365_out0;
wire v$MI_14366_out0;
wire v$MI_2416_out0;
wire v$MI_2417_out0;
wire v$MI_6238_out0;
wire v$MI_6239_out0;
wire v$MI_8450_out0;
wire v$MI_8451_out0;
wire v$MODEEN_15114_out0;
wire v$MODEEN_15115_out0;
wire v$MODEEN_5755_out0;
wire v$MODEEN_5756_out0;
wire v$MODEWRITE_14714_out0;
wire v$MODEWRITE_14715_out0;
wire v$MULTIPLYING$BIT_2849_out0;
wire v$MULTIPLYING$BIT_2850_out0;
wire v$MULTIPLYING$BIT_2851_out0;
wire v$MULTIPLYING$BIT_2852_out0;
wire v$MULTIPLYING$BIT_2853_out0;
wire v$MULTIPLYING$BIT_2854_out0;
wire v$MULTIPLYING$BIT_2855_out0;
wire v$MULTIPLYING$BIT_2856_out0;
wire v$MULTIPLYING$BIT_2857_out0;
wire v$MULTIPLYING$BIT_2858_out0;
wire v$MULTIPLYING$BIT_2859_out0;
wire v$MULTIPLYING$BIT_2860_out0;
wire v$MUL_17034_out0;
wire v$MUL_17035_out0;
wire v$MUX10_15672_out0;
wire v$MUX10_15673_out0;
wire v$MUX10_15674_out0;
wire v$MUX10_15675_out0;
wire v$MUX10_16397_out0;
wire v$MUX10_16398_out0;
wire v$MUX11_1204_out0;
wire v$MUX11_1205_out0;
wire v$MUX11_17933_out0;
wire v$MUX11_17934_out0;
wire v$MUX11_17935_out0;
wire v$MUX11_17936_out0;
wire v$MUX12_17813_out0;
wire v$MUX12_17814_out0;
wire v$MUX12_17815_out0;
wire v$MUX12_17816_out0;
wire v$MUX13_13682_out0;
wire v$MUX13_13683_out0;
wire v$MUX13_13684_out0;
wire v$MUX13_13685_out0;
wire v$MUX14_2957_out0;
wire v$MUX14_2958_out0;
wire v$MUX14_4919_out0;
wire v$MUX14_4920_out0;
wire v$MUX14_4921_out0;
wire v$MUX14_4922_out0;
wire v$MUX15_1317_out0;
wire v$MUX15_1318_out0;
wire v$MUX15_1319_out0;
wire v$MUX15_1320_out0;
wire v$MUX15_15925_out0;
wire v$MUX15_9403_out0;
wire v$MUX16_16762_out0;
wire v$MUX16_16763_out0;
wire v$MUX16_16764_out0;
wire v$MUX16_16765_out0;
wire v$MUX17_16536_out0;
wire v$MUX17_16537_out0;
wire v$MUX17_16538_out0;
wire v$MUX17_16539_out0;
wire v$MUX17_6531_out0;
wire v$MUX18_4858_out0;
wire v$MUX18_4859_out0;
wire v$MUX18_4860_out0;
wire v$MUX18_4861_out0;
wire v$MUX19_6374_out0;
wire v$MUX19_6375_out0;
wire v$MUX19_6376_out0;
wire v$MUX19_6377_out0;
wire v$MUX1_16952_out0;
wire v$MUX1_16953_out0;
wire v$MUX1_16954_out0;
wire v$MUX1_16955_out0;
wire v$MUX1_16956_out0;
wire v$MUX1_16957_out0;
wire v$MUX1_16958_out0;
wire v$MUX1_16959_out0;
wire v$MUX1_16960_out0;
wire v$MUX1_16961_out0;
wire v$MUX1_16962_out0;
wire v$MUX1_2582_out0;
wire v$MUX1_2583_out0;
wire v$MUX1_2584_out0;
wire v$MUX1_2585_out0;
wire v$MUX1_2586_out0;
wire v$MUX1_2587_out0;
wire v$MUX1_2588_out0;
wire v$MUX1_2589_out0;
wire v$MUX1_2590_out0;
wire v$MUX1_2591_out0;
wire v$MUX1_2592_out0;
wire v$MUX1_2593_out0;
wire v$MUX1_2865_out0;
wire v$MUX1_2866_out0;
wire v$MUX1_2867_out0;
wire v$MUX1_2868_out0;
wire v$MUX1_416_out0;
wire v$MUX1_417_out0;
wire v$MUX1_5013_out0;
wire v$MUX1_5014_out0;
wire v$MUX1_7642_out0;
wire v$MUX1_7643_out0;
wire v$MUX20_11364_out0;
wire v$MUX20_11365_out0;
wire v$MUX20_11366_out0;
wire v$MUX20_11367_out0;
wire v$MUX21_4902_out0;
wire v$MUX21_4903_out0;
wire v$MUX21_4904_out0;
wire v$MUX21_4905_out0;
wire v$MUX22_16464_out0;
wire v$MUX22_16465_out0;
wire v$MUX22_16466_out0;
wire v$MUX22_16467_out0;
wire v$MUX23_16223_out0;
wire v$MUX23_16224_out0;
wire v$MUX23_16225_out0;
wire v$MUX23_16226_out0;
wire v$MUX24_18056_out0;
wire v$MUX24_18057_out0;
wire v$MUX24_18058_out0;
wire v$MUX24_18059_out0;
wire v$MUX25_8404_out0;
wire v$MUX25_8405_out0;
wire v$MUX25_8406_out0;
wire v$MUX25_8407_out0;
wire v$MUX2_12234_out0;
wire v$MUX2_12235_out0;
wire v$MUX2_13287_out0;
wire v$MUX2_13288_out0;
wire v$MUX2_13608_out0;
wire v$MUX2_13609_out0;
wire v$MUX2_13610_out0;
wire v$MUX2_13611_out0;
wire v$MUX2_13819_out0;
wire v$MUX2_13820_out0;
wire v$MUX2_13821_out0;
wire v$MUX2_13822_out0;
wire v$MUX2_13823_out0;
wire v$MUX2_13824_out0;
wire v$MUX2_13825_out0;
wire v$MUX2_13826_out0;
wire v$MUX2_13827_out0;
wire v$MUX2_13828_out0;
wire v$MUX2_13829_out0;
wire v$MUX2_13830_out0;
wire v$MUX2_4852_out0;
wire v$MUX2_4853_out0;
wire v$MUX2_6685_out0;
wire v$MUX2_6686_out0;
wire v$MUX3_1428_out0;
wire v$MUX3_1429_out0;
wire v$MUX3_17725_out0;
wire v$MUX3_17726_out0;
wire v$MUX3_6131_out0;
wire v$MUX3_6132_out0;
wire v$MUX3_7600_out0;
wire v$MUX3_7601_out0;
wire v$MUX3_7602_out0;
wire v$MUX3_7603_out0;
wire v$MUX3_9950_out0;
wire v$MUX3_9951_out0;
wire v$MUX3_9952_out0;
wire v$MUX3_9953_out0;
wire v$MUX3_9954_out0;
wire v$MUX3_9955_out0;
wire v$MUX3_9956_out0;
wire v$MUX3_9957_out0;
wire v$MUX3_9958_out0;
wire v$MUX3_9959_out0;
wire v$MUX3_9960_out0;
wire v$MUX3_9961_out0;
wire v$MUX4_11648_out0;
wire v$MUX4_11649_out0;
wire v$MUX4_12637_out0;
wire v$MUX4_12638_out0;
wire v$MUX4_15635_out0;
wire v$MUX4_15636_out0;
wire v$MUX4_16847_out0;
wire v$MUX4_16848_out0;
wire v$MUX4_16849_out0;
wire v$MUX4_16850_out0;
wire v$MUX4_16851_out0;
wire v$MUX4_16852_out0;
wire v$MUX4_16853_out0;
wire v$MUX4_16854_out0;
wire v$MUX4_16855_out0;
wire v$MUX4_16856_out0;
wire v$MUX4_16857_out0;
wire v$MUX4_16858_out0;
wire v$MUX4_17084_out0;
wire v$MUX4_17085_out0;
wire v$MUX4_7799_out0;
wire v$MUX4_7800_out0;
wire v$MUX4_7801_out0;
wire v$MUX4_7802_out0;
wire v$MUX5_11847_out0;
wire v$MUX5_11848_out0;
wire v$MUX5_15500_out0;
wire v$MUX5_15501_out0;
wire v$MUX5_17066_out0;
wire v$MUX5_17067_out0;
wire v$MUX5_18559_out0;
wire v$MUX5_18560_out0;
wire v$MUX5_6928_out0;
wire v$MUX5_6929_out0;
wire v$MUX5_6930_out0;
wire v$MUX5_6931_out0;
wire v$MUX5_9524_out0;
wire v$MUX5_9525_out0;
wire v$MUX5_9526_out0;
wire v$MUX5_9527_out0;
wire v$MUX5_9528_out0;
wire v$MUX5_9529_out0;
wire v$MUX5_9530_out0;
wire v$MUX5_9531_out0;
wire v$MUX5_9532_out0;
wire v$MUX5_9533_out0;
wire v$MUX5_9534_out0;
wire v$MUX5_9535_out0;
wire v$MUX6_10388_out0;
wire v$MUX6_10389_out0;
wire v$MUX6_10390_out0;
wire v$MUX6_10391_out0;
wire v$MUX6_10392_out0;
wire v$MUX6_10393_out0;
wire v$MUX6_10394_out0;
wire v$MUX6_10395_out0;
wire v$MUX6_10396_out0;
wire v$MUX6_10397_out0;
wire v$MUX6_10398_out0;
wire v$MUX6_10399_out0;
wire v$MUX6_13557_out0;
wire v$MUX6_13558_out0;
wire v$MUX6_13737_out0;
wire v$MUX6_13738_out0;
wire v$MUX6_16285_out0;
wire v$MUX6_16286_out0;
wire v$MUX6_16287_out0;
wire v$MUX6_16288_out0;
wire v$MUX6_9130_out0;
wire v$MUX6_9131_out0;
wire v$MUX7_10965_out0;
wire v$MUX7_10966_out0;
wire v$MUX7_1227_out0;
wire v$MUX7_1228_out0;
wire v$MUX7_1229_out0;
wire v$MUX7_1230_out0;
wire v$MUX7_17903_out0;
wire v$MUX7_17904_out0;
wire v$MUX7_17905_out0;
wire v$MUX7_17906_out0;
wire v$MUX7_17907_out0;
wire v$MUX7_17908_out0;
wire v$MUX7_17909_out0;
wire v$MUX7_17910_out0;
wire v$MUX7_17911_out0;
wire v$MUX7_17912_out0;
wire v$MUX7_17913_out0;
wire v$MUX7_17914_out0;
wire v$MUX7_9480_out0;
wire v$MUX7_9481_out0;
wire v$MUX8$OUT_13424_out0;
wire v$MUX8$OUT_13425_out0;
wire v$MUX8_1496_out0;
wire v$MUX8_1497_out0;
wire v$MUX8_2945_out0;
wire v$MUX8_2946_out0;
wire v$MUX8_2947_out0;
wire v$MUX8_2948_out0;
wire v$MUX8_3603_out0;
wire v$MUX8_3604_out0;
wire v$MUX8_3605_out0;
wire v$MUX8_3606_out0;
wire v$MUX8_3607_out0;
wire v$MUX8_3608_out0;
wire v$MUX8_3609_out0;
wire v$MUX8_3610_out0;
wire v$MUX8_3611_out0;
wire v$MUX8_3612_out0;
wire v$MUX8_3613_out0;
wire v$MUX8_3614_out0;
wire v$MUX8_4349_out0;
wire v$MUX8_4350_out0;
wire v$MUX9_8243_out0;
wire v$MUX9_8244_out0;
wire v$MUX9_8245_out0;
wire v$MUX9_8246_out0;
wire v$ModeRegAdd_4007_out0;
wire v$ModeRegAdd_4008_out0;
wire v$ModeWrite_4452_out0;
wire v$ModeWrite_4453_out0;
wire v$NEED$SHIFT$OP1_4821_out0;
wire v$NEED$SHIFT$OP1_4822_out0;
wire v$NEWINTERRUPT_4431_out0;
wire v$NEWINTERRUPT_4432_out0;
wire v$NEWINTERRUPT_5432_out0;
wire v$NEWINTERRUPT_5433_out0;
wire v$NEWINTERRUPT_7025_out0;
wire v$NEWINTERRUPT_7026_out0;
wire v$NEWINT_17801_out0;
wire v$NEWINT_17802_out0;
wire v$NEXTINTERRUPT_12752_out0;
wire v$NEXTINTERRUPT_12753_out0;
wire v$NEXTINTERRUPT_16777_out0;
wire v$NEXTINTERRUPT_16778_out0;
wire v$NEXTINTERRUPT_18433_out0;
wire v$NEXTINTERRUPT_18434_out0;
wire v$NEXTINTERRUPT_18546_out0;
wire v$NEXTINTERRUPT_18547_out0;
wire v$NEXTINT_7001_out0;
wire v$NEXTINT_7002_out0;
wire v$NEXTSTATE_13535_out0;
wire v$NEXTSTATE_13536_out0;
wire v$NEXTSTATE_13537_out0;
wire v$NEXTSTATE_13538_out0;
wire v$NEXTSTATE_13539_out0;
wire v$NE_3429_out0;
wire v$NE_3430_out0;
wire v$NF_14564_out0;
wire v$NF_14565_out0;
wire v$NOT$USED$CARRY_18775_out0;
wire v$NOT$USED$CARRY_18776_out0;
wire v$NOT$USED$CARRY_18777_out0;
wire v$NOT$USED$CARRY_18778_out0;
wire v$NOT$USED1_14378_out0;
wire v$NOT$USED1_14379_out0;
wire v$NOT$USED1_14380_out0;
wire v$NOT$USED1_14381_out0;
wire v$NOT$USED1_14382_out0;
wire v$NOT$USED1_14383_out0;
wire v$NOT$USED1_14384_out0;
wire v$NOT$USED1_14385_out0;
wire v$NOT$USED_15950_out0;
wire v$NOT$USED_15951_out0;
wire v$NOT$USED_15952_out0;
wire v$NOT$USED_15953_out0;
wire v$NOT$USED_2891_out0;
wire v$NOT$USED_2892_out0;
wire v$NOT$USED_5449_out0;
wire v$NOT$USED_5450_out0;
wire v$NP_7258_out0;
wire v$NP_7259_out0;
wire v$NQ0_15381_out0;
wire v$NQ0_15382_out0;
wire v$NQ0_15621_out0;
wire v$NQ0_15622_out0;
wire v$NQ0_7796_out0;
wire v$NQ0_7797_out0;
wire v$NQ1_11038_out0;
wire v$NQ1_11039_out0;
wire v$NQ1_16729_out0;
wire v$NQ1_16730_out0;
wire v$NQ1_254_out0;
wire v$NQ1_255_out0;
wire v$NQ2_16698_out0;
wire v$NQ2_16699_out0;
wire v$NQ2_18563_out0;
wire v$NQ2_18564_out0;
wire v$NQ2_2980_out0;
wire v$NQ2_2981_out0;
wire v$NQ3_1491_out0;
wire v$NQ3_1492_out0;
wire v$NQ3_2998_out0;
wire v$NQ3_2999_out0;
wire v$NR_16656_out0;
wire v$NR_16657_out0;
wire v$NS_18201_out0;
wire v$NS_18202_out0;
wire v$ODDPARITY_15928_out0;
wire v$ODDPARITY_15929_out0;
wire v$OFF_4039_out0;
wire v$OFF_4040_out0;
wire v$OUTPUT_10339_out0;
wire v$OUTPUT_10340_out0;
wire v$OUTPUT_10341_out0;
wire v$OUTPUT_10342_out0;
wire v$OUTPUT_18477_out0;
wire v$OUT_13756_out0;
wire v$OUT_13757_out0;
wire v$OUT_13758_out0;
wire v$OUT_13759_out0;
wire v$OUT_13760_out0;
wire v$OUT_13761_out0;
wire v$OUT_13762_out0;
wire v$OUT_13763_out0;
wire v$OUT_3840_out0;
wire v$OUT_3841_out0;
wire v$OUT_3906_out0;
wire v$OUT_3907_out0;
wire v$OUT_3908_out0;
wire v$OUT_3909_out0;
wire v$OUT_3910_out0;
wire v$OUT_3911_out0;
wire v$OUT_3912_out0;
wire v$OUT_3913_out0;
wire v$OUT_3914_out0;
wire v$OUT_3915_out0;
wire v$OUT_3916_out0;
wire v$OUT_3917_out0;
wire v$OUT_3918_out0;
wire v$OUT_3919_out0;
wire v$OUT_3920_out0;
wire v$OUT_3921_out0;
wire v$OUT_3922_out0;
wire v$OUT_3923_out0;
wire v$OUT_3924_out0;
wire v$OUT_3925_out0;
wire v$OUT_3926_out0;
wire v$OUT_3927_out0;
wire v$OUT_3928_out0;
wire v$OUT_3929_out0;
wire v$OUT_3930_out0;
wire v$OUT_3931_out0;
wire v$OUT_3932_out0;
wire v$OUT_3933_out0;
wire v$OUT_3934_out0;
wire v$OUT_3935_out0;
wire v$OUT_3936_out0;
wire v$OUT_3937_out0;
wire v$OUT_8937_out0;
wire v$OUT_8938_out0;
wire v$OUT_8939_out0;
wire v$OUT_8940_out0;
wire v$OUT_9476_out0;
wire v$OUT_9477_out0;
wire v$OUT_9478_out0;
wire v$OUT_9479_out0;
wire v$OVERFLOW_14976_out0;
wire v$OVERFLOW_14977_out0;
wire v$OVERFLOW_18455_out0;
wire v$OVERFLOW_18456_out0;
wire v$OVERFLOW_18525_out0;
wire v$OVERFLOW_18526_out0;
wire v$OVERFLOW_3630_out0;
wire v$OVERFLOW_3631_out0;
wire v$OVERFLOW_426_out0;
wire v$OVERFLOW_427_out0;
wire v$OddParity_10686_out0;
wire v$OddParity_10687_out0;
wire v$P$AB_2001_out0;
wire v$P$AB_2002_out0;
wire v$P$AB_2003_out0;
wire v$P$AB_2004_out0;
wire v$P$AB_2005_out0;
wire v$P$AB_2006_out0;
wire v$P$AB_2007_out0;
wire v$P$AB_2008_out0;
wire v$P$AB_2009_out0;
wire v$P$AB_2010_out0;
wire v$P$AB_2011_out0;
wire v$P$AB_2012_out0;
wire v$P$AB_2013_out0;
wire v$P$AB_2014_out0;
wire v$P$AB_2015_out0;
wire v$P$AB_2016_out0;
wire v$P$AB_2017_out0;
wire v$P$AB_2018_out0;
wire v$P$AB_2019_out0;
wire v$P$AB_2020_out0;
wire v$P$AB_2021_out0;
wire v$P$AB_2022_out0;
wire v$P$AB_2023_out0;
wire v$P$AB_2024_out0;
wire v$P$AB_2025_out0;
wire v$P$AB_2026_out0;
wire v$P$AB_2027_out0;
wire v$P$AB_2028_out0;
wire v$P$AB_2029_out0;
wire v$P$AB_2030_out0;
wire v$P$AB_2031_out0;
wire v$P$AB_2032_out0;
wire v$P$AB_2033_out0;
wire v$P$AB_2034_out0;
wire v$P$AB_2035_out0;
wire v$P$AB_2036_out0;
wire v$P$AB_2037_out0;
wire v$P$AB_2038_out0;
wire v$P$AB_2039_out0;
wire v$P$AB_2040_out0;
wire v$P$AB_2041_out0;
wire v$P$AB_2042_out0;
wire v$P$AB_2043_out0;
wire v$P$AB_2044_out0;
wire v$P$AB_2045_out0;
wire v$P$AB_2046_out0;
wire v$P$AB_2047_out0;
wire v$P$AB_2048_out0;
wire v$P$AB_2049_out0;
wire v$P$AB_2050_out0;
wire v$P$AB_2051_out0;
wire v$P$AB_2052_out0;
wire v$P$AB_2053_out0;
wire v$P$AB_2054_out0;
wire v$P$AB_2055_out0;
wire v$P$AB_2056_out0;
wire v$P$AB_2057_out0;
wire v$P$AB_2058_out0;
wire v$P$AB_2059_out0;
wire v$P$AB_2060_out0;
wire v$P$AB_2061_out0;
wire v$P$AB_2062_out0;
wire v$P$AB_2063_out0;
wire v$P$AB_2064_out0;
wire v$P$AB_2065_out0;
wire v$P$AB_2066_out0;
wire v$P$AB_2067_out0;
wire v$P$AB_2068_out0;
wire v$P$AB_2069_out0;
wire v$P$AB_2070_out0;
wire v$P$AB_2071_out0;
wire v$P$AB_2072_out0;
wire v$P$AB_2073_out0;
wire v$P$AB_2074_out0;
wire v$P$AB_2075_out0;
wire v$P$AB_2076_out0;
wire v$P$AB_2077_out0;
wire v$P$AB_2078_out0;
wire v$P$AB_2079_out0;
wire v$P$AB_2080_out0;
wire v$P$AB_2081_out0;
wire v$P$AB_2082_out0;
wire v$P$AB_2083_out0;
wire v$P$AB_2084_out0;
wire v$P$AB_2085_out0;
wire v$P$AB_2086_out0;
wire v$P$AB_2087_out0;
wire v$P$AB_2088_out0;
wire v$P$AB_2089_out0;
wire v$P$AB_2090_out0;
wire v$P$AB_2091_out0;
wire v$P$AB_2092_out0;
wire v$P$AB_2093_out0;
wire v$P$AB_2094_out0;
wire v$P$AB_2095_out0;
wire v$P$AB_2096_out0;
wire v$P$AB_2097_out0;
wire v$P$AB_2098_out0;
wire v$P$AB_2099_out0;
wire v$P$AB_2100_out0;
wire v$P$AB_2101_out0;
wire v$P$AB_2102_out0;
wire v$P$AB_2103_out0;
wire v$P$AB_2104_out0;
wire v$P$AB_2105_out0;
wire v$P$AB_2106_out0;
wire v$P$AB_2107_out0;
wire v$P$AB_2108_out0;
wire v$P$AB_2109_out0;
wire v$P$AB_2110_out0;
wire v$P$AB_2111_out0;
wire v$P$AB_2112_out0;
wire v$P$AB_2113_out0;
wire v$P$AB_2114_out0;
wire v$P$AB_2115_out0;
wire v$P$AB_2116_out0;
wire v$P$AB_2117_out0;
wire v$P$AB_2118_out0;
wire v$P$AB_2119_out0;
wire v$P$AB_2120_out0;
wire v$P$AB_2121_out0;
wire v$P$AB_2122_out0;
wire v$P$AB_2123_out0;
wire v$P$AB_2124_out0;
wire v$P$AB_2125_out0;
wire v$P$AB_2126_out0;
wire v$P$AB_2127_out0;
wire v$P$AB_2128_out0;
wire v$P$AB_2129_out0;
wire v$P$AB_2130_out0;
wire v$P$AB_2131_out0;
wire v$P$AB_2132_out0;
wire v$P$AB_2133_out0;
wire v$P$AB_2134_out0;
wire v$P$AB_2135_out0;
wire v$P$AB_2136_out0;
wire v$P$AB_2137_out0;
wire v$P$AB_2138_out0;
wire v$P$AB_2139_out0;
wire v$P$AB_2140_out0;
wire v$P$AB_2141_out0;
wire v$P$AB_2142_out0;
wire v$P$AB_2143_out0;
wire v$P$AB_2144_out0;
wire v$P$AB_2145_out0;
wire v$P$AB_2146_out0;
wire v$P$AB_2147_out0;
wire v$P$AB_2148_out0;
wire v$P$AB_2149_out0;
wire v$P$AB_2150_out0;
wire v$P$AB_2151_out0;
wire v$P$AB_2152_out0;
wire v$P$AB_2153_out0;
wire v$P$AB_2154_out0;
wire v$P$AB_2155_out0;
wire v$P$AB_2156_out0;
wire v$P$AB_2157_out0;
wire v$P$AB_2158_out0;
wire v$P$AB_2159_out0;
wire v$P$AB_2160_out0;
wire v$P$AB_2161_out0;
wire v$P$AB_2162_out0;
wire v$P$AB_2163_out0;
wire v$P$AB_2164_out0;
wire v$P$AB_2165_out0;
wire v$P$AB_2166_out0;
wire v$P$AB_2167_out0;
wire v$P$AB_2168_out0;
wire v$P$AB_2169_out0;
wire v$P$AB_2170_out0;
wire v$P$AB_2171_out0;
wire v$P$AB_2172_out0;
wire v$P$AB_2173_out0;
wire v$P$AB_2174_out0;
wire v$P$AB_2175_out0;
wire v$P$AB_2176_out0;
wire v$P$AB_2177_out0;
wire v$P$AB_2178_out0;
wire v$P$AB_2179_out0;
wire v$P$AB_2180_out0;
wire v$P$AB_2181_out0;
wire v$P$AB_2182_out0;
wire v$P$AB_2183_out0;
wire v$P$AB_2184_out0;
wire v$P$AB_2185_out0;
wire v$P$AB_2186_out0;
wire v$P$AB_2187_out0;
wire v$P$AB_2188_out0;
wire v$P$AB_2189_out0;
wire v$P$AB_2190_out0;
wire v$P$AB_2191_out0;
wire v$P$AB_2192_out0;
wire v$P$AB_2193_out0;
wire v$P$AB_2194_out0;
wire v$P$AB_2195_out0;
wire v$P$AB_2196_out0;
wire v$P$AB_2197_out0;
wire v$P$AB_2198_out0;
wire v$P$AB_2199_out0;
wire v$P$AB_2200_out0;
wire v$P$AB_2201_out0;
wire v$P$AB_2202_out0;
wire v$P$AB_2203_out0;
wire v$P$AB_2204_out0;
wire v$P$AB_2205_out0;
wire v$P$AD_687_out0;
wire v$P$AD_688_out0;
wire v$P$AD_689_out0;
wire v$P$AD_690_out0;
wire v$P$AD_691_out0;
wire v$P$AD_692_out0;
wire v$P$AD_693_out0;
wire v$P$AD_694_out0;
wire v$P$AD_695_out0;
wire v$P$AD_696_out0;
wire v$P$AD_697_out0;
wire v$P$AD_698_out0;
wire v$P$AD_699_out0;
wire v$P$AD_700_out0;
wire v$P$AD_701_out0;
wire v$P$AD_702_out0;
wire v$P$AD_703_out0;
wire v$P$AD_704_out0;
wire v$P$AD_705_out0;
wire v$P$AD_706_out0;
wire v$P$AD_707_out0;
wire v$P$AD_708_out0;
wire v$P$AD_709_out0;
wire v$P$AD_710_out0;
wire v$P$AD_711_out0;
wire v$P$AD_712_out0;
wire v$P$AD_713_out0;
wire v$P$AD_714_out0;
wire v$P$AD_715_out0;
wire v$P$AD_716_out0;
wire v$P$AD_717_out0;
wire v$P$AD_718_out0;
wire v$P$AD_719_out0;
wire v$P$AD_720_out0;
wire v$P$AD_721_out0;
wire v$P$AD_722_out0;
wire v$P$AD_723_out0;
wire v$P$AD_724_out0;
wire v$P$AD_725_out0;
wire v$P$AD_726_out0;
wire v$P$AD_727_out0;
wire v$P$AD_728_out0;
wire v$P$AD_729_out0;
wire v$P$AD_730_out0;
wire v$P$AD_731_out0;
wire v$P$AD_732_out0;
wire v$P$AD_733_out0;
wire v$P$AD_734_out0;
wire v$P$AD_735_out0;
wire v$P$AD_736_out0;
wire v$P$AD_737_out0;
wire v$P$AD_738_out0;
wire v$P$AD_739_out0;
wire v$P$AD_740_out0;
wire v$P$AD_741_out0;
wire v$P$AD_742_out0;
wire v$P$AD_743_out0;
wire v$P$AD_744_out0;
wire v$P$AD_745_out0;
wire v$P$AD_746_out0;
wire v$P$AD_747_out0;
wire v$P$AD_748_out0;
wire v$P$AD_749_out0;
wire v$P$AD_750_out0;
wire v$P$AD_751_out0;
wire v$P$AD_752_out0;
wire v$P$AD_753_out0;
wire v$P$AD_754_out0;
wire v$P$AD_755_out0;
wire v$P$AD_756_out0;
wire v$P$AD_757_out0;
wire v$P$AD_758_out0;
wire v$P$AD_759_out0;
wire v$P$AD_760_out0;
wire v$P$AD_761_out0;
wire v$P$AD_762_out0;
wire v$P$AD_763_out0;
wire v$P$AD_764_out0;
wire v$P$AD_765_out0;
wire v$P$AD_766_out0;
wire v$P$AD_767_out0;
wire v$P$AD_768_out0;
wire v$P$AD_769_out0;
wire v$P$AD_770_out0;
wire v$P$AD_771_out0;
wire v$P$AD_772_out0;
wire v$P$AD_773_out0;
wire v$P$AD_774_out0;
wire v$P$AD_775_out0;
wire v$P$AD_776_out0;
wire v$P$AD_777_out0;
wire v$P$AD_778_out0;
wire v$P$AD_779_out0;
wire v$P$AD_780_out0;
wire v$P$AD_781_out0;
wire v$P$AD_782_out0;
wire v$P$AD_783_out0;
wire v$P$AD_784_out0;
wire v$P$AD_785_out0;
wire v$P$AD_786_out0;
wire v$P$AD_787_out0;
wire v$P$AD_788_out0;
wire v$P$AD_789_out0;
wire v$P$AD_790_out0;
wire v$P$AD_791_out0;
wire v$P$AD_792_out0;
wire v$P$AD_793_out0;
wire v$P$AD_794_out0;
wire v$P$AD_795_out0;
wire v$P$AD_796_out0;
wire v$P$AD_797_out0;
wire v$P$AD_798_out0;
wire v$P$AD_799_out0;
wire v$P$AD_800_out0;
wire v$P$AD_801_out0;
wire v$P$AD_802_out0;
wire v$P$AD_803_out0;
wire v$P$AD_804_out0;
wire v$P$AD_805_out0;
wire v$P$AD_806_out0;
wire v$P$AD_807_out0;
wire v$P$AD_808_out0;
wire v$P$AD_809_out0;
wire v$P$AD_810_out0;
wire v$P$AD_811_out0;
wire v$P$AD_812_out0;
wire v$P$AD_813_out0;
wire v$P$AD_814_out0;
wire v$P$AD_815_out0;
wire v$P$AD_816_out0;
wire v$P$AD_817_out0;
wire v$P$AD_818_out0;
wire v$P$AD_819_out0;
wire v$P$AD_820_out0;
wire v$P$AD_821_out0;
wire v$P$AD_822_out0;
wire v$P$AD_823_out0;
wire v$P$AD_824_out0;
wire v$P$AD_825_out0;
wire v$P$AD_826_out0;
wire v$P$AD_827_out0;
wire v$P$AD_828_out0;
wire v$P$AD_829_out0;
wire v$P$AD_830_out0;
wire v$P$AD_831_out0;
wire v$P$AD_832_out0;
wire v$P$AD_833_out0;
wire v$P$AD_834_out0;
wire v$P$AD_835_out0;
wire v$P$AD_836_out0;
wire v$P$AD_837_out0;
wire v$P$AD_838_out0;
wire v$P$AD_839_out0;
wire v$P$AD_840_out0;
wire v$P$AD_841_out0;
wire v$P$AD_842_out0;
wire v$P$AD_843_out0;
wire v$P$AD_844_out0;
wire v$P$AD_845_out0;
wire v$P$AD_846_out0;
wire v$P$AD_847_out0;
wire v$P$AD_848_out0;
wire v$P$AD_849_out0;
wire v$P$AD_850_out0;
wire v$P$AD_851_out0;
wire v$P$AD_852_out0;
wire v$P$AD_853_out0;
wire v$P$AD_854_out0;
wire v$P$AD_855_out0;
wire v$P$AD_856_out0;
wire v$P$AD_857_out0;
wire v$P$AD_858_out0;
wire v$P$AD_859_out0;
wire v$P$AD_860_out0;
wire v$P$AD_861_out0;
wire v$P$AD_862_out0;
wire v$P$AD_863_out0;
wire v$P$AD_864_out0;
wire v$P$AD_865_out0;
wire v$P$AD_866_out0;
wire v$P$AD_867_out0;
wire v$P$AD_868_out0;
wire v$P$AD_869_out0;
wire v$P$AD_870_out0;
wire v$P$AD_871_out0;
wire v$P$AD_872_out0;
wire v$P$AD_873_out0;
wire v$P$AD_874_out0;
wire v$P$AD_875_out0;
wire v$P$AD_876_out0;
wire v$P$AD_877_out0;
wire v$P$AD_878_out0;
wire v$P$AD_879_out0;
wire v$P$AD_880_out0;
wire v$P$AD_881_out0;
wire v$P$AD_882_out0;
wire v$P$AD_883_out0;
wire v$P$AD_884_out0;
wire v$P$AD_885_out0;
wire v$P$AD_886_out0;
wire v$P$AD_887_out0;
wire v$P$AD_888_out0;
wire v$P$AD_889_out0;
wire v$P$AD_890_out0;
wire v$P$AD_891_out0;
wire v$P$CD_10454_out0;
wire v$P$CD_10455_out0;
wire v$P$CD_10456_out0;
wire v$P$CD_10457_out0;
wire v$P$CD_10458_out0;
wire v$P$CD_10459_out0;
wire v$P$CD_10460_out0;
wire v$P$CD_10461_out0;
wire v$P$CD_10462_out0;
wire v$P$CD_10463_out0;
wire v$P$CD_10464_out0;
wire v$P$CD_10465_out0;
wire v$P$CD_10466_out0;
wire v$P$CD_10467_out0;
wire v$P$CD_10468_out0;
wire v$P$CD_10469_out0;
wire v$P$CD_10470_out0;
wire v$P$CD_10471_out0;
wire v$P$CD_10472_out0;
wire v$P$CD_10473_out0;
wire v$P$CD_10474_out0;
wire v$P$CD_10475_out0;
wire v$P$CD_10476_out0;
wire v$P$CD_10477_out0;
wire v$P$CD_10478_out0;
wire v$P$CD_10479_out0;
wire v$P$CD_10480_out0;
wire v$P$CD_10481_out0;
wire v$P$CD_10482_out0;
wire v$P$CD_10483_out0;
wire v$P$CD_10484_out0;
wire v$P$CD_10485_out0;
wire v$P$CD_10486_out0;
wire v$P$CD_10487_out0;
wire v$P$CD_10488_out0;
wire v$P$CD_10489_out0;
wire v$P$CD_10490_out0;
wire v$P$CD_10491_out0;
wire v$P$CD_10492_out0;
wire v$P$CD_10493_out0;
wire v$P$CD_10494_out0;
wire v$P$CD_10495_out0;
wire v$P$CD_10496_out0;
wire v$P$CD_10497_out0;
wire v$P$CD_10498_out0;
wire v$P$CD_10499_out0;
wire v$P$CD_10500_out0;
wire v$P$CD_10501_out0;
wire v$P$CD_10502_out0;
wire v$P$CD_10503_out0;
wire v$P$CD_10504_out0;
wire v$P$CD_10505_out0;
wire v$P$CD_10506_out0;
wire v$P$CD_10507_out0;
wire v$P$CD_10508_out0;
wire v$P$CD_10509_out0;
wire v$P$CD_10510_out0;
wire v$P$CD_10511_out0;
wire v$P$CD_10512_out0;
wire v$P$CD_10513_out0;
wire v$P$CD_10514_out0;
wire v$P$CD_10515_out0;
wire v$P$CD_10516_out0;
wire v$P$CD_10517_out0;
wire v$P$CD_10518_out0;
wire v$P$CD_10519_out0;
wire v$P$CD_10520_out0;
wire v$P$CD_10521_out0;
wire v$P$CD_10522_out0;
wire v$P$CD_10523_out0;
wire v$P$CD_10524_out0;
wire v$P$CD_10525_out0;
wire v$P$CD_10526_out0;
wire v$P$CD_10527_out0;
wire v$P$CD_10528_out0;
wire v$P$CD_10529_out0;
wire v$P$CD_10530_out0;
wire v$P$CD_10531_out0;
wire v$P$CD_10532_out0;
wire v$P$CD_10533_out0;
wire v$P$CD_10534_out0;
wire v$P$CD_10535_out0;
wire v$P$CD_10536_out0;
wire v$P$CD_10537_out0;
wire v$P$CD_10538_out0;
wire v$P$CD_10539_out0;
wire v$P$CD_10540_out0;
wire v$P$CD_10541_out0;
wire v$P$CD_10542_out0;
wire v$P$CD_10543_out0;
wire v$P$CD_10544_out0;
wire v$P$CD_10545_out0;
wire v$P$CD_10546_out0;
wire v$P$CD_10547_out0;
wire v$P$CD_10548_out0;
wire v$P$CD_10549_out0;
wire v$P$CD_10550_out0;
wire v$P$CD_10551_out0;
wire v$P$CD_10552_out0;
wire v$P$CD_10553_out0;
wire v$P$CD_10554_out0;
wire v$P$CD_10555_out0;
wire v$P$CD_10556_out0;
wire v$P$CD_10557_out0;
wire v$P$CD_10558_out0;
wire v$P$CD_10559_out0;
wire v$P$CD_10560_out0;
wire v$P$CD_10561_out0;
wire v$P$CD_10562_out0;
wire v$P$CD_10563_out0;
wire v$P$CD_10564_out0;
wire v$P$CD_10565_out0;
wire v$P$CD_10566_out0;
wire v$P$CD_10567_out0;
wire v$P$CD_10568_out0;
wire v$P$CD_10569_out0;
wire v$P$CD_10570_out0;
wire v$P$CD_10571_out0;
wire v$P$CD_10572_out0;
wire v$P$CD_10573_out0;
wire v$P$CD_10574_out0;
wire v$P$CD_10575_out0;
wire v$P$CD_10576_out0;
wire v$P$CD_10577_out0;
wire v$P$CD_10578_out0;
wire v$P$CD_10579_out0;
wire v$P$CD_10580_out0;
wire v$P$CD_10581_out0;
wire v$P$CD_10582_out0;
wire v$P$CD_10583_out0;
wire v$P$CD_10584_out0;
wire v$P$CD_10585_out0;
wire v$P$CD_10586_out0;
wire v$P$CD_10587_out0;
wire v$P$CD_10588_out0;
wire v$P$CD_10589_out0;
wire v$P$CD_10590_out0;
wire v$P$CD_10591_out0;
wire v$P$CD_10592_out0;
wire v$P$CD_10593_out0;
wire v$P$CD_10594_out0;
wire v$P$CD_10595_out0;
wire v$P$CD_10596_out0;
wire v$P$CD_10597_out0;
wire v$P$CD_10598_out0;
wire v$P$CD_10599_out0;
wire v$P$CD_10600_out0;
wire v$P$CD_10601_out0;
wire v$P$CD_10602_out0;
wire v$P$CD_10603_out0;
wire v$P$CD_10604_out0;
wire v$P$CD_10605_out0;
wire v$P$CD_10606_out0;
wire v$P$CD_10607_out0;
wire v$P$CD_10608_out0;
wire v$P$CD_10609_out0;
wire v$P$CD_10610_out0;
wire v$P$CD_10611_out0;
wire v$P$CD_10612_out0;
wire v$P$CD_10613_out0;
wire v$P$CD_10614_out0;
wire v$P$CD_10615_out0;
wire v$P$CD_10616_out0;
wire v$P$CD_10617_out0;
wire v$P$CD_10618_out0;
wire v$P$CD_10619_out0;
wire v$P$CD_10620_out0;
wire v$P$CD_10621_out0;
wire v$P$CD_10622_out0;
wire v$P$CD_10623_out0;
wire v$P$CD_10624_out0;
wire v$P$CD_10625_out0;
wire v$P$CD_10626_out0;
wire v$P$CD_10627_out0;
wire v$P$CD_10628_out0;
wire v$P$CD_10629_out0;
wire v$P$CD_10630_out0;
wire v$P$CD_10631_out0;
wire v$P$CD_10632_out0;
wire v$P$CD_10633_out0;
wire v$P$CD_10634_out0;
wire v$P$CD_10635_out0;
wire v$P$CD_10636_out0;
wire v$P$CD_10637_out0;
wire v$P$CD_10638_out0;
wire v$P$CD_10639_out0;
wire v$P$CD_10640_out0;
wire v$P$CD_10641_out0;
wire v$P$CD_10642_out0;
wire v$P$CD_10643_out0;
wire v$P$CD_10644_out0;
wire v$P$CD_10645_out0;
wire v$P$CD_10646_out0;
wire v$P$CD_10647_out0;
wire v$P$CD_10648_out0;
wire v$P$CD_10649_out0;
wire v$P$CD_10650_out0;
wire v$P$CD_10651_out0;
wire v$P$CD_10652_out0;
wire v$P$CD_10653_out0;
wire v$P$CD_10654_out0;
wire v$P$CD_10655_out0;
wire v$P$CD_10656_out0;
wire v$P$CD_10657_out0;
wire v$P$CD_10658_out0;
wire v$P0_4810_out0;
wire v$P0_4811_out0;
wire v$P0_4812_out0;
wire v$P0_4813_out0;
wire v$P0_4814_out0;
wire v$P10_344_out0;
wire v$P10_345_out0;
wire v$P10_346_out0;
wire v$P10_347_out0;
wire v$P10_348_out0;
wire v$P11_9611_out0;
wire v$P11_9612_out0;
wire v$P11_9613_out0;
wire v$P11_9614_out0;
wire v$P11_9615_out0;
wire v$P12_235_out0;
wire v$P12_236_out0;
wire v$P12_237_out0;
wire v$P12_238_out0;
wire v$P12_239_out0;
wire v$P13_3032_out0;
wire v$P13_3033_out0;
wire v$P13_3034_out0;
wire v$P13_3035_out0;
wire v$P13_3036_out0;
wire v$P14_3151_out0;
wire v$P14_3152_out0;
wire v$P14_3153_out0;
wire v$P14_3154_out0;
wire v$P14_3155_out0;
wire v$P15_6904_out0;
wire v$P15_6905_out0;
wire v$P15_6906_out0;
wire v$P15_6907_out0;
wire v$P15_6908_out0;
wire v$P16_6962_out0;
wire v$P16_6963_out0;
wire v$P16_6964_out0;
wire v$P16_6965_out0;
wire v$P16_6966_out0;
wire v$P17_11759_out0;
wire v$P17_11760_out0;
wire v$P17_11761_out0;
wire v$P17_11762_out0;
wire v$P17_11763_out0;
wire v$P18_11722_out0;
wire v$P18_11723_out0;
wire v$P18_11724_out0;
wire v$P18_11725_out0;
wire v$P18_11726_out0;
wire v$P19_16317_out0;
wire v$P19_16318_out0;
wire v$P19_16319_out0;
wire v$P19_16320_out0;
wire v$P19_16321_out0;
wire v$P1_2959_out0;
wire v$P1_2960_out0;
wire v$P1_2961_out0;
wire v$P1_2962_out0;
wire v$P1_2963_out0;
wire v$P20_10659_out0;
wire v$P20_10660_out0;
wire v$P20_10661_out0;
wire v$P20_10662_out0;
wire v$P20_10663_out0;
wire v$P21_4769_out0;
wire v$P21_4770_out0;
wire v$P21_4771_out0;
wire v$P21_4772_out0;
wire v$P21_4773_out0;
wire v$P22_4734_out0;
wire v$P22_4735_out0;
wire v$P22_4736_out0;
wire v$P22_4737_out0;
wire v$P22_4738_out0;
wire v$P23_6386_out0;
wire v$P23_6387_out0;
wire v$P23_6388_out0;
wire v$P23_6389_out0;
wire v$P23_6390_out0;
wire v$P2_2219_out0;
wire v$P2_2220_out0;
wire v$P2_2221_out0;
wire v$P2_2222_out0;
wire v$P2_2223_out0;
wire v$P3_15335_out0;
wire v$P3_15336_out0;
wire v$P3_15337_out0;
wire v$P3_15338_out0;
wire v$P3_15339_out0;
wire v$P4_13636_out0;
wire v$P4_13637_out0;
wire v$P4_13638_out0;
wire v$P4_13639_out0;
wire v$P4_13640_out0;
wire v$P5_221_out0;
wire v$P5_222_out0;
wire v$P5_223_out0;
wire v$P5_224_out0;
wire v$P5_225_out0;
wire v$P6_8104_out0;
wire v$P6_8105_out0;
wire v$P6_8106_out0;
wire v$P6_8107_out0;
wire v$P6_8108_out0;
wire v$P7_11769_out0;
wire v$P7_11770_out0;
wire v$P7_11771_out0;
wire v$P7_11772_out0;
wire v$P7_11773_out0;
wire v$P8_1703_out0;
wire v$P8_1704_out0;
wire v$P8_1705_out0;
wire v$P8_1706_out0;
wire v$P8_1707_out0;
wire v$P9_18445_out0;
wire v$P9_18446_out0;
wire v$P9_18447_out0;
wire v$P9_18448_out0;
wire v$P9_18449_out0;
wire v$PARITY_12073_out0;
wire v$PARITY_12074_out0;
wire v$PCHALTVIEWER_1768_out0;
wire v$PCHALT_12746_out0;
wire v$PCHALT_16563_out0;
wire v$PHALT0$PREV_7612_out0;
wire v$PHALT0_11638_out0;
wire v$PHALT1$PREV_7363_out0;
wire v$PHALT1_8934_out0;
wire v$PHALTVIEWER_2649_out0;
wire v$PHALT_15137_out0;
wire v$PHALT_1636_out0;
wire v$PHALT_17485_out0;
wire v$PIPELINE$RESTART_18625_out0;
wire v$PIPELINE$RESTART_18626_out0;
wire v$PIPELINE$RESTART_6071_out0;
wire v$PIPELINE$RESTART_6072_out0;
wire v$PIPELINEHALT_14816_out0;
wire v$PIPELINEHALT_14817_out0;
wire v$PIPELINERESTART_2418_out0;
wire v$PIPELINERESTART_2419_out0;
wire v$P_13868_out0;
wire v$P_13869_out0;
wire v$P_13870_out0;
wire v$P_13871_out0;
wire v$P_13872_out0;
wire v$P_13873_out0;
wire v$P_13874_out0;
wire v$P_13875_out0;
wire v$P_13876_out0;
wire v$P_13877_out0;
wire v$P_13878_out0;
wire v$P_13879_out0;
wire v$P_13880_out0;
wire v$P_13881_out0;
wire v$P_13882_out0;
wire v$P_13883_out0;
wire v$P_13884_out0;
wire v$P_13885_out0;
wire v$P_13886_out0;
wire v$P_13887_out0;
wire v$P_13888_out0;
wire v$P_13889_out0;
wire v$P_13890_out0;
wire v$P_13891_out0;
wire v$P_13892_out0;
wire v$P_13893_out0;
wire v$P_13894_out0;
wire v$P_13895_out0;
wire v$P_13896_out0;
wire v$P_13897_out0;
wire v$P_13898_out0;
wire v$P_13899_out0;
wire v$P_13900_out0;
wire v$P_13901_out0;
wire v$P_13902_out0;
wire v$P_13903_out0;
wire v$P_13904_out0;
wire v$P_13905_out0;
wire v$P_13906_out0;
wire v$P_13907_out0;
wire v$P_13908_out0;
wire v$P_13909_out0;
wire v$P_13910_out0;
wire v$P_13911_out0;
wire v$P_13912_out0;
wire v$P_13913_out0;
wire v$P_13914_out0;
wire v$P_13915_out0;
wire v$P_13916_out0;
wire v$P_13917_out0;
wire v$P_13918_out0;
wire v$P_13919_out0;
wire v$P_13920_out0;
wire v$P_13921_out0;
wire v$P_13922_out0;
wire v$P_13923_out0;
wire v$P_13924_out0;
wire v$P_13925_out0;
wire v$P_13926_out0;
wire v$P_13927_out0;
wire v$P_13928_out0;
wire v$P_13929_out0;
wire v$P_13930_out0;
wire v$P_13931_out0;
wire v$P_13932_out0;
wire v$P_13933_out0;
wire v$P_13934_out0;
wire v$P_13935_out0;
wire v$P_13936_out0;
wire v$P_13937_out0;
wire v$P_13938_out0;
wire v$P_13939_out0;
wire v$P_13940_out0;
wire v$P_13941_out0;
wire v$P_13942_out0;
wire v$P_13943_out0;
wire v$P_13944_out0;
wire v$P_13945_out0;
wire v$P_13946_out0;
wire v$P_13947_out0;
wire v$P_13948_out0;
wire v$P_13949_out0;
wire v$P_13950_out0;
wire v$P_13951_out0;
wire v$P_13952_out0;
wire v$P_13953_out0;
wire v$P_13954_out0;
wire v$P_13955_out0;
wire v$P_13956_out0;
wire v$P_13957_out0;
wire v$P_13958_out0;
wire v$P_13959_out0;
wire v$P_13960_out0;
wire v$P_13961_out0;
wire v$P_13962_out0;
wire v$P_13963_out0;
wire v$P_13964_out0;
wire v$P_13965_out0;
wire v$P_13966_out0;
wire v$P_13967_out0;
wire v$P_13968_out0;
wire v$P_13969_out0;
wire v$P_13970_out0;
wire v$P_13971_out0;
wire v$P_13972_out0;
wire v$P_13973_out0;
wire v$P_13974_out0;
wire v$P_13975_out0;
wire v$P_13976_out0;
wire v$P_13977_out0;
wire v$P_13978_out0;
wire v$P_13979_out0;
wire v$P_13980_out0;
wire v$P_13981_out0;
wire v$P_13982_out0;
wire v$P_13983_out0;
wire v$P_13984_out0;
wire v$P_13985_out0;
wire v$P_13986_out0;
wire v$P_13987_out0;
wire v$P_8310_out0;
wire v$P_8311_out0;
wire v$ParityCheck_16120_out0;
wire v$ParityCheck_16121_out0;
wire v$ParityEN_15784_out0;
wire v$ParityEN_15785_out0;
wire v$Q0P_12171_out0;
wire v$Q0P_12172_out0;
wire v$Q0P_16773_out0;
wire v$Q0P_16774_out0;
wire v$Q0_13703_out0;
wire v$Q0_13704_out0;
wire v$Q0_18318_out0;
wire v$Q0_18319_out0;
wire v$Q0_75_out0;
wire v$Q0_76_out0;
wire v$Q1P_11007_out0;
wire v$Q1P_11008_out0;
wire v$Q1P_5742_out0;
wire v$Q1P_5743_out0;
wire v$Q1_10923_out0;
wire v$Q1_10924_out0;
wire v$Q1_14326_out0;
wire v$Q1_14327_out0;
wire v$Q1_4450_out0;
wire v$Q1_4451_out0;
wire v$Q2P_4160_out0;
wire v$Q2P_4161_out0;
wire v$Q2P_6039_out0;
wire v$Q2P_6040_out0;
wire v$Q2_17486_out0;
wire v$Q2_17487_out0;
wire v$Q2_3149_out0;
wire v$Q2_3150_out0;
wire v$Q2_5457_out0;
wire v$Q2_5458_out0;
wire v$Q3P_11672_out0;
wire v$Q3P_11673_out0;
wire v$Q3P_13809_out0;
wire v$Q3P_13810_out0;
wire v$Q3_18289_out0;
wire v$Q3_18290_out0;
wire v$Q3_18425_out0;
wire v$Q3_18426_out0;
wire v$Q_14140_out0;
wire v$Q_14141_out0;
wire v$Q_14142_out0;
wire v$Q_14143_out0;
wire v$Q_14144_out0;
wire v$Q_14145_out0;
wire v$Q_14146_out0;
wire v$Q_14147_out0;
wire v$Q_14148_out0;
wire v$Q_14149_out0;
wire v$Q_14150_out0;
wire v$Q_14151_out0;
wire v$Q_14152_out0;
wire v$Q_14153_out0;
wire v$Q_14154_out0;
wire v$Q_14155_out0;
wire v$Q_14156_out0;
wire v$Q_14157_out0;
wire v$Q_14158_out0;
wire v$Q_14159_out0;
wire v$Q_14160_out0;
wire v$Q_14161_out0;
wire v$R0_15192_out0;
wire v$R0_15193_out0;
wire v$R0_2000_out0;
wire v$R0_6676_out0;
wire v$R1_11886_out0;
wire v$R1_15011_out0;
wire v$R1_15012_out0;
wire v$R1_17899_out0;
wire v$R2_3845_out0;
wire v$R2_3846_out0;
wire v$R3_15314_out0;
wire v$R3_15315_out0;
wire v$RAMWEN0_16569_out0;
wire v$RAMWEN1_10766_out0;
wire v$RAMWENVIEWER_17291_out0;
wire v$RAMWEN_15663_out0;
wire v$RAMWEN_15664_out0;
wire v$RAMWEN_17961_out0;
wire v$RAMWEN_7764_out0;
wire v$RAMWEN_7765_out0;
wire v$READ$REQUEST0_11394_out0;
wire v$READ$REQUEST0_18478_out0;
wire v$READ$REQUEST1_16828_out0;
wire v$READ$REQUEST1_6470_out0;
wire v$READ$REQUEST_14458_out0;
wire v$READ$REQUEST_14459_out0;
wire v$READ$REQUEST_16552_out0;
wire v$READ$REQUEST_16553_out0;
wire v$READ$REQUEST_7806_out0;
wire v$READ$REQUEST_7807_out0;
wire v$RECIEVEDPARITY_6224_out0;
wire v$RECIEVEDPARITY_6225_out0;
wire v$RR0VIEWER_14658_out0;
wire v$RR0_8089_out0;
wire v$RR1REGoutVIEWER_7381_out0;
wire v$RR1VIEWER_15032_out0;
wire v$RR1_1947_out0;
wire v$RXBIT_8913_out0;
wire v$RXBIT_8914_out0;
wire v$RXCLK_1240_out0;
wire v$RXCLK_1241_out0;
wire v$RXCLK_15844_out0;
wire v$RXCLK_15845_out0;
wire v$RXDISABLE_7888_out0;
wire v$RXDISABLE_7889_out0;
wire v$RXENABLE_3716_out0;
wire v$RXENABLE_3717_out0;
wire v$RXErrorSet_3480_out0;
wire v$RXErrorSet_3481_out0;
wire v$RXFLAG_12134_out0;
wire v$RXFLAG_12135_out0;
wire v$RXFLAG_15003_out0;
wire v$RXFLAG_15004_out0;
wire v$RXFlagSet_9108_out0;
wire v$RXFlagSet_9109_out0;
wire v$RXINTERRUPT_14845_out0;
wire v$RXINTERRUPT_14846_out0;
wire v$RXINTERRUPT_15347_out0;
wire v$RXINTERRUPT_15348_out0;
wire v$RXINT_12545_out0;
wire v$RXINT_12546_out0;
wire v$RXREAD_15344_out0;
wire v$RXREAD_15345_out0;
wire v$RXREAD_15854_out0;
wire v$RXREAD_15855_out0;
wire v$RXRead_16365_out0;
wire v$RXRead_16366_out0;
wire v$RXRegAdd_12974_out0;
wire v$RXRegAdd_12975_out0;
wire v$RXReset_16530_out0;
wire v$RXReset_16531_out0;
wire v$RXSET_14687_out0;
wire v$RXSET_14688_out0;
wire v$RXSHIFT_674_out0;
wire v$RXSHIFT_675_out0;
wire v$RX_2966_out0;
wire v$RX_2967_out0;
wire v$RX_43_out0;
wire v$RX_44_out0;
wire v$RX_4808_out0;
wire v$RX_4809_out0;
wire v$RX_6186_out0;
wire v$RX_6187_out0;
wire v$RX_6652_out0;
wire v$RX_6653_out0;
wire v$RXflag_15841_out0;
wire v$RXflag_15842_out0;
wire v$RXlast_12821_out0;
wire v$RXlast_12822_out0;
wire v$RXoverflow_9540_out0;
wire v$RXoverflow_9541_out0;
wire v$RXreset_5959_out0;
wire v$RXreset_5960_out0;
wire v$RXset_1701_out0;
wire v$RXset_1702_out0;
wire v$RXset_5101_out0;
wire v$RXset_5102_out0;
wire v$R_1487_out0;
wire v$R_1488_out0;
wire v$R_1489_out0;
wire v$R_1490_out0;
wire v$R_1586_out0;
wire v$R_1587_out0;
wire v$R_1588_out0;
wire v$R_1589_out0;
wire v$R_1590_out0;
wire v$R_16745_out0;
wire v$R_18331_out0;
wire v$R_18332_out0;
wire v$R_18333_out0;
wire v$R_18334_out0;
wire v$R_18335_out0;
wire v$R_18336_out0;
wire v$R_18337_out0;
wire v$R_18338_out0;
wire v$R_18339_out0;
wire v$R_18340_out0;
wire v$R_18341_out0;
wire v$R_18342_out0;
wire v$R_18343_out0;
wire v$R_18344_out0;
wire v$R_18345_out0;
wire v$R_18346_out0;
wire v$R_18347_out0;
wire v$R_18348_out0;
wire v$R_18349_out0;
wire v$R_18350_out0;
wire v$R_18351_out0;
wire v$R_18352_out0;
wire v$R_8778_out0;
wire v$R_8779_out0;
wire v$RceivedParity_18539_out0;
wire v$RceivedParity_18540_out0;
wire v$RecievedParity_9538_out0;
wire v$RecievedParity_9539_out0;
wire v$SAME$H_1156_out0;
wire v$SAME$H_1157_out0;
wire v$SAME$H_8915_out0;
wire v$SAME$H_8916_out0;
wire v$SAME$L_16440_out0;
wire v$SAME$L_16441_out0;
wire v$SAME$L_9463_out0;
wire v$SAME$L_9464_out0;
wire v$SAME_18363_out0;
wire v$SAME_18364_out0;
wire v$SAME_18365_out0;
wire v$SAME_18366_out0;
wire v$SAME_18367_out0;
wire v$SAME_18368_out0;
wire v$SAME_18369_out0;
wire v$SAME_18370_out0;
wire v$SAME_18723_out0;
wire v$SAME_18724_out0;
wire v$SAME_18725_out0;
wire v$SAME_18726_out0;
wire v$SAME_18727_out0;
wire v$SAME_18728_out0;
wire v$SAME_18729_out0;
wire v$SAME_18730_out0;
wire v$SAME_18731_out0;
wire v$SAME_18732_out0;
wire v$SAME_18733_out0;
wire v$SAME_18734_out0;
wire v$SAME_18735_out0;
wire v$SAME_18736_out0;
wire v$SAME_18737_out0;
wire v$SAME_18738_out0;
wire v$SAME_18739_out0;
wire v$SAME_18740_out0;
wire v$SAME_18741_out0;
wire v$SAME_18742_out0;
wire v$SAME_18743_out0;
wire v$SAME_18744_out0;
wire v$SAME_18745_out0;
wire v$SAME_18746_out0;
wire v$SAME_18747_out0;
wire v$SAME_18748_out0;
wire v$SAME_18749_out0;
wire v$SAME_18750_out0;
wire v$SAME_18751_out0;
wire v$SAME_18752_out0;
wire v$SAME_18753_out0;
wire v$SAME_18754_out0;
wire v$SAME_6264_out0;
wire v$SAME_6265_out0;
wire v$SAME_8919_out0;
wire v$SAME_8920_out0;
wire v$SAME_8921_out0;
wire v$SAME_8922_out0;
wire v$SAVES$TO$REG_12526_out0;
wire v$SEL10_12606_out0;
wire v$SEL10_12607_out0;
wire v$SEL10_12608_out0;
wire v$SEL10_12609_out0;
wire v$SEL10_12610_out0;
wire v$SEL10_12611_out0;
wire v$SEL10_12612_out0;
wire v$SEL10_12613_out0;
wire v$SEL10_12614_out0;
wire v$SEL10_12615_out0;
wire v$SEL10_12616_out0;
wire v$SEL10_12617_out0;
wire v$SEL10_12618_out0;
wire v$SEL10_12619_out0;
wire v$SEL10_12620_out0;
wire v$SEL10_12621_out0;
wire v$SEL10_12622_out0;
wire v$SEL10_12623_out0;
wire v$SEL10_12624_out0;
wire v$SEL10_12625_out0;
wire v$SEL10_12626_out0;
wire v$SEL10_12627_out0;
wire v$SEL10_12628_out0;
wire v$SEL10_12629_out0;
wire v$SEL10_1815_out0;
wire v$SEL10_4152_out0;
wire v$SEL10_4153_out0;
wire v$SEL10_7279_out0;
wire v$SEL10_7280_out0;
wire v$SEL10_9506_out0;
wire v$SEL10_9507_out0;
wire v$SEL10_9508_out0;
wire v$SEL10_9509_out0;
wire v$SEL11_12201_out0;
wire v$SEL11_12202_out0;
wire v$SEL11_1500_out0;
wire v$SEL11_15556_out0;
wire v$SEL11_15557_out0;
wire v$SEL11_15890_out0;
wire v$SEL11_15891_out0;
wire v$SEL11_7225_out0;
wire v$SEL11_7226_out0;
wire v$SEL11_7227_out0;
wire v$SEL11_7228_out0;
wire v$SEL11_8352_out0;
wire v$SEL11_8353_out0;
wire v$SEL12_1351_out0;
wire v$SEL12_1352_out0;
wire v$SEL12_13844_out0;
wire v$SEL12_13845_out0;
wire v$SEL12_13846_out0;
wire v$SEL12_13847_out0;
wire v$SEL12_1516_out0;
wire v$SEL13_13249_out0;
wire v$SEL13_14655_out0;
wire v$SEL13_17581_out0;
wire v$SEL13_17582_out0;
wire v$SEL13_3883_out0;
wire v$SEL13_6924_out0;
wire v$SEL13_6925_out0;
wire v$SEL13_6926_out0;
wire v$SEL13_6927_out0;
wire v$SEL14_16347_out0;
wire v$SEL14_16348_out0;
wire v$SEL14_16349_out0;
wire v$SEL14_16350_out0;
wire v$SEL14_4815_out0;
wire v$SEL15_13612_out0;
wire v$SEL15_13613_out0;
wire v$SEL15_4886_out0;
wire v$SEL15_4887_out0;
wire v$SEL15_4888_out0;
wire v$SEL15_4889_out0;
wire v$SEL15_9438_out0;
wire v$SEL16_16894_out0;
wire v$SEL16_16895_out0;
wire v$SEL16_16896_out0;
wire v$SEL16_16897_out0;
wire v$SEL17_16069_out0;
wire v$SEL17_16070_out0;
wire v$SEL17_16071_out0;
wire v$SEL17_16072_out0;
wire v$SEL18_11379_out0;
wire v$SEL18_11380_out0;
wire v$SEL18_11381_out0;
wire v$SEL18_11382_out0;
wire v$SEL19_12815_out0;
wire v$SEL19_12816_out0;
wire v$SEL19_12817_out0;
wire v$SEL19_12818_out0;
wire v$SEL1_11087_out0;
wire v$SEL1_11088_out0;
wire v$SEL1_11089_out0;
wire v$SEL1_11090_out0;
wire v$SEL1_11091_out0;
wire v$SEL1_11092_out0;
wire v$SEL1_11093_out0;
wire v$SEL1_11094_out0;
wire v$SEL1_11095_out0;
wire v$SEL1_11096_out0;
wire v$SEL1_11097_out0;
wire v$SEL1_11098_out0;
wire v$SEL1_1280_out0;
wire v$SEL1_13355_out0;
wire v$SEL1_13356_out0;
wire v$SEL1_13357_out0;
wire v$SEL1_13358_out0;
wire v$SEL1_13459_out0;
wire v$SEL1_13460_out0;
wire v$SEL1_13461_out0;
wire v$SEL1_13462_out0;
wire v$SEL1_13463_out0;
wire v$SEL1_13464_out0;
wire v$SEL1_13465_out0;
wire v$SEL1_13466_out0;
wire v$SEL1_13467_out0;
wire v$SEL1_13468_out0;
wire v$SEL1_13469_out0;
wire v$SEL1_13470_out0;
wire v$SEL1_13471_out0;
wire v$SEL1_13472_out0;
wire v$SEL1_13473_out0;
wire v$SEL1_13474_out0;
wire v$SEL1_13475_out0;
wire v$SEL1_13476_out0;
wire v$SEL1_13477_out0;
wire v$SEL1_13478_out0;
wire v$SEL1_13479_out0;
wire v$SEL1_13480_out0;
wire v$SEL1_13481_out0;
wire v$SEL1_13482_out0;
wire v$SEL1_13483_out0;
wire v$SEL1_13484_out0;
wire v$SEL1_13485_out0;
wire v$SEL1_13486_out0;
wire v$SEL1_13487_out0;
wire v$SEL1_13488_out0;
wire v$SEL1_13489_out0;
wire v$SEL1_13490_out0;
wire v$SEL1_13491_out0;
wire v$SEL1_13492_out0;
wire v$SEL1_13493_out0;
wire v$SEL1_13494_out0;
wire v$SEL1_13495_out0;
wire v$SEL1_13496_out0;
wire v$SEL1_13497_out0;
wire v$SEL1_13498_out0;
wire v$SEL1_13499_out0;
wire v$SEL1_13500_out0;
wire v$SEL1_13501_out0;
wire v$SEL1_13502_out0;
wire v$SEL1_13503_out0;
wire v$SEL1_13504_out0;
wire v$SEL1_13505_out0;
wire v$SEL1_13506_out0;
wire v$SEL1_18044_out0;
wire v$SEL1_18045_out0;
wire v$SEL1_18046_out0;
wire v$SEL1_18047_out0;
wire v$SEL1_2269_out0;
wire v$SEL1_2270_out0;
wire v$SEL1_2271_out0;
wire v$SEL1_2272_out0;
wire v$SEL1_2273_out0;
wire v$SEL1_2274_out0;
wire v$SEL1_2275_out0;
wire v$SEL1_2276_out0;
wire v$SEL1_3515_out0;
wire v$SEL1_3720_out0;
wire v$SEL1_3721_out0;
wire v$SEL1_7005_out0;
wire v$SEL1_7088_out0;
wire v$SEL1_7089_out0;
wire v$SEL1_7090_out0;
wire v$SEL1_7091_out0;
wire v$SEL20_8174_out0;
wire v$SEL20_8175_out0;
wire v$SEL20_8176_out0;
wire v$SEL20_8177_out0;
wire v$SEL21_11048_out0;
wire v$SEL21_11049_out0;
wire v$SEL21_11050_out0;
wire v$SEL21_11051_out0;
wire v$SEL22_7397_out0;
wire v$SEL22_7398_out0;
wire v$SEL22_7399_out0;
wire v$SEL22_7400_out0;
wire v$SEL23_7617_out0;
wire v$SEL23_7618_out0;
wire v$SEL23_7619_out0;
wire v$SEL23_7620_out0;
wire v$SEL24_16922_out0;
wire v$SEL24_16923_out0;
wire v$SEL24_16924_out0;
wire v$SEL24_16925_out0;
wire v$SEL27_16304_out0;
wire v$SEL27_16305_out0;
wire v$SEL27_16306_out0;
wire v$SEL27_16307_out0;
wire v$SEL28_7327_out0;
wire v$SEL28_7328_out0;
wire v$SEL28_7329_out0;
wire v$SEL28_7330_out0;
wire v$SEL29_16594_out0;
wire v$SEL29_16595_out0;
wire v$SEL29_16596_out0;
wire v$SEL29_16597_out0;
wire v$SEL2_11607_out0;
wire v$SEL2_11608_out0;
wire v$SEL2_11609_out0;
wire v$SEL2_11610_out0;
wire v$SEL2_11611_out0;
wire v$SEL2_11612_out0;
wire v$SEL2_11613_out0;
wire v$SEL2_11614_out0;
wire v$SEL2_11615_out0;
wire v$SEL2_11616_out0;
wire v$SEL2_11617_out0;
wire v$SEL2_13321_out0;
wire v$SEL2_13322_out0;
wire v$SEL2_13323_out0;
wire v$SEL2_13324_out0;
wire v$SEL2_13433_out0;
wire v$SEL2_13434_out0;
wire v$SEL2_14411_out0;
wire v$SEL2_15836_out0;
wire v$SEL2_16600_out0;
wire v$SEL2_16601_out0;
wire v$SEL2_16602_out0;
wire v$SEL2_16603_out0;
wire v$SEL2_16604_out0;
wire v$SEL2_16605_out0;
wire v$SEL2_16606_out0;
wire v$SEL2_16607_out0;
wire v$SEL2_16608_out0;
wire v$SEL2_16609_out0;
wire v$SEL2_16610_out0;
wire v$SEL2_16611_out0;
wire v$SEL2_16612_out0;
wire v$SEL2_16613_out0;
wire v$SEL2_16614_out0;
wire v$SEL2_16615_out0;
wire v$SEL2_16616_out0;
wire v$SEL2_16617_out0;
wire v$SEL2_16618_out0;
wire v$SEL2_16619_out0;
wire v$SEL2_16620_out0;
wire v$SEL2_16621_out0;
wire v$SEL2_16622_out0;
wire v$SEL2_16623_out0;
wire v$SEL2_18355_out0;
wire v$SEL2_18356_out0;
wire v$SEL2_18357_out0;
wire v$SEL2_18358_out0;
wire v$SEL2_18359_out0;
wire v$SEL2_18360_out0;
wire v$SEL2_18361_out0;
wire v$SEL2_18362_out0;
wire v$SEL2_18502_out0;
wire v$SEL2_18503_out0;
wire v$SEL2_18504_out0;
wire v$SEL2_18505_out0;
wire v$SEL2_3714_out0;
wire v$SEL2_3715_out0;
wire v$SEL2_7670_out0;
wire v$SEL2_7671_out0;
wire v$SEL2_7672_out0;
wire v$SEL2_7673_out0;
wire v$SEL2_7674_out0;
wire v$SEL2_7675_out0;
wire v$SEL2_7676_out0;
wire v$SEL2_7677_out0;
wire v$SEL2_7678_out0;
wire v$SEL2_7679_out0;
wire v$SEL2_7680_out0;
wire v$SEL2_7681_out0;
wire v$SEL2_7682_out0;
wire v$SEL2_7683_out0;
wire v$SEL2_7684_out0;
wire v$SEL2_7685_out0;
wire v$SEL2_7686_out0;
wire v$SEL2_7687_out0;
wire v$SEL2_7688_out0;
wire v$SEL2_7689_out0;
wire v$SEL2_7690_out0;
wire v$SEL2_7691_out0;
wire v$SEL2_7692_out0;
wire v$SEL2_7693_out0;
wire v$SEL2_7694_out0;
wire v$SEL2_7695_out0;
wire v$SEL2_7696_out0;
wire v$SEL2_7697_out0;
wire v$SEL2_7698_out0;
wire v$SEL2_7699_out0;
wire v$SEL2_7700_out0;
wire v$SEL2_7701_out0;
wire v$SEL2_7702_out0;
wire v$SEL2_7703_out0;
wire v$SEL2_7704_out0;
wire v$SEL2_7705_out0;
wire v$SEL2_7706_out0;
wire v$SEL2_7707_out0;
wire v$SEL2_7708_out0;
wire v$SEL2_7709_out0;
wire v$SEL2_7710_out0;
wire v$SEL2_7711_out0;
wire v$SEL2_7712_out0;
wire v$SEL2_7713_out0;
wire v$SEL2_7714_out0;
wire v$SEL2_7715_out0;
wire v$SEL2_7716_out0;
wire v$SEL2_7717_out0;
wire v$SEL2_9428_out0;
wire v$SEL2_9429_out0;
wire v$SEL3_1137_out0;
wire v$SEL3_1138_out0;
wire v$SEL3_1139_out0;
wire v$SEL3_1140_out0;
wire v$SEL3_1141_out0;
wire v$SEL3_1142_out0;
wire v$SEL3_1143_out0;
wire v$SEL3_1144_out0;
wire v$SEL3_11729_out0;
wire v$SEL3_11730_out0;
wire v$SEL3_11731_out0;
wire v$SEL3_11732_out0;
wire v$SEL3_14006_out0;
wire v$SEL3_14007_out0;
wire v$SEL3_14008_out0;
wire v$SEL3_14009_out0;
wire v$SEL3_1698_out0;
wire v$SEL3_17400_out0;
wire v$SEL3_17401_out0;
wire v$SEL3_18659_out0;
wire v$SEL3_2294_out0;
wire v$SEL3_2295_out0;
wire v$SEL3_2296_out0;
wire v$SEL3_2297_out0;
wire v$SEL3_2298_out0;
wire v$SEL3_2299_out0;
wire v$SEL3_2300_out0;
wire v$SEL3_2301_out0;
wire v$SEL3_2302_out0;
wire v$SEL3_2303_out0;
wire v$SEL3_2304_out0;
wire v$SEL3_2305_out0;
wire v$SEL3_2306_out0;
wire v$SEL3_2307_out0;
wire v$SEL3_2308_out0;
wire v$SEL3_2309_out0;
wire v$SEL3_2310_out0;
wire v$SEL3_2311_out0;
wire v$SEL3_2312_out0;
wire v$SEL3_2313_out0;
wire v$SEL3_2314_out0;
wire v$SEL3_2315_out0;
wire v$SEL3_2316_out0;
wire v$SEL3_2317_out0;
wire v$SEL3_2318_out0;
wire v$SEL3_2319_out0;
wire v$SEL3_2320_out0;
wire v$SEL3_2321_out0;
wire v$SEL3_2322_out0;
wire v$SEL3_2323_out0;
wire v$SEL3_2324_out0;
wire v$SEL3_2325_out0;
wire v$SEL3_2326_out0;
wire v$SEL3_2327_out0;
wire v$SEL3_2328_out0;
wire v$SEL3_2329_out0;
wire v$SEL3_2330_out0;
wire v$SEL3_2331_out0;
wire v$SEL3_2332_out0;
wire v$SEL3_2333_out0;
wire v$SEL3_2334_out0;
wire v$SEL3_2335_out0;
wire v$SEL3_2336_out0;
wire v$SEL3_2337_out0;
wire v$SEL3_2338_out0;
wire v$SEL3_2339_out0;
wire v$SEL3_2340_out0;
wire v$SEL3_2341_out0;
wire v$SEL3_3126_out0;
wire v$SEL3_8424_out0;
wire v$SEL3_8425_out0;
wire v$SEL3_8426_out0;
wire v$SEL3_8427_out0;
wire v$SEL3_8428_out0;
wire v$SEL3_8429_out0;
wire v$SEL3_8430_out0;
wire v$SEL3_8431_out0;
wire v$SEL3_8432_out0;
wire v$SEL3_8433_out0;
wire v$SEL3_8434_out0;
wire v$SEL3_8435_out0;
wire v$SEL3_8436_out0;
wire v$SEL3_8437_out0;
wire v$SEL3_8438_out0;
wire v$SEL3_8439_out0;
wire v$SEL3_8440_out0;
wire v$SEL3_8441_out0;
wire v$SEL3_8442_out0;
wire v$SEL3_8443_out0;
wire v$SEL3_8444_out0;
wire v$SEL3_8445_out0;
wire v$SEL3_8446_out0;
wire v$SEL3_8447_out0;
wire v$SEL4_1186_out0;
wire v$SEL4_16422_out0;
wire v$SEL4_1845_out0;
wire v$SEL4_1846_out0;
wire v$SEL4_1847_out0;
wire v$SEL4_1848_out0;
wire v$SEL4_4937_out0;
wire v$SEL4_4938_out0;
wire v$SEL4_4939_out0;
wire v$SEL4_4940_out0;
wire v$SEL4_4941_out0;
wire v$SEL4_4942_out0;
wire v$SEL4_4943_out0;
wire v$SEL4_4944_out0;
wire v$SEL4_6079_out0;
wire v$SEL4_6080_out0;
wire v$SEL4_6081_out0;
wire v$SEL4_6082_out0;
wire v$SEL4_6083_out0;
wire v$SEL4_6084_out0;
wire v$SEL4_6085_out0;
wire v$SEL4_6086_out0;
wire v$SEL4_6087_out0;
wire v$SEL4_6088_out0;
wire v$SEL4_6089_out0;
wire v$SEL4_6090_out0;
wire v$SEL4_6091_out0;
wire v$SEL4_6092_out0;
wire v$SEL4_6093_out0;
wire v$SEL4_6094_out0;
wire v$SEL4_6095_out0;
wire v$SEL4_6096_out0;
wire v$SEL4_6097_out0;
wire v$SEL4_6098_out0;
wire v$SEL4_6099_out0;
wire v$SEL4_6100_out0;
wire v$SEL4_6101_out0;
wire v$SEL4_6102_out0;
wire v$SEL4_6103_out0;
wire v$SEL4_6104_out0;
wire v$SEL4_6105_out0;
wire v$SEL4_6106_out0;
wire v$SEL4_6107_out0;
wire v$SEL4_6108_out0;
wire v$SEL4_6109_out0;
wire v$SEL4_6110_out0;
wire v$SEL4_6111_out0;
wire v$SEL4_6112_out0;
wire v$SEL4_6113_out0;
wire v$SEL4_6114_out0;
wire v$SEL4_6115_out0;
wire v$SEL4_6116_out0;
wire v$SEL4_6117_out0;
wire v$SEL4_6118_out0;
wire v$SEL4_6119_out0;
wire v$SEL4_6120_out0;
wire v$SEL4_6121_out0;
wire v$SEL4_6122_out0;
wire v$SEL4_6123_out0;
wire v$SEL4_6124_out0;
wire v$SEL4_6125_out0;
wire v$SEL4_6126_out0;
wire v$SEL4_7053_out0;
wire v$SEL4_7054_out0;
wire v$SEL4_7321_out0;
wire v$SEL4_7322_out0;
wire v$SEL4_7323_out0;
wire v$SEL4_7324_out0;
wire v$SEL4_7334_out0;
wire v$SEL4_7335_out0;
wire v$SEL4_7336_out0;
wire v$SEL4_7337_out0;
wire v$SEL4_7338_out0;
wire v$SEL4_7339_out0;
wire v$SEL4_7340_out0;
wire v$SEL4_7341_out0;
wire v$SEL4_7342_out0;
wire v$SEL4_7343_out0;
wire v$SEL4_7344_out0;
wire v$SEL4_7345_out0;
wire v$SEL4_7346_out0;
wire v$SEL4_7347_out0;
wire v$SEL4_7348_out0;
wire v$SEL4_7349_out0;
wire v$SEL4_7350_out0;
wire v$SEL4_7351_out0;
wire v$SEL4_7352_out0;
wire v$SEL4_7353_out0;
wire v$SEL4_7354_out0;
wire v$SEL4_7355_out0;
wire v$SEL4_7356_out0;
wire v$SEL4_7357_out0;
wire v$SEL5_11625_out0;
wire v$SEL5_11667_out0;
wire v$SEL5_11668_out0;
wire v$SEL5_11669_out0;
wire v$SEL5_11670_out0;
wire v$SEL5_12215_out0;
wire v$SEL5_12216_out0;
wire v$SEL5_12217_out0;
wire v$SEL5_12218_out0;
wire v$SEL5_12219_out0;
wire v$SEL5_12220_out0;
wire v$SEL5_12221_out0;
wire v$SEL5_12222_out0;
wire v$SEL5_12776_out0;
wire v$SEL5_12777_out0;
wire v$SEL5_12778_out0;
wire v$SEL5_12779_out0;
wire v$SEL5_12780_out0;
wire v$SEL5_12781_out0;
wire v$SEL5_12782_out0;
wire v$SEL5_12783_out0;
wire v$SEL5_12784_out0;
wire v$SEL5_12785_out0;
wire v$SEL5_12786_out0;
wire v$SEL5_12787_out0;
wire v$SEL5_12788_out0;
wire v$SEL5_12789_out0;
wire v$SEL5_12790_out0;
wire v$SEL5_12791_out0;
wire v$SEL5_12792_out0;
wire v$SEL5_12793_out0;
wire v$SEL5_12794_out0;
wire v$SEL5_12795_out0;
wire v$SEL5_12796_out0;
wire v$SEL5_12797_out0;
wire v$SEL5_12798_out0;
wire v$SEL5_12799_out0;
wire v$SEL5_15451_out0;
wire v$SEL5_15452_out0;
wire v$SEL5_15453_out0;
wire v$SEL5_15454_out0;
wire v$SEL5_1581_out0;
wire v$SEL5_313_out0;
wire v$SEL5_314_out0;
wire v$SEL6_12472_out0;
wire v$SEL6_12473_out0;
wire v$SEL6_12474_out0;
wire v$SEL6_12475_out0;
wire v$SEL6_13779_out0;
wire v$SEL6_13780_out0;
wire v$SEL6_13781_out0;
wire v$SEL6_13782_out0;
wire v$SEL6_13783_out0;
wire v$SEL6_13784_out0;
wire v$SEL6_13785_out0;
wire v$SEL6_13786_out0;
wire v$SEL6_14244_out0;
wire v$SEL6_14456_out0;
wire v$SEL6_14457_out0;
wire v$SEL6_5805_out0;
wire v$SEL6_5806_out0;
wire v$SEL6_5807_out0;
wire v$SEL6_5808_out0;
wire v$SEL6_8932_out0;
wire v$SEL6_8933_out0;
wire v$SEL7_1223_out0;
wire v$SEL7_14332_out0;
wire v$SEL7_14333_out0;
wire v$SEL7_14334_out0;
wire v$SEL7_14335_out0;
wire v$SEL7_15615_out0;
wire v$SEL7_15616_out0;
wire v$SEL7_17010_out0;
wire v$SEL7_4166_out0;
wire v$SEL7_4167_out0;
wire v$SEL7_4168_out0;
wire v$SEL7_4169_out0;
wire v$SEL7_4170_out0;
wire v$SEL7_4171_out0;
wire v$SEL7_4172_out0;
wire v$SEL7_4173_out0;
wire v$SEL7_4174_out0;
wire v$SEL7_4175_out0;
wire v$SEL7_4176_out0;
wire v$SEL7_4177_out0;
wire v$SEL7_4178_out0;
wire v$SEL7_4179_out0;
wire v$SEL7_4180_out0;
wire v$SEL7_4181_out0;
wire v$SEL7_4182_out0;
wire v$SEL7_4183_out0;
wire v$SEL7_4184_out0;
wire v$SEL7_4185_out0;
wire v$SEL7_4186_out0;
wire v$SEL7_4187_out0;
wire v$SEL7_4188_out0;
wire v$SEL7_4189_out0;
wire v$SEL7_6345_out0;
wire v$SEL7_6346_out0;
wire v$SEL7_6347_out0;
wire v$SEL7_6348_out0;
wire v$SEL7_6349_out0;
wire v$SEL7_6350_out0;
wire v$SEL7_6351_out0;
wire v$SEL7_6352_out0;
wire v$SEL8_12914_out0;
wire v$SEL8_12915_out0;
wire v$SEL8_12916_out0;
wire v$SEL8_12917_out0;
wire v$SEL8_12918_out0;
wire v$SEL8_12919_out0;
wire v$SEL8_12920_out0;
wire v$SEL8_12921_out0;
wire v$SEL8_12922_out0;
wire v$SEL8_12923_out0;
wire v$SEL8_12924_out0;
wire v$SEL8_12925_out0;
wire v$SEL8_12926_out0;
wire v$SEL8_12927_out0;
wire v$SEL8_12928_out0;
wire v$SEL8_12929_out0;
wire v$SEL8_12930_out0;
wire v$SEL8_12931_out0;
wire v$SEL8_12932_out0;
wire v$SEL8_12933_out0;
wire v$SEL8_12934_out0;
wire v$SEL8_12935_out0;
wire v$SEL8_12936_out0;
wire v$SEL8_12937_out0;
wire v$SEL8_16570_out0;
wire v$SEL8_16571_out0;
wire v$SEL8_16572_out0;
wire v$SEL8_16573_out0;
wire v$SEL8_16574_out0;
wire v$SEL8_16575_out0;
wire v$SEL8_16576_out0;
wire v$SEL8_16577_out0;
wire v$SEL8_17683_out0;
wire v$SEL8_17684_out0;
wire v$SEL8_17685_out0;
wire v$SEL8_17686_out0;
wire v$SEL8_1968_out0;
wire v$SEL9_10263_out0;
wire v$SEL9_10264_out0;
wire v$SEL9_10265_out0;
wire v$SEL9_10266_out0;
wire v$SEL9_10837_out0;
wire v$SEL9_10838_out0;
wire v$SEL9_10839_out0;
wire v$SEL9_10840_out0;
wire v$SEL9_10841_out0;
wire v$SEL9_10842_out0;
wire v$SEL9_10843_out0;
wire v$SEL9_10844_out0;
wire v$SEL9_10845_out0;
wire v$SEL9_10846_out0;
wire v$SEL9_10847_out0;
wire v$SEL9_10848_out0;
wire v$SEL9_10849_out0;
wire v$SEL9_10850_out0;
wire v$SEL9_10851_out0;
wire v$SEL9_10852_out0;
wire v$SEL9_10853_out0;
wire v$SEL9_10854_out0;
wire v$SEL9_10855_out0;
wire v$SEL9_10856_out0;
wire v$SEL9_10857_out0;
wire v$SEL9_10858_out0;
wire v$SEL9_10859_out0;
wire v$SEL9_10860_out0;
wire v$SEL9_5394_out0;
wire v$SELIN$VIEWER_11070_out0;
wire v$SELIN_18215_out0;
wire v$SELOUTVIEWER_7278_out0;
wire v$SELOUT_1720_out0;
wire v$SERIALIN_5728_out0;
wire v$SERIALIN_5729_out0;
wire v$SHIFTEN_10282_out0;
wire v$SHIFTEN_10283_out0;
wire v$SHIFTEN_12766_out0;
wire v$SHIFTEN_12767_out0;
wire v$SHIFTEN_7092_out0;
wire v$SHIFTEN_7093_out0;
wire v$SHIFTEN_9406_out0;
wire v$SHIFTEN_9407_out0;
wire v$SHIFTEN_9408_out0;
wire v$SHIFTEN_9409_out0;
wire v$SHIFTEN_9410_out0;
wire v$SHIFTEN_9411_out0;
wire v$SHIFTEN_9412_out0;
wire v$SHIFTEN_9413_out0;
wire v$SHIFTEN_9414_out0;
wire v$SHIFTEN_9415_out0;
wire v$SHIFTEN_9416_out0;
wire v$SHIFTEN_9417_out0;
wire v$SHOULD$STORE_12710_out0;
wire v$SIGN_12760_out0;
wire v$SIGN_12761_out0;
wire v$SIGN_1366_out0;
wire v$SIGN_1367_out0;
wire v$SIGN_1368_out0;
wire v$SIGN_1369_out0;
wire v$SIN_100_out0;
wire v$SIN_101_out0;
wire v$SIN_102_out0;
wire v$SIN_91_out0;
wire v$SIN_92_out0;
wire v$SIN_93_out0;
wire v$SIN_94_out0;
wire v$SIN_95_out0;
wire v$SIN_96_out0;
wire v$SIN_97_out0;
wire v$SIN_98_out0;
wire v$SIN_99_out0;
wire v$SOUT1_1917_out0;
wire v$SOUT1_1918_out0;
wire v$SOUT1_1919_out0;
wire v$SOUT1_1920_out0;
wire v$SOUT1_1921_out0;
wire v$SOUT1_1922_out0;
wire v$SOUT1_1923_out0;
wire v$SOUT1_1924_out0;
wire v$SOUT1_1925_out0;
wire v$SOUT1_1926_out0;
wire v$SOUT1_1927_out0;
wire v$SOUT1_1928_out0;
wire v$SOUT_18193_out0;
wire v$SOUT_18194_out0;
wire v$STALL$FETCH$OCCURRED_2647_out0;
wire v$STALL$FETCH$OCCURRED_2648_out0;
wire v$STALL$IN$PREV_13214_out0;
wire v$STALL$IN$PREV_13215_out0;
wire v$STALL$PREV$CYCLE_5772_out0;
wire v$STALL$PREV$CYCLE_5773_out0;
wire v$STALL$PREV$PREV_5809_out0;
wire v$STALL$PREV$PREV_5810_out0;
wire v$STALL$VIEWER_18065_out0;
wire v$STALL$VIEWER_18066_out0;
wire v$STALL_12230_out0;
wire v$STALL_12231_out0;
wire v$STALL_13145_out0;
wire v$STALL_13146_out0;
wire v$STALL_15494_out0;
wire v$STALL_15495_out0;
wire v$STALL_17890_out0;
wire v$STALL_17891_out0;
wire v$START$PIPELINED$VIEWER_6398_out0;
wire v$START_14012_out0;
wire v$START_16352_out0;
wire v$START_18718_out0;
wire v$START_3700_out0;
wire v$START_4238_out0;
wire v$START_5492_out0;
wire v$STATE_16013_out0;
wire v$STATE_16014_out0;
wire v$STATE_16015_out0;
wire v$STATE_16016_out0;
wire v$STATE_16017_out0;
wire v$STATUSCLR_5953_out0;
wire v$STATUSCLR_5954_out0;
wire v$STATUSREAD_1637_out0;
wire v$STATUSREAD_1638_out0;
wire v$STClr_10217_out0;
wire v$STClr_10218_out0;
wire v$STOP$1_7810_out0;
wire v$STOP$1_7811_out0;
wire v$STOP$2_8234_out0;
wire v$STOP$2_8235_out0;
wire v$STOPBITERROR_11727_out0;
wire v$STOPBITERROR_11728_out0;
wire v$STOPERROR_294_out0;
wire v$STOPERROR_295_out0;
wire v$STP$DECODED_16534_out0;
wire v$STP$DECODED_16535_out0;
wire v$STP$SAVED_7560_out0;
wire v$STP$SAVED_7561_out0;
wire v$STPHALT_12943_out0;
wire v$STPHALT_12944_out0;
wire v$STPHALT_18124_out0;
wire v$STPHALT_18125_out0;
wire v$STPHALT_4317_out0;
wire v$STPHALT_4318_out0;
wire v$STP_10818_out0;
wire v$STP_10819_out0;
wire v$STP_11714_out0;
wire v$STP_11715_out0;
wire v$STP_17762_out0;
wire v$STP_17763_out0;
wire v$STP_6205_out0;
wire v$STP_6206_out0;
wire v$STRead_9925_out0;
wire v$STRead_9926_out0;
wire v$SUBEN_12858_out0;
wire v$SUBEN_12859_out0;
wire v$SUBTRACTION$SIGN_11872_out0;
wire v$SUBTRACTION$SIGN_11873_out0;
wire v$SUB_13790_out0;
wire v$SUB_13791_out0;
wire v$SUM$0_12330_out0;
wire v$SUM$10_14308_out0;
wire v$SUM$11_17033_out0;
wire v$SUM$1_10360_out0;
wire v$SUM$2_9082_out0;
wire v$SUM$3_7904_out0;
wire v$SUM$4_15246_out0;
wire v$SUM$5_7817_out0;
wire v$SUM$6_12912_out0;
wire v$SUM$7_7743_out0;
wire v$SUM$8_15776_out0;
wire v$SUM$9_197_out0;
wire v$S_10347_out0;
wire v$S_10348_out0;
wire v$S_10442_out0;
wire v$S_10443_out0;
wire v$S_10699_out0;
wire v$S_10700_out0;
wire v$S_1226_out0;
wire v$S_12649_out0;
wire v$S_12650_out0;
wire v$S_12819_out0;
wire v$S_12820_out0;
wire v$S_15475_out0;
wire v$S_15476_out0;
wire v$S_15477_out0;
wire v$S_15478_out0;
wire v$S_16383_out0;
wire v$S_16384_out0;
wire v$S_16930_out0;
wire v$S_16931_out0;
wire v$S_16932_out0;
wire v$S_16933_out0;
wire v$S_16934_out0;
wire v$S_16935_out0;
wire v$S_16936_out0;
wire v$S_16937_out0;
wire v$S_16938_out0;
wire v$S_16939_out0;
wire v$S_16940_out0;
wire v$S_16941_out0;
wire v$S_16942_out0;
wire v$S_16943_out0;
wire v$S_16944_out0;
wire v$S_16945_out0;
wire v$S_16946_out0;
wire v$S_16947_out0;
wire v$S_16948_out0;
wire v$S_16949_out0;
wire v$S_16950_out0;
wire v$S_16951_out0;
wire v$S_17947_out0;
wire v$S_17948_out0;
wire v$S_2443_out0;
wire v$S_2444_out0;
wire v$S_4025_out0;
wire v$S_4026_out0;
wire v$S_4239_out0;
wire v$S_4240_out0;
wire v$S_5733_out0;
wire v$S_5734_out0;
wire v$S_8017_out0;
wire v$S_8018_out0;
wire v$S_8019_out0;
wire v$S_8020_out0;
wire v$S_8021_out0;
wire v$S_8167_out0;
wire v$S_8168_out0;
wire v$S_901_out0;
wire v$S_902_out0;
wire v$S_9424_out0;
wire v$S_9425_out0;
wire v$SetError_17573_out0;
wire v$SetError_17574_out0;
wire v$ShiftEN_5827_out0;
wire v$ShiftEN_5828_out0;
wire v$ShiftEN_7722_out0;
wire v$ShiftEN_7723_out0;
wire v$ShiftOut_16343_out0;
wire v$ShiftOut_16344_out0;
wire v$Shift_9605_out0;
wire v$Shift_9606_out0;
wire v$StatRegAdd1_14555_out0;
wire v$StatRegAdd1_14556_out0;
wire v$StatRegAdd_7741_out0;
wire v$StatRegAdd_7742_out0;
wire v$TAKEJUMP_10799_out0;
wire v$TAKEJUMP_10800_out0;
wire v$THRESHOLD$WRITE_7236_out0;
wire v$THRESHOLD$WRITE_7237_out0;
wire v$TWOS$COMPLEMENT$ADDER$COUT_3431_out0;
wire v$TWOS$COMPLEMENT$ADDER$COUT_3432_out0;
wire v$TXFLAG_14691_out0;
wire v$TXFLAG_14692_out0;
wire v$TXFLAG_3878_out0;
wire v$TXFLAG_3879_out0;
wire v$TXFlag_15247_out0;
wire v$TXFlag_15248_out0;
wire v$TXFlag_7718_out0;
wire v$TXFlag_7719_out0;
wire v$TXINTERRUPT_3634_out0;
wire v$TXINTERRUPT_3635_out0;
wire v$TXINT_4911_out0;
wire v$TXINT_4912_out0;
wire v$TXLast_11385_out0;
wire v$TXLast_11386_out0;
wire v$TXRST_16379_out0;
wire v$TXRST_16380_out0;
wire v$TXRST_8044_out0;
wire v$TXRST_8045_out0;
wire v$TXRegAdd_15600_out0;
wire v$TXRegAdd_15601_out0;
wire v$TXReset_17834_out0;
wire v$TXReset_17835_out0;
wire v$TXSet_12652_out0;
wire v$TXSet_12653_out0;
wire v$TXSet_14337_out0;
wire v$TXSet_14338_out0;
wire v$TXWRITE_11109_out0;
wire v$TXWRITE_11110_out0;
wire v$TXWRITE_16093_out0;
wire v$TXWRITE_16094_out0;
wire v$TXWrite_17496_out0;
wire v$TXWrite_17497_out0;
wire v$TX_11681_out0;
wire v$TX_11682_out0;
wire v$TX_1298_out0;
wire v$TX_1299_out0;
wire v$TX_18258_out0;
wire v$TX_18259_out0;
wire v$TX_420_out0;
wire v$TX_421_out0;
wire v$TXoverflow_4108_out0;
wire v$TXoverflow_4109_out0;
wire v$V0_7423_out0;
wire v$V0_9351_out0;
wire v$V1_16703_out0;
wire v$V1_17836_out0;
wire v$VALID$PREV_13429_out0;
wire v$VALID$PREV_13430_out0;
wire v$VALID0_13405_out0;
wire v$VALID1_8806_out0;
wire v$VALID_14495_out0;
wire v$VALID_14496_out0;
wire v$VALID_17917_out0;
wire v$VALID_17918_out0;
wire v$VALID_18670_out0;
wire v$VALID_18671_out0;
wire v$VALID_3712_out0;
wire v$VALID_3713_out0;
wire v$WB$HAZARD_8892_out0;
wire v$WB$HAZARD_8893_out0;
wire v$WEN$FPU_8312_out0;
wire v$WEN$FPU_8313_out0;
wire v$WEN3_1849_out0;
wire v$WEN3_1850_out0;
wire v$WEN3_3284_out0;
wire v$WEN3_3285_out0;
wire v$WENALU_16372_out0;
wire v$WENALU_16373_out0;
wire v$WENALU_18660_out0;
wire v$WENALU_18661_out0;
wire v$WENALU_4072_out0;
wire v$WENALU_4073_out0;
wire v$WENFPU_13739_out0;
wire v$WENFPU_13740_out0;
wire v$WENFPU_3498_out0;
wire v$WENFPU_3499_out0;
wire v$WENLDST_12484_out0;
wire v$WENLDST_12485_out0;
wire v$WENLDST_18629_out0;
wire v$WENLDST_18630_out0;
wire v$WENLDST_6687_out0;
wire v$WENLDST_6688_out0;
wire v$WENRAM0_9919_out0;
wire v$WENRAM1_1719_out0;
wire v$WENRAM_17082_out0;
wire v$WENRAM_17083_out0;
wire v$WENRAM_2342_out0;
wire v$WENRAM_2343_out0;
wire v$WENRAM_4969_out0;
wire v$WENRAM_4970_out0;
wire v$WEN_12173_out0;
wire v$WEN_12174_out0;
wire v$WEN_12333_out0;
wire v$WEN_12334_out0;
wire v$WEN_14218_out0;
wire v$WEN_14219_out0;
wire v$WEN_18392_out0;
wire v$WEN_18393_out0;
wire v$WEN_3683_out0;
wire v$WEN_3684_out0;
wire v$WEN_3801_out0;
wire v$WEN_3802_out0;
wire v$WR0VIEWER_15892_out0;
wire v$WR0_1316_out0;
wire v$WR0_14268_out0;
wire v$WR1VIEWER_15905_out0;
wire v$WR1_14336_out0;
wire v$WR1_303_out0;
wire v$WREN_10997_out0;
wire v$WREN_10998_out0;
wire v$WREN_2534_out0;
wire v$WREN_2535_out0;
wire v$Wordlength_5140_out0;
wire v$Wordlength_5141_out0;
wire v$Write_3255_out0;
wire v$Write_3256_out0;
wire v$Write_3257_out0;
wire v$Write_3258_out0;
wire v$Write_3259_out0;
wire v$Write_3260_out0;
wire v$Write_3261_out0;
wire v$Write_3262_out0;
wire v$Write_3263_out0;
wire v$Write_3264_out0;
wire v$Write_3265_out0;
wire v$Write_3266_out0;
wire v$Z1_16994_out0;
wire v$Z1_16995_out0;
wire v$Z1_16996_out0;
wire v$Z1_16997_out0;
wire v$Z1_16998_out0;
wire v$Z1_16999_out0;
wire v$Z1_17000_out0;
wire v$Z1_17001_out0;
wire v$Z1_17002_out0;
wire v$Z1_17003_out0;
wire v$Z1_17004_out0;
wire v$Z1_17005_out0;
wire v$Z1_17723_out0;
wire v$Z1_17724_out0;
wire v$Z1_5764_out0;
wire v$Z1_5765_out0;
wire v$Z1_5766_out0;
wire v$Z1_5767_out0;
wire v$Z1_5768_out0;
wire v$Z1_5769_out0;
wire v$Z1_5770_out0;
wire v$Z1_5771_out0;
wire v$Z2_179_out0;
wire v$Z2_180_out0;
wire v$Z2_181_out0;
wire v$Z2_182_out0;
wire v$Z2_183_out0;
wire v$Z2_184_out0;
wire v$Z2_185_out0;
wire v$Z2_186_out0;
wire v$Z2_2256_out0;
wire v$Z2_2257_out0;
wire v$Z2_6320_out0;
wire v$Z2_6321_out0;
wire v$Z2_6322_out0;
wire v$Z2_6323_out0;
wire v$Z2_6324_out0;
wire v$Z2_6325_out0;
wire v$Z2_6326_out0;
wire v$Z2_6327_out0;
wire v$Z2_6328_out0;
wire v$Z2_6329_out0;
wire v$Z2_6330_out0;
wire v$Z2_6331_out0;
wire v$Z3_11986_out0;
wire v$Z3_11987_out0;
wire v$Z3_17777_out0;
wire v$Z3_17778_out0;
wire v$Z3_17779_out0;
wire v$Z3_17780_out0;
wire v$Z3_17781_out0;
wire v$Z3_17782_out0;
wire v$Z3_17783_out0;
wire v$Z3_17784_out0;
wire v$Z3_17785_out0;
wire v$Z3_17786_out0;
wire v$Z4_7919_out0;
wire v$Z4_7920_out0;
wire v$Z4_7921_out0;
wire v$Z4_7922_out0;
wire v$Z4_7923_out0;
wire v$Z4_7924_out0;
wire v$Z4_7925_out0;
wire v$Z4_7926_out0;
wire v$Z_10329_out0;
wire v$Z_10330_out0;
wire v$Z_10331_out0;
wire v$Z_10332_out0;
wire v$Z_10333_out0;
wire v$Z_10334_out0;
wire v$Z_10335_out0;
wire v$Z_10336_out0;
wire v$Z_12553_out0;
wire v$Z_12554_out0;
wire v$Z_12555_out0;
wire v$Z_12556_out0;
wire v$Z_12557_out0;
wire v$Z_12558_out0;
wire v$Z_12559_out0;
wire v$Z_12560_out0;
wire v$Z_12561_out0;
wire v$Z_12562_out0;
wire v$Z_12563_out0;
wire v$Z_12564_out0;
wire v$Z_12565_out0;
wire v$Z_12566_out0;
wire v$Z_12567_out0;
wire v$Z_12568_out0;
wire v$Z_12569_out0;
wire v$Z_12570_out0;
wire v$Z_12571_out0;
wire v$Z_12572_out0;
wire v$Z_12573_out0;
wire v$Z_12574_out0;
wire v$Z_12575_out0;
wire v$Z_12576_out0;
wire v$Z_12577_out0;
wire v$Z_12578_out0;
wire v$Z_12579_out0;
wire v$Z_12580_out0;
wire v$Z_12581_out0;
wire v$Z_12582_out0;
wire v$Z_12583_out0;
wire v$Z_12584_out0;
wire v$Z_12585_out0;
wire v$Z_12586_out0;
wire v$Z_12587_out0;
wire v$Z_12588_out0;
wire v$Z_12589_out0;
wire v$Z_12590_out0;
wire v$Z_12591_out0;
wire v$Z_12592_out0;
wire v$Z_12593_out0;
wire v$Z_12594_out0;
wire v$Z_12595_out0;
wire v$Z_12596_out0;
wire v$Z_12597_out0;
wire v$Z_12598_out0;
wire v$Z_12599_out0;
wire v$Z_12600_out0;
wire v$Z_13551_out0;
wire v$Z_13552_out0;
wire v$Z_15808_out0;
wire v$Z_15809_out0;
wire v$Z_15810_out0;
wire v$Z_15811_out0;
wire v$Z_2551_out0;
wire v$Z_2552_out0;
wire v$Z_2553_out0;
wire v$Z_2554_out0;
wire v$Z_2555_out0;
wire v$Z_2556_out0;
wire v$Z_2557_out0;
wire v$Z_2558_out0;
wire v$Z_2559_out0;
wire v$Z_2560_out0;
wire v$Z_2561_out0;
wire v$Z_2562_out0;
wire v$_10244_out0;
wire v$_10244_out1;
wire v$_10245_out0;
wire v$_10245_out1;
wire v$_10278_out0;
wire v$_10279_out0;
wire v$_10284_out0;
wire v$_10284_out1;
wire v$_10285_out0;
wire v$_10285_out1;
wire v$_10286_out0;
wire v$_10286_out1;
wire v$_10287_out0;
wire v$_10287_out1;
wire v$_10288_out0;
wire v$_10288_out1;
wire v$_10416_out0;
wire v$_10417_out0;
wire v$_10446_out0;
wire v$_10447_out0;
wire v$_10448_out0;
wire v$_10449_out0;
wire v$_10450_out0;
wire v$_10772_out0;
wire v$_10773_out0;
wire v$_10774_out0;
wire v$_10775_out0;
wire v$_10776_out0;
wire v$_10787_out0;
wire v$_10788_out0;
wire v$_10910_out0;
wire v$_10911_out0;
wire v$_10912_out0;
wire v$_10913_out0;
wire v$_10914_out0;
wire v$_11022_out0;
wire v$_11022_out1;
wire v$_11023_out0;
wire v$_11023_out1;
wire v$_11024_out0;
wire v$_11024_out1;
wire v$_11025_out0;
wire v$_11025_out1;
wire v$_11026_out0;
wire v$_11026_out1;
wire v$_11056_out0;
wire v$_11056_out1;
wire v$_11057_out0;
wire v$_11057_out1;
wire v$_11099_out0;
wire v$_11100_out0;
wire v$_11101_out0;
wire v$_11102_out0;
wire v$_11103_out0;
wire v$_11391_out0;
wire v$_11392_out0;
wire v$_11618_out0;
wire v$_11618_out1;
wire v$_11619_out0;
wire v$_11619_out1;
wire v$_11620_out0;
wire v$_11620_out1;
wire v$_11621_out0;
wire v$_11621_out1;
wire v$_11622_out0;
wire v$_11622_out1;
wire v$_11765_out0;
wire v$_11766_out0;
wire v$_11858_out0;
wire v$_11858_out1;
wire v$_11859_out0;
wire v$_11859_out1;
wire v$_11860_out0;
wire v$_11860_out1;
wire v$_11861_out0;
wire v$_11861_out1;
wire v$_11862_out0;
wire v$_11862_out1;
wire v$_11863_out0;
wire v$_11863_out1;
wire v$_11864_out0;
wire v$_11864_out1;
wire v$_11865_out0;
wire v$_11865_out1;
wire v$_11866_out0;
wire v$_11866_out1;
wire v$_11867_out0;
wire v$_11867_out1;
wire v$_11868_out0;
wire v$_11868_out1;
wire v$_11869_out0;
wire v$_11869_out1;
wire v$_1197_out0;
wire v$_1198_out0;
wire v$_12077_out0;
wire v$_12077_out1;
wire v$_12078_out0;
wire v$_12078_out1;
wire v$_12080_out0;
wire v$_12080_out1;
wire v$_12081_out0;
wire v$_12081_out1;
wire v$_12764_out0;
wire v$_12765_out0;
wire v$_12772_out0;
wire v$_12773_out0;
wire v$_1302_out0;
wire v$_1303_out0;
wire v$_1304_out0;
wire v$_1305_out0;
wire v$_1306_out0;
wire v$_13180_out0;
wire v$_13180_out1;
wire v$_13181_out0;
wire v$_13181_out1;
wire v$_13182_out0;
wire v$_13182_out1;
wire v$_13183_out0;
wire v$_13183_out1;
wire v$_13184_out0;
wire v$_13184_out1;
wire v$_13269_out0;
wire v$_13272_out0;
wire v$_13289_out0;
wire v$_13290_out0;
wire v$_1353_out0;
wire v$_13542_out0;
wire v$_13543_out0;
wire v$_1354_out0;
wire v$_1355_out0;
wire v$_1356_out0;
wire v$_1357_out0;
wire v$_13691_out0;
wire v$_13692_out0;
wire v$_13842_out0;
wire v$_13842_out1;
wire v$_13843_out0;
wire v$_13843_out1;
wire v$_14078_out0;
wire v$_14078_out1;
wire v$_14079_out0;
wire v$_14079_out1;
wire v$_14247_out0;
wire v$_14247_out1;
wire v$_14248_out0;
wire v$_14248_out1;
wire v$_14324_out0;
wire v$_14325_out0;
wire v$_14509_out0;
wire v$_14509_out1;
wire v$_14510_out0;
wire v$_14510_out1;
wire v$_14511_out0;
wire v$_14511_out1;
wire v$_14512_out0;
wire v$_14512_out1;
wire v$_14513_out0;
wire v$_14513_out1;
wire v$_14514_out0;
wire v$_14514_out1;
wire v$_14515_out0;
wire v$_14515_out1;
wire v$_14516_out0;
wire v$_14516_out1;
wire v$_14517_out0;
wire v$_14517_out1;
wire v$_14518_out0;
wire v$_14518_out1;
wire v$_14519_out0;
wire v$_14519_out1;
wire v$_14520_out0;
wire v$_14520_out1;
wire v$_14521_out0;
wire v$_14521_out1;
wire v$_14522_out0;
wire v$_14522_out1;
wire v$_14645_out0;
wire v$_14645_out1;
wire v$_14646_out0;
wire v$_14646_out1;
wire v$_15138_out0;
wire v$_15139_out0;
wire v$_15148_out0;
wire v$_15149_out0;
wire v$_15150_out0;
wire v$_15151_out0;
wire v$_15152_out0;
wire v$_15186_out0;
wire v$_15186_out1;
wire v$_15187_out0;
wire v$_15187_out1;
wire v$_15188_out0;
wire v$_15188_out1;
wire v$_15189_out0;
wire v$_15189_out1;
wire v$_15320_out0;
wire v$_15320_out1;
wire v$_15321_out0;
wire v$_15321_out1;
wire v$_1553_out0;
wire v$_1554_out0;
wire v$_15741_out0;
wire v$_15741_out1;
wire v$_15742_out0;
wire v$_15742_out1;
wire v$_15743_out0;
wire v$_15743_out1;
wire v$_15744_out0;
wire v$_15744_out1;
wire v$_15745_out0;
wire v$_15745_out1;
wire v$_15839_out0;
wire v$_15839_out1;
wire v$_15840_out0;
wire v$_15840_out1;
wire v$_16130_out0;
wire v$_16131_out0;
wire v$_16132_out0;
wire v$_16133_out0;
wire v$_16134_out0;
wire v$_16137_out0;
wire v$_16137_out1;
wire v$_16138_out0;
wire v$_16138_out1;
wire v$_16182_out0;
wire v$_16182_out1;
wire v$_16183_out0;
wire v$_16183_out1;
wire v$_16184_out0;
wire v$_16184_out1;
wire v$_16185_out0;
wire v$_16185_out1;
wire v$_16186_out0;
wire v$_16186_out1;
wire v$_16265_out0;
wire v$_16266_out0;
wire v$_16267_out0;
wire v$_16268_out0;
wire v$_16269_out0;
wire v$_1639_out0;
wire v$_1639_out1;
wire v$_1640_out0;
wire v$_1640_out1;
wire v$_1641_out0;
wire v$_1641_out1;
wire v$_1642_out0;
wire v$_1642_out1;
wire v$_1643_out0;
wire v$_1643_out1;
wire v$_1644_out0;
wire v$_1644_out1;
wire v$_1645_out0;
wire v$_1645_out1;
wire v$_1646_out0;
wire v$_1646_out1;
wire v$_1647_out0;
wire v$_1647_out1;
wire v$_1648_out0;
wire v$_1648_out1;
wire v$_1649_out0;
wire v$_1649_out1;
wire v$_1650_out0;
wire v$_1650_out1;
wire v$_16550_out0;
wire v$_16550_out1;
wire v$_16551_out0;
wire v$_16551_out1;
wire v$_16589_out0;
wire v$_16589_out1;
wire v$_16590_out0;
wire v$_16590_out1;
wire v$_16591_out0;
wire v$_16591_out1;
wire v$_16592_out0;
wire v$_16592_out1;
wire v$_16593_out0;
wire v$_16593_out1;
wire v$_16704_out0;
wire v$_16704_out1;
wire v$_16705_out0;
wire v$_16705_out1;
wire v$_16706_out0;
wire v$_16706_out1;
wire v$_16707_out0;
wire v$_16707_out1;
wire v$_16708_out0;
wire v$_16708_out1;
wire v$_16740_out0;
wire v$_16741_out0;
wire v$_16742_out0;
wire v$_16743_out0;
wire v$_16744_out0;
wire v$_16980_out0;
wire v$_16980_out1;
wire v$_16981_out0;
wire v$_16981_out1;
wire v$_17325_out0;
wire v$_17325_out1;
wire v$_17326_out0;
wire v$_17326_out1;
wire v$_17327_out0;
wire v$_17327_out1;
wire v$_17328_out0;
wire v$_17328_out1;
wire v$_17329_out0;
wire v$_17329_out1;
wire v$_17755_out0;
wire v$_17755_out1;
wire v$_17756_out0;
wire v$_17756_out1;
wire v$_17757_out0;
wire v$_17757_out1;
wire v$_17758_out0;
wire v$_17758_out1;
wire v$_17759_out0;
wire v$_17759_out1;
wire v$_17981_out0;
wire v$_17981_out1;
wire v$_17982_out0;
wire v$_17982_out1;
wire v$_18018_out0;
wire v$_18019_out0;
wire v$_18188_out0;
wire v$_18189_out0;
wire v$_18190_out0;
wire v$_18191_out0;
wire v$_18192_out0;
wire v$_18297_out0;
wire v$_18298_out0;
wire v$_1854_out0;
wire v$_1855_out0;
wire v$_1856_out0;
wire v$_1857_out0;
wire v$_1858_out0;
wire v$_1966_out0;
wire v$_1967_out0;
wire v$_2447_out0;
wire v$_2448_out0;
wire v$_2652_out0;
wire v$_2653_out0;
wire v$_2922_out0;
wire v$_2923_out0;
wire v$_2924_out0;
wire v$_2925_out0;
wire v$_2926_out0;
wire v$_2982_out0;
wire v$_2983_out0;
wire v$_3109_out0;
wire v$_3109_out1;
wire v$_3110_out0;
wire v$_3110_out1;
wire v$_3118_out0;
wire v$_3118_out1;
wire v$_3119_out0;
wire v$_3119_out1;
wire v$_330_out0;
wire v$_330_out1;
wire v$_331_out0;
wire v$_331_out1;
wire v$_3486_out0;
wire v$_3486_out1;
wire v$_3487_out0;
wire v$_3487_out1;
wire v$_3685_out0;
wire v$_3685_out1;
wire v$_3686_out0;
wire v$_3686_out1;
wire v$_3787_out0;
wire v$_3787_out1;
wire v$_3788_out0;
wire v$_3788_out1;
wire v$_3992_out0;
wire v$_3992_out1;
wire v$_3993_out0;
wire v$_3993_out1;
wire v$_4015_out0;
wire v$_4015_out1;
wire v$_4016_out0;
wire v$_4016_out1;
wire v$_4019_out0;
wire v$_4019_out1;
wire v$_4020_out0;
wire v$_4020_out1;
wire v$_41_out0;
wire v$_42_out0;
wire v$_4774_out0;
wire v$_4774_out1;
wire v$_4775_out0;
wire v$_4775_out1;
wire v$_4892_out0;
wire v$_4892_out1;
wire v$_4893_out0;
wire v$_4893_out1;
wire v$_4896_out1;
wire v$_4897_out1;
wire v$_5040_out0;
wire v$_5040_out1;
wire v$_5041_out0;
wire v$_5041_out1;
wire v$_5074_out0;
wire v$_5074_out1;
wire v$_5075_out0;
wire v$_5075_out1;
wire v$_5405_out0;
wire v$_5405_out1;
wire v$_5406_out0;
wire v$_5406_out1;
wire v$_5786_out0;
wire v$_5786_out1;
wire v$_5787_out0;
wire v$_5787_out1;
wire v$_5948_out0;
wire v$_5948_out1;
wire v$_5949_out0;
wire v$_5949_out1;
wire v$_5950_out0;
wire v$_5950_out1;
wire v$_5951_out0;
wire v$_5951_out1;
wire v$_5952_out0;
wire v$_5952_out1;
wire v$_6075_out0;
wire v$_6076_out0;
wire v$_6898_out0;
wire v$_6898_out1;
wire v$_6899_out0;
wire v$_6899_out1;
wire v$_6900_out0;
wire v$_6900_out1;
wire v$_6901_out0;
wire v$_6901_out1;
wire v$_6902_out0;
wire v$_6902_out1;
wire v$_6977_out0;
wire v$_6977_out1;
wire v$_6978_out0;
wire v$_6978_out1;
wire v$_6979_out0;
wire v$_6979_out1;
wire v$_6980_out0;
wire v$_6980_out1;
wire v$_6981_out0;
wire v$_6981_out1;
wire v$_6982_out0;
wire v$_6982_out1;
wire v$_6983_out0;
wire v$_6983_out1;
wire v$_7067_out0;
wire v$_7068_out0;
wire v$_7069_out0;
wire v$_7070_out0;
wire v$_7071_out0;
wire v$_7245_out0;
wire v$_7245_out1;
wire v$_7246_out0;
wire v$_7246_out1;
wire v$_7287_out0;
wire v$_7287_out1;
wire v$_7288_out0;
wire v$_7288_out1;
wire v$_7289_out0;
wire v$_7290_out0;
wire v$_7358_out0;
wire v$_7358_out1;
wire v$_7359_out0;
wire v$_7359_out1;
wire v$_7360_out0;
wire v$_7360_out1;
wire v$_7361_out0;
wire v$_7361_out1;
wire v$_7362_out0;
wire v$_7362_out1;
wire v$_7395_out0;
wire v$_7395_out1;
wire v$_7396_out0;
wire v$_7396_out1;
wire v$_7476_out0;
wire v$_7477_out0;
wire v$_7656_out0;
wire v$_7656_out1;
wire v$_7657_out0;
wire v$_7657_out1;
wire v$_7658_out0;
wire v$_7658_out1;
wire v$_7659_out0;
wire v$_7659_out1;
wire v$_7660_out0;
wire v$_7660_out1;
wire v$_7661_out0;
wire v$_7661_out1;
wire v$_7662_out0;
wire v$_7662_out1;
wire v$_7663_out0;
wire v$_7663_out1;
wire v$_7664_out0;
wire v$_7664_out1;
wire v$_7665_out0;
wire v$_7665_out1;
wire v$_7666_out0;
wire v$_7666_out1;
wire v$_7667_out0;
wire v$_7667_out1;
wire v$_7768_out0;
wire v$_7769_out0;
wire v$_7770_out0;
wire v$_7771_out0;
wire v$_7772_out0;
wire v$_7981_out0;
wire v$_7981_out1;
wire v$_7982_out0;
wire v$_7982_out1;
wire v$_8090_out0;
wire v$_8090_out1;
wire v$_8091_out0;
wire v$_8091_out1;
wire v$_8232_out0;
wire v$_8233_out0;
wire v$_8774_out0;
wire v$_8775_out0;
wire v$_8776_out0;
wire v$_8776_out1;
wire v$_8777_out0;
wire v$_8777_out1;
wire v$_8812_out0;
wire v$_8812_out1;
wire v$_8813_out0;
wire v$_8813_out1;
wire v$_893_out0;
wire v$_894_out0;
wire v$_9062_out0;
wire v$_9063_out0;
wire v$_9064_out0;
wire v$_9065_out0;
wire v$_9066_out0;
wire v$_9070_out0;
wire v$_9070_out1;
wire v$_9071_out0;
wire v$_9071_out1;
wire v$_9110_out0;
wire v$_9110_out1;
wire v$_9111_out0;
wire v$_9111_out1;
wire v$_9372_out0;
wire v$_9372_out1;
wire v$_9373_out0;
wire v$_9373_out1;
wire v$_9381_out0;
wire v$_9381_out1;
wire v$_9382_out0;
wire v$_9382_out1;
wire v$_9383_out0;
wire v$_9383_out1;
wire v$_9384_out0;
wire v$_9384_out1;
wire v$_9385_out0;
wire v$_9385_out1;
wire v$_9482_out0;
wire v$_9482_out1;
wire v$_9483_out0;
wire v$_9483_out1;
wire v$_9497_out0;
wire v$_9497_out1;
wire v$_9498_out0;
wire v$_9498_out1;
wire v$_9499_out0;
wire v$_9499_out1;
wire v$_9500_out0;
wire v$_9500_out1;
wire v$_9501_out0;
wire v$_9501_out1;
wire v$_9580_out0;
wire v$_9581_out0;
wire v$increment_17844_out0;
wire v$increment_17845_out0;

always @(posedge clk) v$FF1_2_out0 <= v$NEWINTERRUPT_7025_out0;
always @(posedge clk) v$FF1_3_out0 <= v$NEWINTERRUPT_7026_out0;
always @(posedge clk) v$FF1_191_out0 <= v$G3_8040_out0;
always @(posedge clk) v$FF1_192_out0 <= v$G3_8041_out0;
always @(posedge clk) v$INT2_256_out0 <= v$I2EN_15746_out0 ? v$SEL1_11971_out0 : v$INT2_256_out0;
always @(posedge clk) v$INT2_257_out0 <= v$I2EN_15747_out0 ? v$SEL1_11972_out0 : v$INT2_257_out0;
always @(posedge clk) v$FF3_262_out0 <= v$ShiftEN_7722_out0 ? v$MUX3_17725_out0 : v$FF3_262_out0;
always @(posedge clk) v$FF3_263_out0 <= v$ShiftEN_7723_out0 ? v$MUX3_17726_out0 : v$FF3_263_out0;
always @(posedge clk) v$INT3_271_out0 <= v$I3EN_17775_out0 ? v$SEL1_11971_out0 : v$INT3_271_out0;
always @(posedge clk) v$INT3_272_out0 <= v$I3EN_17776_out0 ? v$SEL1_11972_out0 : v$INT3_272_out0;
always @(posedge clk) v$REG13_296_out0 <= v$HALT0_361_out0;
always @(posedge clk) v$FF0_655_out0 <= v$CLK4_12213_out0 ? v$G1_15293_out0 : v$FF0_655_out0;
always @(posedge clk) v$FF0_656_out0 <= v$CLK4_12214_out0 ? v$G1_15294_out0 : v$FF0_656_out0;
always @(posedge clk) v$REG2_657_out0 <= v$increment_17844_out0 ? v$A2_14825_out0 : v$REG2_657_out0;
always @(posedge clk) v$REG2_658_out0 <= v$increment_17845_out0 ? v$A2_14826_out0 : v$REG2_658_out0;
always @(posedge clk) v$REG1_1163_out0 <= v$G14_15815_out0 ? v$A_11042_out0 : v$REG1_1163_out0;
always @(posedge clk) v$REG1_1164_out0 <= v$G14_15816_out0 ? v$A_11043_out0 : v$REG1_1164_out0;
always @(posedge clk) v$FF1_1178_out0 <= v$CLK4_12213_out0 ? v$G21_17674_out0 : v$FF1_1178_out0;
always @(posedge clk) v$FF1_1179_out0 <= v$CLK4_12214_out0 ? v$G21_17675_out0 : v$FF1_1179_out0;
always @(posedge clk) v$FF2_1180_out0 <= v$LDMAIN_13807_out0;
always @(posedge clk) v$FF2_1181_out0 <= v$LDMAIN_13808_out0;
always @(posedge clk) v$FF3_1296_out0 <= v$Shift_9605_out0 ? v$FF1_16187_out0 : v$FF3_1296_out0;
always @(posedge clk) v$FF3_1297_out0 <= v$Shift_9606_out0 ? v$FF1_16188_out0 : v$FF3_1297_out0;
always @(posedge clk) v$FF1_1376_out0 <= v$NEWINTERRUPT_4431_out0;
always @(posedge clk) v$FF1_1377_out0 <= v$NEWINTERRUPT_4432_out0;
always @(posedge clk) v$FF2_1572_out0 <= v$Shift_9605_out0 ? v$FF7_14553_out0 : v$FF2_1572_out0;
always @(posedge clk) v$FF2_1573_out0 <= v$Shift_9606_out0 ? v$FF7_14554_out0 : v$FF2_1573_out0;
always @(posedge clk) v$FF5_1754_out0 <= v$SHIFTEN_9406_out0 ? v$MUX1_2582_out0 : v$FF5_1754_out0;
always @(posedge clk) v$FF5_1755_out0 <= v$SHIFTEN_9407_out0 ? v$MUX1_2583_out0 : v$FF5_1755_out0;
always @(posedge clk) v$FF5_1756_out0 <= v$SHIFTEN_9408_out0 ? v$MUX1_2584_out0 : v$FF5_1756_out0;
always @(posedge clk) v$FF5_1757_out0 <= v$SHIFTEN_9409_out0 ? v$MUX1_2585_out0 : v$FF5_1757_out0;
always @(posedge clk) v$FF5_1758_out0 <= v$SHIFTEN_9410_out0 ? v$MUX1_2586_out0 : v$FF5_1758_out0;
always @(posedge clk) v$FF5_1759_out0 <= v$SHIFTEN_9411_out0 ? v$MUX1_2587_out0 : v$FF5_1759_out0;
always @(posedge clk) v$FF5_1760_out0 <= v$SHIFTEN_9412_out0 ? v$MUX1_2588_out0 : v$FF5_1760_out0;
always @(posedge clk) v$FF5_1761_out0 <= v$SHIFTEN_9413_out0 ? v$MUX1_2589_out0 : v$FF5_1761_out0;
always @(posedge clk) v$FF5_1762_out0 <= v$SHIFTEN_9414_out0 ? v$MUX1_2590_out0 : v$FF5_1762_out0;
always @(posedge clk) v$FF5_1763_out0 <= v$SHIFTEN_9415_out0 ? v$MUX1_2591_out0 : v$FF5_1763_out0;
always @(posedge clk) v$FF5_1764_out0 <= v$SHIFTEN_9416_out0 ? v$MUX1_2592_out0 : v$FF5_1764_out0;
always @(posedge clk) v$FF5_1765_out0 <= v$SHIFTEN_9417_out0 ? v$MUX1_2593_out0 : v$FF5_1765_out0;
always @(posedge clk) v$FF4_2347_out0 <= v$ShiftEN_7722_out0 ? v$MUX4_15635_out0 : v$FF4_2347_out0;
always @(posedge clk) v$FF4_2348_out0 <= v$ShiftEN_7723_out0 ? v$MUX4_15636_out0 : v$FF4_2348_out0;
always @(posedge clk) v$FF11_2449_out0 <= v$G50_16361_out0;
always @(posedge clk) v$FF11_2450_out0 <= v$G50_16362_out0;
always @(posedge clk) v$FF1_2525_out0 <= v$G4_14683_out0;
always @(posedge clk) v$FF1_2526_out0 <= v$G4_14684_out0;
always @(posedge clk) v$FF6_2621_out0 <= v$SHIFTEN_9406_out0 ? v$MUX3_9950_out0 : v$FF6_2621_out0;
always @(posedge clk) v$FF6_2622_out0 <= v$SHIFTEN_9407_out0 ? v$MUX3_9951_out0 : v$FF6_2622_out0;
always @(posedge clk) v$FF6_2623_out0 <= v$SHIFTEN_9408_out0 ? v$MUX3_9952_out0 : v$FF6_2623_out0;
always @(posedge clk) v$FF6_2624_out0 <= v$SHIFTEN_9409_out0 ? v$MUX3_9953_out0 : v$FF6_2624_out0;
always @(posedge clk) v$FF6_2625_out0 <= v$SHIFTEN_9410_out0 ? v$MUX3_9954_out0 : v$FF6_2625_out0;
always @(posedge clk) v$FF6_2626_out0 <= v$SHIFTEN_9411_out0 ? v$MUX3_9955_out0 : v$FF6_2626_out0;
always @(posedge clk) v$FF6_2627_out0 <= v$SHIFTEN_9412_out0 ? v$MUX3_9956_out0 : v$FF6_2627_out0;
always @(posedge clk) v$FF6_2628_out0 <= v$SHIFTEN_9413_out0 ? v$MUX3_9957_out0 : v$FF6_2628_out0;
always @(posedge clk) v$FF6_2629_out0 <= v$SHIFTEN_9414_out0 ? v$MUX3_9958_out0 : v$FF6_2629_out0;
always @(posedge clk) v$FF6_2630_out0 <= v$SHIFTEN_9415_out0 ? v$MUX3_9959_out0 : v$FF6_2630_out0;
always @(posedge clk) v$FF6_2631_out0 <= v$SHIFTEN_9416_out0 ? v$MUX3_9960_out0 : v$FF6_2631_out0;
always @(posedge clk) v$FF6_2632_out0 <= v$SHIFTEN_9417_out0 ? v$MUX3_9961_out0 : v$FF6_2632_out0;
always @(posedge clk) v$REG3_2822_out0 <= v$G55_18199_out0 ? v$MUX5_11943_out0 : v$REG3_2822_out0;
always @(posedge clk) v$REG3_2823_out0 <= v$G55_18200_out0 ? v$MUX5_11944_out0 : v$REG3_2823_out0;
always @(posedge clk) v$FF2_2951_out0 <= v$ShiftEN_7722_out0 ? v$MUX2_13287_out0 : v$FF2_2951_out0;
always @(posedge clk) v$FF2_2952_out0 <= v$ShiftEN_7723_out0 ? v$MUX2_13288_out0 : v$FF2_2952_out0;
always @(posedge clk) v$REG12_3330_out0 <= v$HALT1_4159_out0 ? v$RAMADDR1_12657_out0 : v$REG12_3330_out0;
always @(posedge clk) v$FF3_3378_out0 <= v$G53_17493_out0;
always @(posedge clk) v$FF4_3781_out0 <= v$CAPTURE_242_out0 ? v$G6_12126_out0 : v$FF4_3781_out0;
always @(posedge clk) v$FF4_3782_out0 <= v$CAPTURE_243_out0 ? v$G6_12127_out0 : v$FF4_3782_out0;
always @(posedge clk) v$REG1_4043_out0 <= v$EN_15897_out0 ? v$MODE_10801_out0 : v$REG1_4043_out0;
always @(posedge clk) v$REG1_4044_out0 <= v$EN_15898_out0 ? v$MODE_10802_out0 : v$REG1_4044_out0;
always @(posedge clk) v$REG2_4047_out0 <= v$START_5492_out0 ? v$_1852_out0 : v$REG2_4047_out0;
always @(posedge clk) v$REG8_4106_out0 <= v$SELIN_18215_out0;
always @(posedge clk) v$FF0_4326_out0 <= v$CLK4_17983_out0 ? v$MUX1_7642_out0 : v$FF0_4326_out0;
always @(posedge clk) v$FF0_4327_out0 <= v$CLK4_17984_out0 ? v$MUX1_7643_out0 : v$FF0_4327_out0;
always @(posedge clk) v$FF1_4339_out0 <= v$START_5492_out0 ? v$IS$32$BITS_14038_out0 : v$FF1_4339_out0;
always @(posedge clk) v$FF2_4345_out0 <= v$CLK4_17983_out0 ? v$MUX3_6131_out0 : v$FF2_4345_out0;
always @(posedge clk) v$FF2_4346_out0 <= v$CLK4_17984_out0 ? v$MUX3_6132_out0 : v$FF2_4346_out0;
always @(posedge clk) v$FF5_4744_out0 <= v$EQ2_11605_out0;
always @(posedge clk) v$FF5_4745_out0 <= v$EQ2_11606_out0;
always @(posedge clk) v$REG1_4894_out0 <= v$D1_14097_out1 ? v$DIN3_14418_out0 : v$REG1_4894_out0;
always @(posedge clk) v$REG1_4895_out0 <= v$D1_14098_out1 ? v$DIN3_14419_out0 : v$REG1_4895_out0;
always @(posedge clk) v$FF0_5007_out0 <= v$G1_13147_out0;
always @(posedge clk) v$FF0_5008_out0 <= v$G1_13148_out0;
always @(posedge clk) v$REG2_5128_out0 <= v$HALT_16371_out0 ? v$G8_15731_out0 : v$REG2_5128_out0;
always @(posedge clk) v$FF1_5226_out0 <= v$NEXTSTATE_13535_out0;
always @(posedge clk) v$FF1_5227_out0 <= v$NEXTSTATE_13536_out0;
always @(posedge clk) v$FF1_5228_out0 <= v$NEXTSTATE_13537_out0;
always @(posedge clk) v$FF1_5229_out0 <= v$NEXTSTATE_13538_out0;
always @(posedge clk) v$FF1_5448_out0 <= v$G45_15360_out0;
always @(posedge clk) v$REG14_5459_out0 <= v$HALT1_4159_out0;
always @(posedge clk) v$FF1_6026_out0 <= v$INTERRUPT0_11700_out0;
always @(posedge clk) v$FF1_6027_out0 <= v$INTERRUPT0_11701_out0;
always @(posedge clk) v$FF1_6149_out0 <= v$CAPTURE_242_out0 ? v$I3_4823_out0 : v$FF1_6149_out0;
always @(posedge clk) v$FF1_6150_out0 <= v$CAPTURE_243_out0 ? v$I3_4824_out0 : v$FF1_6150_out0;
always @(posedge clk) v$REG7_6181_out0 <= v$G84_1235_out0;
always @(posedge clk) v$REG4_6650_out0 <= v$G66_8673_out0 ? v$MUX1_15262_out0 : v$REG4_6650_out0;
always @(posedge clk) v$REG4_6651_out0 <= v$G66_8674_out0 ? v$MUX1_15263_out0 : v$REG4_6651_out0;
always @(posedge clk) v$REG3_6998_out0 <= v$EXEC1_18513_out0 ? v$_1606_out0 : v$REG3_6998_out0;
always @(posedge clk) v$FF4_7017_out0 <= v$EQ1_14322_out0;
always @(posedge clk) v$FF4_7018_out0 <= v$EQ1_14323_out0;
always @(posedge clk) v$REG1_7074_out0 <= v$HALTVALID_7744_out0 ? v$NEXTSTATE_13539_out0 : v$REG1_7074_out0;
always @(posedge clk) v$FF3_7331_out0 <= v$RX_43_out0;
always @(posedge clk) v$FF3_7332_out0 <= v$RX_44_out0;
always @(posedge clk) v$FF3_7563_out0 <= v$CAPTURE_242_out0 ? v$G9_15531_out0 : v$FF3_7563_out0;
always @(posedge clk) v$FF3_7564_out0 <= v$CAPTURE_243_out0 ? v$G9_15532_out0 : v$FF3_7564_out0;
always @(posedge clk) v$REG1_7848_out0 <= v$START_5492_out0 ? v$_12523_out0 : v$REG1_7848_out0;
always @(posedge clk) v$FF10_7890_out0 <= v$HALT_12900_out0;
always @(posedge clk) v$FF10_7891_out0 <= v$HALT_12901_out0;
always @(posedge clk) v$FF8_8026_out0 <= v$ShiftEN_7722_out0 ? v$MUX8_1496_out0 : v$FF8_8026_out0;
always @(posedge clk) v$FF8_8027_out0 <= v$ShiftEN_7723_out0 ? v$MUX8_1497_out0 : v$FF8_8027_out0;
always @(posedge clk) v$FF4_8055_out0 <= v$G68_15184_out0;
always @(posedge clk) v$FF4_8056_out0 <= v$G68_15185_out0;
always @(posedge clk) v$FF7_8087_out0 <= v$G62_11755_out0 ? v$R_8778_out0 : v$FF7_8087_out0;
always @(posedge clk) v$FF7_8088_out0 <= v$G62_11756_out0 ? v$R_8779_out0 : v$FF7_8088_out0;
always @(posedge clk) v$FF1_8223_out0 <= v$EXEC2_8048_out0 ? v$S_17947_out0 : v$FF1_8223_out0;
always @(posedge clk) v$FF1_8224_out0 <= v$EXEC2_8049_out0 ? v$S_17948_out0 : v$FF1_8224_out0;
always @(posedge clk) v$FF4_8252_out0 <= v$Shift_9605_out0 ? v$RX_2966_out0 : v$FF4_8252_out0;
always @(posedge clk) v$FF4_8253_out0 <= v$Shift_9606_out0 ? v$RX_2967_out0 : v$FF4_8253_out0;
always @(posedge clk) v$FF7_8298_out0 <= v$SHIFTEN_9406_out0 ? v$MUX8_3603_out0 : v$FF7_8298_out0;
always @(posedge clk) v$FF7_8299_out0 <= v$SHIFTEN_9407_out0 ? v$MUX8_3604_out0 : v$FF7_8299_out0;
always @(posedge clk) v$FF7_8300_out0 <= v$SHIFTEN_9408_out0 ? v$MUX8_3605_out0 : v$FF7_8300_out0;
always @(posedge clk) v$FF7_8301_out0 <= v$SHIFTEN_9409_out0 ? v$MUX8_3606_out0 : v$FF7_8301_out0;
always @(posedge clk) v$FF7_8302_out0 <= v$SHIFTEN_9410_out0 ? v$MUX8_3607_out0 : v$FF7_8302_out0;
always @(posedge clk) v$FF7_8303_out0 <= v$SHIFTEN_9411_out0 ? v$MUX8_3608_out0 : v$FF7_8303_out0;
always @(posedge clk) v$FF7_8304_out0 <= v$SHIFTEN_9412_out0 ? v$MUX8_3609_out0 : v$FF7_8304_out0;
always @(posedge clk) v$FF7_8305_out0 <= v$SHIFTEN_9413_out0 ? v$MUX8_3610_out0 : v$FF7_8305_out0;
always @(posedge clk) v$FF7_8306_out0 <= v$SHIFTEN_9414_out0 ? v$MUX8_3611_out0 : v$FF7_8306_out0;
always @(posedge clk) v$FF7_8307_out0 <= v$SHIFTEN_9415_out0 ? v$MUX8_3612_out0 : v$FF7_8307_out0;
always @(posedge clk) v$FF7_8308_out0 <= v$SHIFTEN_9416_out0 ? v$MUX8_3613_out0 : v$FF7_8308_out0;
always @(posedge clk) v$FF7_8309_out0 <= v$SHIFTEN_9417_out0 ? v$MUX8_3614_out0 : v$FF7_8309_out0;
always @(posedge clk) v$REG1_8824_out0 <= v$G6_3503_out0;
always @(posedge clk) v$REG1_8890_out0 <= v$EXEC2_9439_out0 ? v$MUX5_14489_out0 : v$REG1_8890_out0;
always @(posedge clk) v$REG1_8891_out0 <= v$EXEC2_9440_out0 ? v$MUX5_14490_out0 : v$REG1_8891_out0;
always @(posedge clk) v$FF6_8963_out0 <= v$Shift_9605_out0 ? v$FF8_16727_out0 : v$FF6_8963_out0;
always @(posedge clk) v$FF6_8964_out0 <= v$Shift_9606_out0 ? v$FF8_16728_out0 : v$FF6_8964_out0;
always @(posedge clk) v$FF0_9401_out0 <= v$G12_2215_out0;
always @(posedge clk) v$FF0_9402_out0 <= v$G12_2216_out0;
always @(posedge clk) v$FF2_9418_out0 <= v$STATUSREAD_1637_out0;
always @(posedge clk) v$FF2_9419_out0 <= v$STATUSREAD_1638_out0;
always @(posedge clk) v$FF1_9422_out0 <= v$ShiftEN_7722_out0 ? v$MUX1_416_out0 : v$FF1_9422_out0;
always @(posedge clk) v$FF1_9423_out0 <= v$ShiftEN_7723_out0 ? v$MUX1_417_out0 : v$FF1_9423_out0;
always @(posedge clk) v$FF1_9607_out0 <= v$CLK4_17983_out0 ? v$MUX2_6685_out0 : v$FF1_9607_out0;
always @(posedge clk) v$FF1_9608_out0 <= v$CLK4_17984_out0 ? v$MUX2_6686_out0 : v$FF1_9608_out0;
always @(posedge clk) v$REG11_9622_out0 <= v$HALT1_4159_out0 ? v$DATAIN1_9634_out0 : v$REG11_9622_out0;
always @(posedge clk) v$FF1_9630_out0 <= v$G2_5253_out0;
always @(posedge clk) v$FF1_9631_out0 <= v$G2_5254_out0;
always @(posedge clk) v$FF3_9971_out0 <= v$SHIFTEN_9406_out0 ? v$MUX5_9524_out0 : v$FF3_9971_out0;
always @(posedge clk) v$FF3_9972_out0 <= v$SHIFTEN_9407_out0 ? v$MUX5_9525_out0 : v$FF3_9972_out0;
always @(posedge clk) v$FF3_9973_out0 <= v$SHIFTEN_9408_out0 ? v$MUX5_9526_out0 : v$FF3_9973_out0;
always @(posedge clk) v$FF3_9974_out0 <= v$SHIFTEN_9409_out0 ? v$MUX5_9527_out0 : v$FF3_9974_out0;
always @(posedge clk) v$FF3_9975_out0 <= v$SHIFTEN_9410_out0 ? v$MUX5_9528_out0 : v$FF3_9975_out0;
always @(posedge clk) v$FF3_9976_out0 <= v$SHIFTEN_9411_out0 ? v$MUX5_9529_out0 : v$FF3_9976_out0;
always @(posedge clk) v$FF3_9977_out0 <= v$SHIFTEN_9412_out0 ? v$MUX5_9530_out0 : v$FF3_9977_out0;
always @(posedge clk) v$FF3_9978_out0 <= v$SHIFTEN_9413_out0 ? v$MUX5_9531_out0 : v$FF3_9978_out0;
always @(posedge clk) v$FF3_9979_out0 <= v$SHIFTEN_9414_out0 ? v$MUX5_9532_out0 : v$FF3_9979_out0;
always @(posedge clk) v$FF3_9980_out0 <= v$SHIFTEN_9415_out0 ? v$MUX5_9533_out0 : v$FF3_9980_out0;
always @(posedge clk) v$FF3_9981_out0 <= v$SHIFTEN_9416_out0 ? v$MUX5_9534_out0 : v$FF3_9981_out0;
always @(posedge clk) v$FF3_9982_out0 <= v$SHIFTEN_9417_out0 ? v$MUX5_9535_out0 : v$FF3_9982_out0;
always @(posedge clk) v$REG1_10302_out0 <= v$EXEC2_8048_out0 ? v$MUX6_13706_out0 : v$REG1_10302_out0;
always @(posedge clk) v$REG1_10303_out0 <= v$EXEC2_8049_out0 ? v$MUX6_13707_out0 : v$REG1_10303_out0;
always @(posedge clk) v$FF1_10306_out0 <= v$G5_7583_out0 ? v$A1_9430_out1 : v$FF1_10306_out0;
always @(posedge clk) v$FF1_10307_out0 <= v$G5_7584_out0 ? v$A1_9431_out1 : v$FF1_10307_out0;
always @(posedge clk) v$FF8_10337_out0 <= v$EQ3_4203_out0;
always @(posedge clk) v$FF8_10338_out0 <= v$EQ3_4204_out0;
always @(posedge clk) v$FF9_10664_out0 <= v$STP$DECODED_16534_out0;
always @(posedge clk) v$FF9_10665_out0 <= v$STP$DECODED_16535_out0;
always @(posedge clk) v$REG4_10777_out0 <= v$START_3700_out0 ? v$RD_11793_out0 : v$REG4_10777_out0;
always @(posedge clk) v$S$FF_10816_out0 <= v$EXEC2_1167_out0 ? v$S_10699_out0 : v$S$FF_10816_out0;
always @(posedge clk) v$S$FF_10817_out0 <= v$EXEC2_1168_out0 ? v$S_10700_out0 : v$S$FF_10817_out0;
always @(posedge clk) v$REG1_10904_out0 <= v$EXEC2_1469_out0 ? v$MUX5_7954_out0 : v$REG1_10904_out0;
always @(posedge clk) v$REG1_10905_out0 <= v$EXEC2_1470_out0 ? v$MUX5_7955_out0 : v$REG1_10905_out0;
always @(posedge clk) v$FF14_10906_out0 <= v$VALID_3712_out0;
always @(posedge clk) v$FF14_10907_out0 <= v$VALID_3713_out0;
always @(posedge clk) v$FF3_10915_out0 <= v$CLK4_17983_out0 ? v$MUX4_17084_out0 : v$FF3_10915_out0;
always @(posedge clk) v$FF3_10916_out0 <= v$CLK4_17984_out0 ? v$MUX4_17085_out0 : v$FF3_10916_out0;
always @(posedge clk) v$REG4_10994_out0 <= v$G88_7401_out0;
always @(posedge clk) v$REG3_11001_out0 <= v$D1_14097_out3 ? v$DIN3_14418_out0 : v$REG3_11001_out0;
always @(posedge clk) v$REG3_11002_out0 <= v$D1_14098_out3 ? v$DIN3_14419_out0 : v$REG3_11002_out0;
always @(posedge clk) v$FF1_11054_out0 <= v$G1_4213_out0;
always @(posedge clk) v$FF1_11055_out0 <= v$G1_4214_out0;
always @(posedge clk) v$REG3_11767_out0 <= v$G33_324_out0 ? v$SEL4_9556_out0 : v$REG3_11767_out0;
always @(posedge clk) v$REG3_11768_out0 <= v$G18_7510_out0 ? v$SEL4_9557_out0 : v$REG3_11768_out0;
always @(posedge clk) v$REG2_11798_out0 <= v$IR2$VALID_13250_out0 ? v$_8774_out0 : v$REG2_11798_out0;
always @(posedge clk) v$REG2_11799_out0 <= v$IR2$VALID_13251_out0 ? v$_8775_out0 : v$REG2_11799_out0;
always @(posedge clk) v$REG1_12089_out0 <= v$OUT_14931_out0;
always @(posedge clk) v$FF15_12716_out0 <= v$HALT$PREV$PREV_18074_out0;
always @(posedge clk) v$FF15_12717_out0 <= v$HALT$PREV$PREV_18075_out0;
always @(posedge clk) v$FF7_12756_out0 <= v$STALL_17890_out0;
always @(posedge clk) v$FF7_12757_out0 <= v$STALL_17891_out0;
always @(posedge clk) v$PCNORMAL_12768_out0 <= v$G33_10750_out0 ? v$SUM_13667_out0 : v$PCNORMAL_12768_out0;
always @(posedge clk) v$PCNORMAL_12769_out0 <= v$G33_10751_out0 ? v$SUM_13668_out0 : v$PCNORMAL_12769_out0;
v$RAM1_12913 I12913 (v$RAM1_12913_out0, v$RAMADDR_13607_out0, v$MUX2_15843_out0, v$RAMWEN_17961_out0, clk);
always @(posedge clk) v$FF2_13039_out0 <= v$G7_14122_out0;
always @(posedge clk) v$FF2_13040_out0 <= v$G7_14123_out0;
always @(posedge clk) v$FF2_13041_out0 <= v$G7_14124_out0;
always @(posedge clk) v$FF2_13042_out0 <= v$G7_14125_out0;
always @(posedge clk) v$FF2_13043_out0 <= v$G7_14126_out0;
always @(posedge clk) v$FF2_13044_out0 <= v$G7_14127_out0;
always @(posedge clk) v$FF2_13045_out0 <= v$G4_11833_out0;
always @(posedge clk) v$FF2_13046_out0 <= v$G4_11834_out0;
always @(posedge clk) v$FF2_13047_out0 <= v$G4_11835_out0;
always @(posedge clk) v$FF2_13048_out0 <= v$G4_11836_out0;
always @(posedge clk) v$FF2_13049_out0 <= v$G4_11837_out0;
always @(posedge clk) v$FF2_13050_out0 <= v$G7_14128_out0;
always @(posedge clk) v$FF2_13051_out0 <= v$G7_14129_out0;
always @(posedge clk) v$FF2_13052_out0 <= v$G7_14130_out0;
always @(posedge clk) v$FF2_13053_out0 <= v$G7_14131_out0;
always @(posedge clk) v$FF2_13054_out0 <= v$G7_14132_out0;
always @(posedge clk) v$FF2_13055_out0 <= v$G7_14133_out0;
always @(posedge clk) v$FF2_13056_out0 <= v$G4_11838_out0;
always @(posedge clk) v$FF2_13057_out0 <= v$G4_11839_out0;
always @(posedge clk) v$FF2_13058_out0 <= v$G4_11840_out0;
always @(posedge clk) v$FF2_13059_out0 <= v$G4_11841_out0;
always @(posedge clk) v$FF2_13060_out0 <= v$G4_11842_out0;
always @(posedge clk) v$FF1_13095_out0 <= v$G16_6391_out0 ? v$G7_1831_out0 : v$FF1_13095_out0;
always @(posedge clk) v$FF1_13096_out0 <= v$G16_6392_out0 ? v$G7_1832_out0 : v$FF1_13096_out0;
always @(posedge clk) v$FF2_13458_out0 <= v$G51_18762_out0;
always @(posedge clk) v$FF4_13548_out0 <= v$G54_13285_out0;
always @(posedge clk) v$REG1_13592_out0 <= v$MUX1_18328_out0;
always @(posedge clk) v$REG1_13593_out0 <= v$MUX1_18329_out0;
always @(posedge clk) v$FF1_13680_out0 <= v$EXEC2_9439_out0 ? v$S_10347_out0 : v$FF1_13680_out0;
always @(posedge clk) v$FF1_13681_out0 <= v$EXEC2_9440_out0 ? v$S_10348_out0 : v$FF1_13681_out0;
always @(posedge clk) v$REG1_14090_out0 <= v$G1_12223_out0 ? v$MUX1_5137_out0 : v$REG1_14090_out0;
always @(posedge clk) v$REG1_14099_out0 <= v$IR1$VALID_61_out0 ? v$RM_18197_out0 : v$REG1_14099_out0;
always @(posedge clk) v$REG1_14100_out0 <= v$IR1$VALID_62_out0 ? v$RM_18198_out0 : v$REG1_14100_out0;
always @(posedge clk) v$FF10_14203_out0 <= v$WREN_10997_out0;
always @(posedge clk) v$FF10_14204_out0 <= v$WREN_10998_out0;
always @(posedge clk) v$FF8_14460_out0 <= v$SHIFTEN_9406_out0 ? v$MUX4_16847_out0 : v$FF8_14460_out0;
always @(posedge clk) v$FF8_14461_out0 <= v$SHIFTEN_9407_out0 ? v$MUX4_16848_out0 : v$FF8_14461_out0;
always @(posedge clk) v$FF8_14462_out0 <= v$SHIFTEN_9408_out0 ? v$MUX4_16849_out0 : v$FF8_14462_out0;
always @(posedge clk) v$FF8_14463_out0 <= v$SHIFTEN_9409_out0 ? v$MUX4_16850_out0 : v$FF8_14463_out0;
always @(posedge clk) v$FF8_14464_out0 <= v$SHIFTEN_9410_out0 ? v$MUX4_16851_out0 : v$FF8_14464_out0;
always @(posedge clk) v$FF8_14465_out0 <= v$SHIFTEN_9411_out0 ? v$MUX4_16852_out0 : v$FF8_14465_out0;
always @(posedge clk) v$FF8_14466_out0 <= v$SHIFTEN_9412_out0 ? v$MUX4_16853_out0 : v$FF8_14466_out0;
always @(posedge clk) v$FF8_14467_out0 <= v$SHIFTEN_9413_out0 ? v$MUX4_16854_out0 : v$FF8_14467_out0;
always @(posedge clk) v$FF8_14468_out0 <= v$SHIFTEN_9414_out0 ? v$MUX4_16855_out0 : v$FF8_14468_out0;
always @(posedge clk) v$FF8_14469_out0 <= v$SHIFTEN_9415_out0 ? v$MUX4_16856_out0 : v$FF8_14469_out0;
always @(posedge clk) v$FF8_14470_out0 <= v$SHIFTEN_9416_out0 ? v$MUX4_16857_out0 : v$FF8_14470_out0;
always @(posedge clk) v$FF8_14471_out0 <= v$SHIFTEN_9417_out0 ? v$MUX4_16858_out0 : v$FF8_14471_out0;
always @(posedge clk) v$FF7_14553_out0 <= v$Shift_9605_out0 ? v$FF6_8963_out0 : v$FF7_14553_out0;
always @(posedge clk) v$FF7_14554_out0 <= v$Shift_9606_out0 ? v$FF6_8964_out0 : v$FF7_14554_out0;
always @(posedge clk) v$FF2_14629_out0 <= v$CLK4_12213_out0 ? v$G24_9618_out0 : v$FF2_14629_out0;
always @(posedge clk) v$FF2_14630_out0 <= v$CLK4_12214_out0 ? v$G24_9619_out0 : v$FF2_14630_out0;
always @(posedge clk) v$FF2_14782_out0 <= v$SHIFTEN_9406_out0 ? v$MUX6_10388_out0 : v$FF2_14782_out0;
always @(posedge clk) v$FF2_14783_out0 <= v$SHIFTEN_9407_out0 ? v$MUX6_10389_out0 : v$FF2_14783_out0;
always @(posedge clk) v$FF2_14784_out0 <= v$SHIFTEN_9408_out0 ? v$MUX6_10390_out0 : v$FF2_14784_out0;
always @(posedge clk) v$FF2_14785_out0 <= v$SHIFTEN_9409_out0 ? v$MUX6_10391_out0 : v$FF2_14785_out0;
always @(posedge clk) v$FF2_14786_out0 <= v$SHIFTEN_9410_out0 ? v$MUX6_10392_out0 : v$FF2_14786_out0;
always @(posedge clk) v$FF2_14787_out0 <= v$SHIFTEN_9411_out0 ? v$MUX6_10393_out0 : v$FF2_14787_out0;
always @(posedge clk) v$FF2_14788_out0 <= v$SHIFTEN_9412_out0 ? v$MUX6_10394_out0 : v$FF2_14788_out0;
always @(posedge clk) v$FF2_14789_out0 <= v$SHIFTEN_9413_out0 ? v$MUX6_10395_out0 : v$FF2_14789_out0;
always @(posedge clk) v$FF2_14790_out0 <= v$SHIFTEN_9414_out0 ? v$MUX6_10396_out0 : v$FF2_14790_out0;
always @(posedge clk) v$FF2_14791_out0 <= v$SHIFTEN_9415_out0 ? v$MUX6_10397_out0 : v$FF2_14791_out0;
always @(posedge clk) v$FF2_14792_out0 <= v$SHIFTEN_9416_out0 ? v$MUX6_10398_out0 : v$FF2_14792_out0;
always @(posedge clk) v$FF2_14793_out0 <= v$SHIFTEN_9417_out0 ? v$MUX6_10399_out0 : v$FF2_14793_out0;
always @(posedge clk) v$REG1_14834_out0 <= v$MUX1_9915_out0;
always @(posedge clk) v$REG1_14835_out0 <= v$MUX1_9916_out0;
always @(posedge clk) v$REG2_15005_out0 <= v$R_18353_out0;
always @(posedge clk) v$REG2_15006_out0 <= v$R_18354_out0;
always @(posedge clk) v$FF3_15030_out0 <= v$INTERRUPT2_1663_out0;
always @(posedge clk) v$FF3_15031_out0 <= v$INTERRUPT2_1664_out0;
always @(posedge clk) v$FF6_15324_out0 <= v$ShiftEN_7722_out0 ? v$MUX6_9130_out0 : v$FF6_15324_out0;
always @(posedge clk) v$FF6_15325_out0 <= v$ShiftEN_7723_out0 ? v$MUX6_9131_out0 : v$FF6_15325_out0;
always @(posedge clk) v$FF2_15481_out0 <= v$G1_5421_out0;
always @(posedge clk) v$FF2_15482_out0 <= v$G1_5422_out0;
always @(posedge clk) v$REG2_15617_out0 <= v$G13_7894_out0 ? v$B_3366_out0 : v$REG2_15617_out0;
always @(posedge clk) v$REG2_15618_out0 <= v$G13_7895_out0 ? v$B_3367_out0 : v$REG2_15618_out0;
always @(posedge clk) v$INT0_15885_out0 <= v$I0EN_8042_out0 ? v$SEL1_11971_out0 : v$INT0_15885_out0;
always @(posedge clk) v$INT0_15886_out0 <= v$I0EN_8043_out0 ? v$SEL1_11972_out0 : v$INT0_15886_out0;
always @(posedge clk) v$FF3_15956_out0 <= v$CLK4_12213_out0 ? v$G32_16334_out0 : v$FF3_15956_out0;
always @(posedge clk) v$FF3_15957_out0 <= v$CLK4_12214_out0 ? v$G32_16335_out0 : v$FF3_15957_out0;
always @(posedge clk) v$FF4_15974_out0 <= v$SHIFTEN_9406_out0 ? v$MUX2_13819_out0 : v$FF4_15974_out0;
always @(posedge clk) v$FF4_15975_out0 <= v$SHIFTEN_9407_out0 ? v$MUX2_13820_out0 : v$FF4_15975_out0;
always @(posedge clk) v$FF4_15976_out0 <= v$SHIFTEN_9408_out0 ? v$MUX2_13821_out0 : v$FF4_15976_out0;
always @(posedge clk) v$FF4_15977_out0 <= v$SHIFTEN_9409_out0 ? v$MUX2_13822_out0 : v$FF4_15977_out0;
always @(posedge clk) v$FF4_15978_out0 <= v$SHIFTEN_9410_out0 ? v$MUX2_13823_out0 : v$FF4_15978_out0;
always @(posedge clk) v$FF4_15979_out0 <= v$SHIFTEN_9411_out0 ? v$MUX2_13824_out0 : v$FF4_15979_out0;
always @(posedge clk) v$FF4_15980_out0 <= v$SHIFTEN_9412_out0 ? v$MUX2_13825_out0 : v$FF4_15980_out0;
always @(posedge clk) v$FF4_15981_out0 <= v$SHIFTEN_9413_out0 ? v$MUX2_13826_out0 : v$FF4_15981_out0;
always @(posedge clk) v$FF4_15982_out0 <= v$SHIFTEN_9414_out0 ? v$MUX2_13827_out0 : v$FF4_15982_out0;
always @(posedge clk) v$FF4_15983_out0 <= v$SHIFTEN_9415_out0 ? v$MUX2_13828_out0 : v$FF4_15983_out0;
always @(posedge clk) v$FF4_15984_out0 <= v$SHIFTEN_9416_out0 ? v$MUX2_13829_out0 : v$FF4_15984_out0;
always @(posedge clk) v$FF4_15985_out0 <= v$SHIFTEN_9417_out0 ? v$MUX2_13830_out0 : v$FF4_15985_out0;
always @(posedge clk) v$FF9_16021_out0 <= v$FF10_14203_out0 ? v$G26_16019_out0 : v$FF9_16021_out0;
always @(posedge clk) v$FF9_16022_out0 <= v$FF10_14204_out0 ? v$G26_16020_out0 : v$FF9_16022_out0;
always @(posedge clk) v$FF1_16074_out0 <= v$SHIFTEN_9406_out0 ? v$MUX7_17903_out0 : v$FF1_16074_out0;
always @(posedge clk) v$FF1_16075_out0 <= v$SHIFTEN_9407_out0 ? v$MUX7_17904_out0 : v$FF1_16075_out0;
always @(posedge clk) v$FF1_16076_out0 <= v$SHIFTEN_9408_out0 ? v$MUX7_17905_out0 : v$FF1_16076_out0;
always @(posedge clk) v$FF1_16077_out0 <= v$SHIFTEN_9409_out0 ? v$MUX7_17906_out0 : v$FF1_16077_out0;
always @(posedge clk) v$FF1_16078_out0 <= v$SHIFTEN_9410_out0 ? v$MUX7_17907_out0 : v$FF1_16078_out0;
always @(posedge clk) v$FF1_16079_out0 <= v$SHIFTEN_9411_out0 ? v$MUX7_17908_out0 : v$FF1_16079_out0;
always @(posedge clk) v$FF1_16080_out0 <= v$SHIFTEN_9412_out0 ? v$MUX7_17909_out0 : v$FF1_16080_out0;
always @(posedge clk) v$FF1_16081_out0 <= v$SHIFTEN_9413_out0 ? v$MUX7_17910_out0 : v$FF1_16081_out0;
always @(posedge clk) v$FF1_16082_out0 <= v$SHIFTEN_9414_out0 ? v$MUX7_17911_out0 : v$FF1_16082_out0;
always @(posedge clk) v$FF1_16083_out0 <= v$SHIFTEN_9415_out0 ? v$MUX7_17912_out0 : v$FF1_16083_out0;
always @(posedge clk) v$FF1_16084_out0 <= v$SHIFTEN_9416_out0 ? v$MUX7_17913_out0 : v$FF1_16084_out0;
always @(posedge clk) v$FF1_16085_out0 <= v$SHIFTEN_9417_out0 ? v$MUX7_17914_out0 : v$FF1_16085_out0;
always @(posedge clk) v$REG9_16088_out0 <= v$HALT0_361_out0 ? v$RAMADDR0_16982_out0 : v$REG9_16088_out0;
always @(posedge clk) v$FF6_16171_out0 <= v$PHALT1_8934_out0;
always @(posedge clk) v$FF1_16187_out0 <= v$Shift_9605_out0 ? v$FF2_1572_out0 : v$FF1_16187_out0;
always @(posedge clk) v$FF1_16188_out0 <= v$Shift_9606_out0 ? v$FF2_1573_out0 : v$FF1_16188_out0;
always @(posedge clk) v$REG0_16254_out0 <= v$D1_14097_out0 ? v$DIN3_14418_out0 : v$REG0_16254_out0;
always @(posedge clk) v$REG0_16255_out0 <= v$D1_14098_out0 ? v$DIN3_14419_out0 : v$REG0_16255_out0;
always @(posedge clk) v$FF1_16315_out0 <= v$EXEC2_1469_out0 ? v$S_10442_out0 : v$FF1_16315_out0;
always @(posedge clk) v$FF1_16316_out0 <= v$EXEC2_1470_out0 ? v$S_10443_out0 : v$FF1_16316_out0;
always @(posedge clk) v$FF2_16336_out0 <= v$CAPTURE_242_out0 ? v$G1_13546_out0 : v$FF2_16336_out0;
always @(posedge clk) v$FF2_16337_out0 <= v$CAPTURE_243_out0 ? v$G1_13547_out0 : v$FF2_16337_out0;
always @(posedge clk) v$FF5_16338_out0 <= v$ShiftEN_7722_out0 ? v$MUX5_18559_out0 : v$FF5_16338_out0;
always @(posedge clk) v$FF5_16339_out0 <= v$ShiftEN_7723_out0 ? v$MUX5_18560_out0 : v$FF5_16339_out0;
always @(posedge clk) v$REG2_16345_out0 <= v$THRESHOLD$WRITE_7236_out0 ? v$THRESHOLD_15533_out0 : v$REG2_16345_out0;
always @(posedge clk) v$REG2_16346_out0 <= v$THRESHOLD$WRITE_7237_out0 ? v$THRESHOLD_15534_out0 : v$REG2_16346_out0;
always @(posedge clk) v$FF5_16426_out0 <= v$PHALT0_11638_out0;
always @(posedge clk) v$FF12_16427_out0 <= v$FF10_7890_out0;
always @(posedge clk) v$FF12_16428_out0 <= v$FF10_7891_out0;
always @(posedge clk) v$REG10_16463_out0 <= v$HALT0_361_out0 ? v$DATAIN0_11058_out0 : v$REG10_16463_out0;
always @(posedge clk) v$FF2_16652_out0 <= v$INTERRUPT1_17700_out0;
always @(posedge clk) v$FF2_16653_out0 <= v$INTERRUPT1_17701_out0;
always @(posedge clk) v$FF8_16727_out0 <= v$Shift_9605_out0 ? v$FF4_8252_out0 : v$FF8_16727_out0;
always @(posedge clk) v$FF8_16728_out0 <= v$Shift_9606_out0 ? v$FF4_8253_out0 : v$FF8_16728_out0;
always @(posedge clk) v$REG2_16798_out0 <= v$_7380_out0;
v$ROM1_17450 I17450 (v$ROM1_17450_out0, v$ADDRESS_15194_out0, clk);
v$ROM1_17451 I17451 (v$ROM1_17451_out0, v$ADDRESS_15195_out0, clk);
always @(posedge clk) v$REG2_17480_out0 <= v$D1_14097_out2 ? v$DIN3_14418_out0 : v$REG2_17480_out0;
always @(posedge clk) v$REG2_17481_out0 <= v$D1_14098_out2 ? v$DIN3_14419_out0 : v$REG2_17481_out0;
always @(posedge clk) v$REG3_17753_out0 <= v$IR2$VALID_13250_out0 ? v$EQ1_16270_out0 : v$REG3_17753_out0;
always @(posedge clk) v$REG3_17754_out0 <= v$IR2$VALID_13251_out0 ? v$EQ1_16271_out0 : v$REG3_17754_out0;
always @(posedge clk) v$PCINTERRUPT_17807_out0 <= v$ININTERRUPT_1133_out0 ? v$SUM_13667_out0 : v$PCINTERRUPT_17807_out0;
always @(posedge clk) v$PCINTERRUPT_17808_out0 <= v$ININTERRUPT_1134_out0 ? v$SUM_13668_out0 : v$PCINTERRUPT_17808_out0;
always @(posedge clk) v$FF4_17846_out0 <= v$C1_5434_out0;
always @(posedge clk) v$FF4_17847_out0 <= v$C1_5435_out0;
always @(posedge clk) v$FF3_18116_out0 <= v$G29_7851_out0;
always @(posedge clk) v$FF3_18117_out0 <= v$G29_7852_out0;
always @(posedge clk) v$FF7_18120_out0 <= v$ShiftEN_7722_out0 ? v$MUX7_9480_out0 : v$FF7_18120_out0;
always @(posedge clk) v$FF7_18121_out0 <= v$ShiftEN_7723_out0 ? v$MUX7_9481_out0 : v$FF7_18121_out0;
always @(posedge clk) v$REG2_18373_out0 <= v$EXEC1_18513_out0 ? v$COUT$EXEC1_1594_out0 : v$REG2_18373_out0;
always @(posedge clk) v$FF4_18438_out0 <= v$INTERRUPT3_2816_out0;
always @(posedge clk) v$FF4_18439_out0 <= v$INTERRUPT3_2817_out0;
always @(posedge clk) v$FF5_18473_out0 <= v$Shift_9605_out0 ? v$FF3_1296_out0 : v$FF5_18473_out0;
always @(posedge clk) v$FF5_18474_out0 <= v$Shift_9606_out0 ? v$FF3_1297_out0 : v$FF5_18474_out0;
always @(posedge clk) v$LSB$FF_18514_out0 <= v$EXEC2_1167_out0 ? v$MUX5_17066_out0 : v$LSB$FF_18514_out0;
always @(posedge clk) v$LSB$FF_18515_out0 <= v$EXEC2_1168_out0 ? v$MUX5_17067_out0 : v$LSB$FF_18515_out0;
always @(posedge clk) v$INT1_18533_out0 <= v$I1EN_18402_out0 ? v$SEL1_11971_out0 : v$INT1_18533_out0;
always @(posedge clk) v$INT1_18534_out0 <= v$I1EN_18403_out0 ? v$SEL1_11972_out0 : v$INT1_18534_out0;
always @(posedge clk) v$FF13_18541_out0 <= v$FF7_12756_out0;
always @(posedge clk) v$FF13_18542_out0 <= v$FF7_12757_out0;
always @(posedge clk) v$REG1_18662_out0 <= v$MODEWRITE_14714_out0 ? v$SEL1_18247_out0 : v$REG1_18662_out0;
always @(posedge clk) v$REG1_18663_out0 <= v$MODEWRITE_14715_out0 ? v$SEL1_18248_out0 : v$REG1_18663_out0;
assign v$C9_18761_out0 = 16'h0;
assign v$C9_18760_out0 = 16'h0;
assign v$C3_18553_out0 = 1'h0;
assign v$C3_18552_out0 = 1'h0;
assign v$C3_18437_out0 = 24'h0;
assign v$C2_18321_out0 = 1'h0;
assign v$C2_18320_out0 = 1'h0;
assign v$CIN_18232_out0 = 1'h1;
assign v$CIN_18231_out0 = 1'h1;
assign v$CIN_18230_out0 = 1'h1;
assign v$CIN_18229_out0 = 1'h1;
assign v$CIN_18228_out0 = 1'h1;
assign v$CIN_18227_out0 = 1'h1;
assign v$CIN_18226_out0 = 1'h1;
assign v$CIN_18225_out0 = 1'h1;
assign v$C1_18209_out0 = 16'h0;
assign v$C1_18208_out0 = 16'h0;
assign v$C3_18130_out0 = 1'h0;
assign v$C3_18129_out0 = 1'h0;
assign v$C3_18128_out0 = 1'h0;
assign v$C2_18013_out0 = 15'h0;
assign v$C2_18012_out0 = 15'h0;
assign v$C4_17973_out0 = 24'h0;
assign v$C1_17673_out0 = 1'h0;
assign v$C1_17672_out0 = 1'h0;
assign v$C1_17671_out0 = 1'h0;
assign v$C1_17670_out0 = 1'h0;
assign v$C1_17669_out0 = 1'h0;
assign v$C1_17668_out0 = 1'h0;
assign v$C1_17667_out0 = 1'h0;
assign v$C1_17666_out0 = 1'h0;
assign v$C1_17341_out0 = 1'h1;
assign v$C1_17340_out0 = 1'h1;
assign v$C1_17339_out0 = 1'h1;
assign v$C1_17338_out0 = 1'h1;
assign v$C2_17021_out0 = 1'h0;
assign v$C2_17020_out0 = 1'h0;
assign v$C5_16919_out0 = 2'h2;
assign v$C5_16918_out0 = 2'h2;
assign v$C5_16917_out0 = 2'h2;
assign v$C5_16916_out0 = 2'h1;
assign v$C5_16915_out0 = 2'h2;
assign v$C5_16914_out0 = 2'h2;
assign v$C5_16913_out0 = 2'h2;
assign v$C5_16912_out0 = 2'h1;
assign v$C5_16911_out0 = 2'h2;
assign v$C5_16910_out0 = 1'h0;
assign v$C5_16909_out0 = 2'h2;
assign v$C5_16908_out0 = 1'h0;
assign v$C1_16843_out0 = 3'h0;
assign v$C1_16842_out0 = 3'h0;
assign v$C4_16518_out0 = 2'h1;
assign v$C4_16517_out0 = 2'h1;
assign v$C4_16516_out0 = 2'h1;
assign v$C4_16515_out0 = 2'h0;
assign v$C4_16514_out0 = 2'h1;
assign v$C4_16513_out0 = 2'h1;
assign v$C4_16512_out0 = 2'h1;
assign v$C4_16511_out0 = 2'h0;
assign v$C4_16510_out0 = 2'h1;
assign v$C4_16509_out0 = 2'h1;
assign v$CON4_16439_out0 = 1'h0;
assign v$CON4_16438_out0 = 1'h0;
assign v$CON4_16437_out0 = 1'h0;
assign v$CON4_16436_out0 = 1'h0;
assign v$CON4_16435_out0 = 1'h0;
assign v$C2_16332_out0 = 1'h1;
assign v$C2_16331_out0 = 1'h1;
assign v$C2_16330_out0 = 1'h1;
assign v$C2_16329_out0 = 1'h1;
assign v$C1_16323_out0 = 16'h0;
assign v$C1_16322_out0 = 16'h0;
assign v$C4_16303_out0 = 2'h0;
assign v$C4_16302_out0 = 2'h0;
assign v$C2_16284_out0 = 1'h0;
assign v$C2_16283_out0 = 1'h0;
assign v$C2_16282_out0 = 1'h0;
assign v$C2_16281_out0 = 1'h0;
assign v$C2_16241_out0 = 1'h1;
assign v$C2_16240_out0 = 1'h1;
assign v$C1_16234_out0 = 24'h0;
assign v$C1_16233_out0 = 24'h0;
assign v$C5_16095_out0 = 1'h0;
assign v$C2_15987_out0 = 6'h1;
assign v$C2_15986_out0 = 6'h1;
assign v$C1_15941_out0 = 12'h0;
assign v$C1_15940_out0 = 12'h0;
assign v$C1_15922_out0 = 1'h1;
assign v$C1_15921_out0 = 1'h1;
assign v$C4_15907_out0 = 12'h0;
assign v$C4_15906_out0 = 12'h0;
assign v$C1_15805_out0 = 11'h0;
assign v$C1_15804_out0 = 11'h0;
assign v$C1_15735_out0 = 5'h1f;
assign v$C1_15734_out0 = 5'h1f;
assign v$C1_15723_out0 = 1'h0;
assign v$C1_15722_out0 = 1'h0;
assign v$C1_15721_out0 = 1'h0;
assign v$C1_15720_out0 = 1'h0;
assign v$C1_15678_out0 = 5'h0;
assign v$C5_15620_out0 = 23'h0;
assign v$C5_15619_out0 = 23'h0;
assign v$C9_15265_out0 = 24'hffffff;
assign v$C9_15264_out0 = 24'hffffff;
assign v$C1_15227_out0 = 32'h0;
assign v$C1_15226_out0 = 32'h0;
assign v$C2_15181_out0 = 1'h0;
assign v$C2_15180_out0 = 1'h0;
assign v$C2_15179_out0 = 1'h0;
assign v$C2_15178_out0 = 1'h0;
assign v$C4_14833_out0 = 1'h1;
assign v$C4_14832_out0 = 1'h1;
assign v$C4_14831_out0 = 1'h1;
assign v$C4_14830_out0 = 1'h1;
assign v$C1_14813_out0 = 8'h0;
assign v$C1_14812_out0 = 8'h0;
assign v$C4_14657_out0 = 5'h0;
assign v$C7_14644_out0 = 24'h0;
assign v$C7_14643_out0 = 24'h0;
assign v$CON2_14371_out0 = 1'h0;
assign v$CON2_14370_out0 = 1'h0;
assign v$CON2_14369_out0 = 1'h0;
assign v$CON2_14368_out0 = 1'h0;
assign v$CON2_14367_out0 = 1'h0;
assign v$C1_14254_out0 = 2'h3;
assign v$C1_14253_out0 = 2'h3;
assign v$C1_14029_out0 = 1'h0;
assign v$C4_14027_out0 = 32'h0;
assign v$C4_14026_out0 = 32'h0;
assign v$C1_13992_out0 = 8'h0;
assign v$C1_13991_out0 = 8'h0;
assign v$C8_13622_out0 = 24'hffffff;
assign v$C8_13621_out0 = 24'hffffff;
assign v$C1_13581_out0 = 8'hff;
assign v$C1_13580_out0 = 5'h1f;
assign v$C1_13579_out0 = 8'hff;
assign v$C1_13578_out0 = 5'h1f;
assign v$C1_13577_out0 = 8'hff;
assign v$C1_13576_out0 = 5'h1f;
assign v$C1_13575_out0 = 8'hff;
assign v$C1_13574_out0 = 5'h1f;
assign v$C10_13541_out0 = 3'h0;
assign v$C10_13540_out0 = 3'h0;
assign v$C3_13519_out0 = 1'h1;
assign v$C3_13518_out0 = 1'h1;
assign v$C3_13517_out0 = 1'h1;
assign v$C3_13516_out0 = 1'h1;
assign v$C2_13510_out0 = 1'h0;
assign v$C2_13509_out0 = 1'h0;
assign v$C1_13449_out0 = 8'h0;
assign v$C1_13448_out0 = 8'h0;
assign v$C2_13387_out0 = 2'h1;
assign v$C2_13386_out0 = 2'h1;
assign v$C2_13326_out0 = 3'h0;
assign v$C2_13325_out0 = 3'h0;
assign v$C3_13164_out0 = 6'h0;
assign v$C3_13163_out0 = 6'h0;
assign v$CON6_13001_out0 = 1'h0;
assign v$CON6_13000_out0 = 1'h0;
assign v$CON6_12999_out0 = 1'h0;
assign v$CON6_12998_out0 = 1'h0;
assign v$CON6_12997_out0 = 1'h0;
assign v$C1_12853_out0 = 1'h0;
assign v$C1_12852_out0 = 1'h0;
assign v$C1_12826_out0 = 4'h0;
assign v$C1_12825_out0 = 4'h0;
assign v$C6_12552_out0 = 1'h1;
assign v$C6_12551_out0 = 1'h1;
assign v$C2_12208_out0 = 16'hffff;
assign v$C2_12207_out0 = 16'hffff;
assign v$C3_12206_out0 = 16'h0;
assign v$C3_12205_out0 = 16'h0;
assign v$C6_11361_out0 = 1'h0;
assign v$C6_11360_out0 = 1'h0;
assign v$C6_11359_out0 = 1'h0;
assign v$C6_11358_out0 = 1'h0;
assign v$C6_11357_out0 = 1'h0;
assign v$C6_11356_out0 = 1'h0;
assign v$C6_11355_out0 = 1'h0;
assign v$C6_11354_out0 = 1'h0;
assign v$C6_11353_out0 = 1'h0;
assign v$C6_11352_out0 = 1'h0;
assign v$C6_11351_out0 = 1'h0;
assign v$C6_11350_out0 = 1'h0;
assign v$C2_10701_out0 = 1'h1;
assign v$CON5_10685_out0 = 1'h0;
assign v$CON5_10684_out0 = 1'h0;
assign v$CON5_10683_out0 = 1'h0;
assign v$CON5_10682_out0 = 1'h0;
assign v$CON5_10681_out0 = 1'h0;
assign v$C2_10010_out0 = 16'hffff;
assign v$C2_10009_out0 = 16'hffff;
assign v$C7_9496_out0 = 1'h1;
assign v$C10_8950_out0 = 13'h0;
assign v$C10_8949_out0 = 13'h0;
assign v$C6_8836_out0 = 1'h0;
assign v$C5_8765_out0 = 1'h1;
assign v$C5_8764_out0 = 1'h1;
assign v$C5_8763_out0 = 1'h1;
assign v$C5_8762_out0 = 1'h1;
assign v$C4_8259_out0 = 31'h0;
assign v$C4_8258_out0 = 15'h0;
assign v$C4_8257_out0 = 31'h0;
assign v$C4_8256_out0 = 15'h0;
assign v$C8_8207_out0 = 13'h0;
assign v$C8_8206_out0 = 13'h0;
assign v$C6_8047_out0 = 6'h1;
assign v$C6_8046_out0 = 6'h1;
assign v$C1_7978_out0 = 8'h0;
assign v$C1_7977_out0 = 4'h0;
assign v$C1_7976_out0 = 2'h0;
assign v$C1_7975_out0 = 1'h0;
assign v$C1_7974_out0 = 8'h0;
assign v$C1_7973_out0 = 4'h0;
assign v$C1_7972_out0 = 2'h0;
assign v$C1_7971_out0 = 1'h0;
assign v$CON3_7916_out0 = 1'h0;
assign v$CON3_7915_out0 = 1'h0;
assign v$CON3_7914_out0 = 1'h0;
assign v$CON3_7913_out0 = 1'h0;
assign v$CON3_7912_out0 = 1'h0;
assign v$C2_7814_out0 = 24'h0;
assign v$C1_7725_out0 = 2'h2;
assign v$C1_7724_out0 = 2'h2;
assign v$C2_7631_out0 = 1'h1;
assign v$C2_7630_out0 = 1'h1;
assign v$C2_7629_out0 = 1'h1;
assign v$C2_7628_out0 = 1'h1;
assign v$C2_7627_out0 = 1'h1;
assign v$C2_7626_out0 = 1'h1;
assign v$C2_7625_out0 = 1'h1;
assign v$C2_7624_out0 = 1'h1;
assign v$C1_7425_out0 = 5'h0;
assign v$C1_7424_out0 = 5'h0;
assign v$C8_7282_out0 = 4'h0;
assign v$C8_7281_out0 = 4'h0;
assign v$C3_7014_out0 = 5'h17;
assign v$C4_6626_out0 = 3'h0;
assign v$C4_6625_out0 = 3'h0;
assign v$C6_6545_out0 = 2'h3;
assign v$C6_6544_out0 = 2'h3;
assign v$C6_6543_out0 = 2'h3;
assign v$C6_6542_out0 = 2'h2;
assign v$C6_6541_out0 = 2'h3;
assign v$C6_6540_out0 = 2'h3;
assign v$C6_6539_out0 = 2'h3;
assign v$C6_6538_out0 = 2'h2;
assign v$C6_6537_out0 = 2'h3;
assign v$C6_6536_out0 = 2'h2;
assign v$C6_6535_out0 = 2'h3;
assign v$C6_6534_out0 = 2'h2;
assign v$C1_6458_out0 = 1'h0;
assign v$C1_6457_out0 = 1'h0;
assign v$C10_6385_out0 = 16'h0;
assign v$C10_6384_out0 = 16'h0;
assign v$C4_6368_out0 = 1'h0;
assign v$C4_6367_out0 = 1'h0;
assign v$C7_6038_out0 = 13'h0;
assign v$C7_6037_out0 = 13'h0;
assign v$C1_6023_out0 = 2'h0;
assign v$C1_6022_out0 = 4'h0;
assign v$C1_6021_out0 = 1'h0;
assign v$C1_6020_out0 = 8'h0;
assign v$C1_6019_out0 = 16'h0;
assign v$C1_6018_out0 = 2'h0;
assign v$C1_6017_out0 = 4'h0;
assign v$C1_6016_out0 = 1'h0;
assign v$C1_6015_out0 = 8'h0;
assign v$C1_6014_out0 = 16'h0;
assign v$C1_6013_out0 = 2'h0;
assign v$C1_6012_out0 = 4'h0;
assign v$C1_6011_out0 = 1'h0;
assign v$C1_6010_out0 = 8'h0;
assign v$C1_6009_out0 = 16'h0;
assign v$C1_6008_out0 = 4'h0;
assign v$C1_6007_out0 = 1'h0;
assign v$C1_6006_out0 = 16'h0;
assign v$C1_6005_out0 = 2'h0;
assign v$C1_6004_out0 = 8'h0;
assign v$C1_6003_out0 = 32'h0;
assign v$C1_6002_out0 = 4'h0;
assign v$C1_6001_out0 = 1'h0;
assign v$C1_6000_out0 = 16'h0;
assign v$C1_5999_out0 = 2'h0;
assign v$C1_5998_out0 = 8'h0;
assign v$C1_5997_out0 = 32'h0;
assign v$C1_5996_out0 = 2'h0;
assign v$C1_5995_out0 = 4'h0;
assign v$C1_5994_out0 = 1'h0;
assign v$C1_5993_out0 = 8'h0;
assign v$C1_5992_out0 = 16'h0;
assign v$C1_5991_out0 = 1'h0;
assign v$C1_5990_out0 = 2'h0;
assign v$C1_5989_out0 = 16'h0;
assign v$C1_5988_out0 = 4'h0;
assign v$C1_5987_out0 = 8'h0;
assign v$C1_5986_out0 = 1'h0;
assign v$C1_5985_out0 = 2'h0;
assign v$C1_5984_out0 = 4'h0;
assign v$C1_5983_out0 = 1'h0;
assign v$C1_5982_out0 = 8'h0;
assign v$C1_5981_out0 = 16'h0;
assign v$C1_5980_out0 = 2'h0;
assign v$C1_5979_out0 = 16'h0;
assign v$C1_5978_out0 = 4'h0;
assign v$C1_5977_out0 = 8'h0;
assign v$C1_5976_out0 = 1'h0;
assign v$C1_5975_out0 = 2'h0;
assign v$C1_5974_out0 = 4'h0;
assign v$C1_5973_out0 = 1'h0;
assign v$C1_5972_out0 = 8'h0;
assign v$C1_5971_out0 = 16'h0;
assign v$C1_5970_out0 = 2'h0;
assign v$C1_5969_out0 = 4'h0;
assign v$C1_5968_out0 = 1'h0;
assign v$C1_5967_out0 = 8'h0;
assign v$C1_5966_out0 = 16'h0;
assign v$C1_5965_out0 = 2'h0;
assign v$C1_5964_out0 = 4'h0;
assign v$C1_5963_out0 = 1'h0;
assign v$C1_5962_out0 = 8'h0;
assign v$C1_5961_out0 = 16'h0;
assign v$C1_5958_out0 = 8'h81;
assign v$C1_5957_out0 = 5'h11;
assign v$C1_5956_out0 = 8'h81;
assign v$C1_5955_out0 = 5'h11;
assign v$C1_5435_out0 = 1'h1;
assign v$C1_5434_out0 = 1'h1;
assign v$C1_5413_out0 = 4'h0;
assign v$C1_5412_out0 = 4'h0;
assign v$C3_5387_out0 = 1'h1;
assign v$C3_5386_out0 = 1'h1;
assign v$C1_5239_out0 = 5'h0;
assign v$C1_4468_out0 = 1'h0;
assign v$C1_4467_out0 = 1'h0;
assign v$C1_4466_out0 = 1'h0;
assign v$C1_4465_out0 = 1'h0;
assign v$C1_4464_out0 = 1'h0;
assign v$C1_4461_out0 = 24'h0;
assign v$C1_4460_out0 = 24'h0;
assign v$C1_4459_out0 = 24'h0;
assign v$C1_4458_out0 = 24'h0;
assign v$C1_4457_out0 = 24'h0;
assign v$C1_4456_out0 = 24'h0;
assign v$C1_4455_out0 = 24'h0;
assign v$C1_4454_out0 = 24'h0;
assign v$C1_4357_out0 = 1'h1;
assign v$C1_4356_out0 = 1'h1;
assign v$C5_4113_out0 = 32'h0;
assign v$C5_4112_out0 = 32'h0;
assign v$CON1_4084_out0 = 1'h0;
assign v$CON1_4083_out0 = 1'h0;
assign v$CON1_4082_out0 = 1'h0;
assign v$CON1_4081_out0 = 1'h0;
assign v$CON1_4080_out0 = 1'h0;
assign v$C5_3972_out0 = 24'h0;
assign v$C5_3971_out0 = 24'h0;
assign v$C5_3970_out0 = 24'h0;
assign v$C5_3969_out0 = 24'h0;
assign v$C5_3968_out0 = 24'h0;
assign v$C5_3967_out0 = 24'h0;
assign v$C5_3966_out0 = 24'h0;
assign v$C5_3965_out0 = 24'h0;
assign v$C5_3964_out0 = 24'h0;
assign v$C5_3963_out0 = 24'h0;
assign v$C5_3962_out0 = 24'h0;
assign v$C5_3961_out0 = 24'h0;
assign v$C4_3755_out0 = 1'h1;
assign v$C4_3754_out0 = 1'h1;
assign v$C11_3633_out0 = 1'h0;
assign v$C11_3632_out0 = 1'h0;
assign v$C2_3629_out0 = 1'h1;
assign v$C2_3628_out0 = 1'h1;
assign v$C3_3309_out0 = 2'h0;
assign v$C3_3308_out0 = 2'h0;
assign v$C3_3307_out0 = 2'h0;
assign v$C3_3306_out0 = 2'h0;
assign v$C3_3305_out0 = 2'h0;
assign v$C3_3304_out0 = 2'h0;
assign v$C3_3303_out0 = 2'h0;
assign v$C3_3302_out0 = 2'h0;
assign v$C9_3301_out0 = 16'h0;
assign v$C9_3300_out0 = 16'h0;
assign v$C1_3019_out0 = 2'h0;
assign v$C1_3018_out0 = 2'h0;
assign v$C2_2976_out0 = 1'h1;
assign v$C2_2975_out0 = 1'h1;
assign v$C4_2921_out0 = 1'h1;
assign v$C4_2920_out0 = 1'h1;
assign v$C2_2667_out0 = 1'h0;
assign v$C2_2666_out0 = 1'h0;
assign v$C1_2644_out0 = 1'h1;
assign v$C1_2643_out0 = 1'h1;
assign v$C1_2642_out0 = 1'h1;
assign v$C1_2641_out0 = 1'h1;
assign v$C1_2640_out0 = 1'h1;
assign v$C1_2639_out0 = 1'h1;
assign v$C1_2638_out0 = 1'h1;
assign v$C1_2637_out0 = 1'h1;
assign v$C1_2636_out0 = 1'h1;
assign v$C1_2635_out0 = 1'h1;
assign v$C1_2634_out0 = 1'h1;
assign v$C1_2633_out0 = 1'h1;
assign v$C4_2452_out0 = 13'h0;
assign v$C4_2451_out0 = 13'h0;
assign v$C6_2433_out0 = 1'h1;
assign v$C6_2432_out0 = 1'h1;
assign v$CON7_2424_out0 = 1'h0;
assign v$CON7_2423_out0 = 1'h0;
assign v$CON7_2422_out0 = 1'h0;
assign v$CON7_2421_out0 = 1'h0;
assign v$CON7_2420_out0 = 1'h0;
assign v$C7_1709_out0 = 16'h0;
assign v$C7_1708_out0 = 16'h0;
assign v$C6_1569_out0 = 1'h1;
assign v$C6_1568_out0 = 1'h1;
assign v$C1_1556_out0 = 8'hff;
assign v$C1_1555_out0 = 8'hff;
assign v$C6_1536_out0 = 13'h0;
assign v$C6_1535_out0 = 13'h0;
assign v$C1_1515_out0 = 1'h0;
assign v$C1_1514_out0 = 1'h0;
assign v$C1_1472_out0 = 1'h0;
assign v$C1_1471_out0 = 1'h0;
assign v$C2_1457_out0 = 1'h1;
assign v$C2_1456_out0 = 1'h1;
assign v$C3_1363_out0 = 1'h1;
assign v$C3_1362_out0 = 1'h1;
assign v$C2_1172_out0 = 1'h1;
assign v$C2_1171_out0 = 1'h1;
assign v$C7_339_out0 = 1'h0;
assign v$C7_338_out0 = 1'h0;
assign v$C2_165_out0 = 2'h0;
assign v$C2_164_out0 = 4'h0;
assign v$C2_163_out0 = 1'h0;
assign v$C2_162_out0 = 8'h0;
assign v$C2_161_out0 = 16'h0;
assign v$C2_160_out0 = 2'h0;
assign v$C2_159_out0 = 4'h0;
assign v$C2_158_out0 = 1'h0;
assign v$C2_157_out0 = 8'h0;
assign v$C2_156_out0 = 16'h0;
assign v$C2_155_out0 = 2'h0;
assign v$C2_154_out0 = 4'h0;
assign v$C2_153_out0 = 1'h0;
assign v$C2_152_out0 = 8'h0;
assign v$C2_151_out0 = 16'h0;
assign v$C2_150_out0 = 4'h0;
assign v$C2_149_out0 = 1'h0;
assign v$C2_148_out0 = 16'h0;
assign v$C2_147_out0 = 2'h0;
assign v$C2_146_out0 = 8'h0;
assign v$C2_145_out0 = 32'h0;
assign v$C2_144_out0 = 4'h0;
assign v$C2_143_out0 = 1'h0;
assign v$C2_142_out0 = 16'h0;
assign v$C2_141_out0 = 2'h0;
assign v$C2_140_out0 = 8'h0;
assign v$C2_139_out0 = 32'h0;
assign v$C2_138_out0 = 2'h0;
assign v$C2_137_out0 = 4'h0;
assign v$C2_136_out0 = 1'h0;
assign v$C2_135_out0 = 8'h0;
assign v$C2_134_out0 = 16'h0;
assign v$C2_133_out0 = 1'h0;
assign v$C2_132_out0 = 2'h0;
assign v$C2_131_out0 = 16'h0;
assign v$C2_130_out0 = 4'h0;
assign v$C2_129_out0 = 8'h0;
assign v$C2_128_out0 = 1'h0;
assign v$C2_127_out0 = 2'h0;
assign v$C2_126_out0 = 4'h0;
assign v$C2_125_out0 = 1'h0;
assign v$C2_124_out0 = 8'h0;
assign v$C2_123_out0 = 16'h0;
assign v$C2_122_out0 = 2'h0;
assign v$C2_121_out0 = 16'h0;
assign v$C2_120_out0 = 4'h0;
assign v$C2_119_out0 = 8'h0;
assign v$C2_118_out0 = 1'h0;
assign v$C2_117_out0 = 2'h0;
assign v$C2_116_out0 = 4'h0;
assign v$C2_115_out0 = 1'h0;
assign v$C2_114_out0 = 8'h0;
assign v$C2_113_out0 = 16'h0;
assign v$C2_112_out0 = 2'h0;
assign v$C2_111_out0 = 4'h0;
assign v$C2_110_out0 = 1'h0;
assign v$C2_109_out0 = 8'h0;
assign v$C2_108_out0 = 16'h0;
assign v$C2_107_out0 = 2'h0;
assign v$C2_106_out0 = 4'h0;
assign v$C2_105_out0 = 1'h0;
assign v$C2_104_out0 = 8'h0;
assign v$C2_103_out0 = 16'h0;
assign v$G3_20_out0 = !(v$FF0_5007_out0 || v$FF1_9630_out0);
assign v$G3_21_out0 = !(v$FF0_5008_out0 || v$FF1_9631_out0);
assign v$G2_65_out0 = ! v$FF1_191_out0;
assign v$G2_66_out0 = ! v$FF1_192_out0;
assign v$Q0_75_out0 = v$FF0_9401_out0;
assign v$Q0_76_out0 = v$FF0_9402_out0;
assign v$SIN_94_out0 = v$C7_338_out0;
assign v$SIN_100_out0 = v$C7_339_out0;
assign v$G58_168_out0 = ! v$FF5_4744_out0;
assign v$G58_169_out0 = ! v$FF5_4745_out0;
assign v$_1273_out0 = { v$FF0_9401_out0,v$FF1_2525_out0 };
assign v$_1274_out0 = { v$FF0_9402_out0,v$FF1_2526_out0 };
assign v$G2_1288_out0 = ((v$FF5_18473_out0 && !v$FF3_1296_out0) || (!v$FF5_18473_out0) && v$FF3_1296_out0);
assign v$G2_1289_out0 = ((v$FF5_18474_out0 && !v$FF3_1297_out0) || (!v$FF5_18474_out0) && v$FF3_1297_out0);
assign v$INITIAL$FETCH$OCCURRED_1537_out0 = v$FF4_17846_out0;
assign v$INITIAL$FETCH$OCCURRED_1538_out0 = v$FF4_17847_out0;
assign v$CIN$EXEC1_1591_out0 = v$REG2_18373_out0;
assign v$PHALT_1636_out0 = v$REG2_5128_out0;
assign v$SELOUT_1720_out0 = v$REG8_4106_out0;
assign v$SOUT1_1917_out0 = v$FF4_15974_out0;
assign v$SOUT1_1918_out0 = v$FF4_15975_out0;
assign v$SOUT1_1919_out0 = v$FF4_15976_out0;
assign v$SOUT1_1920_out0 = v$FF4_15977_out0;
assign v$SOUT1_1921_out0 = v$FF4_15978_out0;
assign v$SOUT1_1922_out0 = v$FF4_15979_out0;
assign v$SOUT1_1923_out0 = v$FF4_15980_out0;
assign v$SOUT1_1924_out0 = v$FF4_15981_out0;
assign v$SOUT1_1925_out0 = v$FF4_15982_out0;
assign v$SOUT1_1926_out0 = v$FF4_15983_out0;
assign v$SOUT1_1927_out0 = v$FF4_15984_out0;
assign v$SOUT1_1928_out0 = v$FF4_15985_out0;
assign v$I2P_2258_out0 = v$FF2_16336_out0;
assign v$I2P_2259_out0 = v$FF2_16337_out0;
assign v$_2264_out0 = { v$FF7_18120_out0,v$FF8_8026_out0 };
assign v$_2265_out0 = { v$FF7_18121_out0,v$FF8_8027_out0 };
assign v$PIPELINERESTART_2418_out0 = v$FF1_2_out0;
assign v$PIPELINERESTART_2419_out0 = v$FF1_3_out0;
assign v$G4_2889_out0 = ((v$FF7_14553_out0 && !v$FF6_8963_out0) || (!v$FF7_14553_out0) && v$FF6_8963_out0);
assign v$G4_2890_out0 = ((v$FF7_14554_out0 && !v$FF6_8964_out0) || (!v$FF7_14554_out0) && v$FF6_8964_out0);
assign v$LEFT$SHIT_3056_out0 = v$C1_17338_out0;
assign v$LEFT$SHIT_3057_out0 = v$C4_14830_out0;
assign v$LEFT$SHIT_3058_out0 = v$C3_13516_out0;
assign v$LEFT$SHIT_3059_out0 = v$C5_8762_out0;
assign v$LEFT$SHIT_3060_out0 = v$C2_16329_out0;
assign v$LEFT$SHIT_3066_out0 = v$C1_17339_out0;
assign v$LEFT$SHIT_3067_out0 = v$C4_14831_out0;
assign v$LEFT$SHIT_3068_out0 = v$C3_13517_out0;
assign v$LEFT$SHIT_3069_out0 = v$C5_8763_out0;
assign v$LEFT$SHIT_3070_out0 = v$C2_16330_out0;
assign v$LEFT$SHIT_3071_out0 = v$C1_14029_out0;
assign v$LEFT$SHIT_3077_out0 = v$C6_2432_out0;
assign v$LEFT$SHIT_3078_out0 = v$C4_14832_out0;
assign v$LEFT$SHIT_3079_out0 = v$C2_16331_out0;
assign v$LEFT$SHIT_3080_out0 = v$C5_8764_out0;
assign v$LEFT$SHIT_3081_out0 = v$C1_17340_out0;
assign v$LEFT$SHIT_3082_out0 = v$C3_13518_out0;
assign v$LEFT$SHIT_3083_out0 = v$C6_2433_out0;
assign v$LEFT$SHIT_3084_out0 = v$C4_14833_out0;
assign v$LEFT$SHIT_3085_out0 = v$C2_16332_out0;
assign v$LEFT$SHIT_3086_out0 = v$C5_8765_out0;
assign v$LEFT$SHIT_3087_out0 = v$C1_17341_out0;
assign v$LEFT$SHIT_3088_out0 = v$C3_13519_out0;
assign v$Q2_3149_out0 = v$FF2_15481_out0;
assign v$Q2_3150_out0 = v$FF2_15482_out0;
assign v$R0_3278_out0 = v$REG0_16254_out0;
assign v$R0_3279_out0 = v$REG0_16255_out0;
assign v$S$REG_3443_out0 = v$REG1_10904_out0;
assign v$S$REG_3444_out0 = v$REG1_10905_out0;
assign v$A$SAVED_3698_out0 = v$REG1_1163_out0;
assign v$A$SAVED_3699_out0 = v$REG1_1164_out0;
assign v$_3785_out0 = { v$FF7_14553_out0,v$FF6_8963_out0 };
assign v$_3786_out0 = { v$FF7_14554_out0,v$FF6_8964_out0 };
assign v$EN_3877_out0 = v$C7_9496_out0;
assign {v$A1_4011_out1,v$A1_4011_out0 } = v$REG1_14834_out0 + v$C2_15986_out0 + v$C1_1514_out0;
assign {v$A1_4012_out1,v$A1_4012_out0 } = v$REG1_14835_out0 + v$C2_15987_out0 + v$C1_1515_out0;
assign v$Q1_4450_out0 = v$FF1_9607_out0;
assign v$Q1_4451_out0 = v$FF1_9608_out0;
assign v$B$SAVED_4748_out0 = v$REG2_15617_out0;
assign v$B$SAVED_4749_out0 = v$REG2_15618_out0;
assign v$_4896_out0 = v$REG1_18662_out0[2:0];
assign v$_4896_out1 = v$REG1_18662_out0[3:1];
assign v$_4897_out0 = v$REG1_18663_out0[2:0];
assign v$_4897_out1 = v$REG1_18663_out0[3:1];
assign v$RESULT_5062_out0 = v$REG2_16798_out0;
assign v$Wordlength_5140_out0 = v$REG1_14834_out0 == 6'h27;
assign v$Wordlength_5141_out0 = v$REG1_14835_out0 == 6'h27;
assign v$G2_5253_out0 = ((v$FF0_5007_out0 && !v$FF1_9630_out0) || (!v$FF0_5007_out0) && v$FF1_9630_out0);
assign v$G2_5254_out0 = ((v$FF0_5008_out0 && !v$FF1_9631_out0) || (!v$FF0_5008_out0) && v$FF1_9631_out0);
assign v$OUT_5259_out0 = v$ROM1_17450_out0;
assign v$OUT_5260_out0 = v$ROM1_17451_out0;
assign v$Q2_5457_out0 = v$FF2_14629_out0;
assign v$Q2_5458_out0 = v$FF2_14630_out0;
assign v$G17_5476_out0 = ! v$FF2_16652_out0;
assign v$G17_5477_out0 = ! v$FF2_16653_out0;
assign v$D_5727_out0 = v$REG1_14090_out0;
assign v$STALL$PREV$CYCLE_5772_out0 = v$FF7_12756_out0;
assign v$STALL$PREV$CYCLE_5773_out0 = v$FF7_12757_out0;
assign v$STALL$PREV$PREV_5809_out0 = v$FF13_18541_out0;
assign v$STALL$PREV$PREV_5810_out0 = v$FF13_18542_out0;
assign v$IR$READ$IN$PREV$CYCLE_6188_out0 = v$REG2_15005_out0;
assign v$IR$READ$IN$PREV$CYCLE_6189_out0 = v$REG2_15006_out0;
assign v$I1P_6440_out0 = v$FF3_7563_out0;
assign v$I1P_6441_out0 = v$FF3_7564_out0;
assign v$EQ1_6932_out0 = v$REG2_16345_out0 == 16'h0;
assign v$EQ1_6933_out0 = v$REG2_16346_out0 == 16'h0;
assign v$PHALT1$PREV_7363_out0 = v$FF6_16171_out0;
assign v$G20_7402_out0 = ((v$FF7_18120_out0 && !v$FF8_8026_out0) || (!v$FF7_18120_out0) && v$FF8_8026_out0);
assign v$G20_7403_out0 = ((v$FF7_18121_out0 && !v$FF8_8027_out0) || (!v$FF7_18121_out0) && v$FF8_8027_out0);
assign v$PHALT0$PREV_7612_out0 = v$FF5_16426_out0;
assign v$HALT$PREV$PREV$PREV_7732_out0 = v$FF15_12716_out0;
assign v$HALT$PREV$PREV$PREV_7733_out0 = v$FF15_12717_out0;
assign v$_7734_out0 = { v$FF3_262_out0,v$FF4_2347_out0 };
assign v$_7735_out0 = { v$FF3_263_out0,v$FF4_2348_out0 };
assign v$LSB_7815_out0 = v$LSB$FF_18514_out0;
assign v$LSB_7816_out0 = v$LSB$FF_18515_out0;
assign v$LSBS_7937_out0 = v$REG1_10302_out0;
assign v$LSBS_7938_out0 = v$REG1_10303_out0;
assign v$R2_7958_out0 = v$REG2_17480_out0;
assign v$R2_7959_out0 = v$REG2_17481_out0;
assign v$B2_8415_out0 = v$C7_14643_out0;
assign v$B2_8418_out0 = v$C7_14644_out0;
assign v$CINA_8471_out0 = v$CON6_12997_out0;
assign v$CINA_8472_out0 = v$CON7_2420_out0;
assign v$CINA_8484_out0 = v$CON4_16435_out0;
assign v$CINA_8486_out0 = v$CON5_10681_out0;
assign v$CINA_8489_out0 = v$CON2_14367_out0;
assign v$CINA_8495_out0 = v$CON1_4080_out0;
assign v$CINA_8500_out0 = v$CON3_7912_out0;
assign v$CINA_8512_out0 = v$CON6_12998_out0;
assign v$CINA_8513_out0 = v$CON7_2421_out0;
assign v$CINA_8525_out0 = v$CON4_16436_out0;
assign v$CINA_8527_out0 = v$CON5_10682_out0;
assign v$CINA_8530_out0 = v$CON2_14368_out0;
assign v$CINA_8536_out0 = v$CON1_4081_out0;
assign v$CINA_8541_out0 = v$CON3_7913_out0;
assign v$CINA_8553_out0 = v$CON6_12999_out0;
assign v$CINA_8554_out0 = v$CON7_2422_out0;
assign v$CINA_8566_out0 = v$CON4_16437_out0;
assign v$CINA_8568_out0 = v$CON5_10683_out0;
assign v$CINA_8571_out0 = v$CON2_14369_out0;
assign v$CINA_8577_out0 = v$CON1_4082_out0;
assign v$CINA_8582_out0 = v$CON3_7914_out0;
assign v$CINA_8594_out0 = v$CON6_13000_out0;
assign v$CINA_8595_out0 = v$CON7_2423_out0;
assign v$CINA_8607_out0 = v$CON4_16438_out0;
assign v$CINA_8609_out0 = v$CON5_10684_out0;
assign v$CINA_8612_out0 = v$CON2_14370_out0;
assign v$CINA_8618_out0 = v$CON1_4083_out0;
assign v$CINA_8623_out0 = v$CON3_7915_out0;
assign v$CINA_8635_out0 = v$CON6_13001_out0;
assign v$CINA_8636_out0 = v$CON7_2424_out0;
assign v$CINA_8648_out0 = v$CON4_16439_out0;
assign v$CINA_8650_out0 = v$CON5_10685_out0;
assign v$CINA_8653_out0 = v$CON2_14371_out0;
assign v$CINA_8659_out0 = v$CON1_4084_out0;
assign v$CINA_8664_out0 = v$CON3_7916_out0;
assign v$PHALT1_8934_out0 = v$REG14_5459_out0;
assign v$I3P_8969_out0 = v$FF1_6149_out0;
assign v$I3P_8970_out0 = v$FF1_6150_out0;
assign v$G23_9360_out0 = ((v$FF1_9422_out0 && !v$FF2_2951_out0) || (!v$FF1_9422_out0) && v$FF2_2951_out0);
assign v$G23_9361_out0 = ((v$FF1_9423_out0 && !v$FF2_2952_out0) || (!v$FF1_9423_out0) && v$FF2_2952_out0);
assign v$SHIFTEN_9406_out0 = v$C1_2633_out0;
assign v$SHIFTEN_9407_out0 = v$C1_2634_out0;
assign v$SHIFTEN_9408_out0 = v$C1_2635_out0;
assign v$SHIFTEN_9409_out0 = v$C1_2636_out0;
assign v$SHIFTEN_9410_out0 = v$C1_2637_out0;
assign v$SHIFTEN_9411_out0 = v$C1_2638_out0;
assign v$SHIFTEN_9412_out0 = v$C1_2639_out0;
assign v$SHIFTEN_9413_out0 = v$C1_2640_out0;
assign v$SHIFTEN_9414_out0 = v$C1_2641_out0;
assign v$SHIFTEN_9415_out0 = v$C1_2642_out0;
assign v$SHIFTEN_9416_out0 = v$C1_2643_out0;
assign v$SHIFTEN_9417_out0 = v$C1_2644_out0;
assign v$_9436_out0 = { v$FF8_16727_out0,v$FF4_8252_out0 };
assign v$_9437_out0 = { v$FF8_16728_out0,v$FF4_8253_out0 };
assign v$RecievedParity_9538_out0 = v$FF7_8087_out0;
assign v$RecievedParity_9539_out0 = v$FF7_8088_out0;
assign v$G31_9632_out0 = ! v$FF4_18438_out0;
assign v$G31_9633_out0 = ! v$FF4_18439_out0;
assign v$G63_10019_out0 = ! v$FF8_10337_out0;
assign v$G63_10020_out0 = ! v$FF8_10338_out0;
assign v$I0P_10308_out0 = v$FF4_3781_out0;
assign v$I0P_10309_out0 = v$FF4_3782_out0;
assign v$OUTPUT_10339_out0 = v$FF1_5226_out0;
assign v$OUTPUT_10340_out0 = v$FF1_5227_out0;
assign v$OUTPUT_10341_out0 = v$FF1_5228_out0;
assign v$OUTPUT_10342_out0 = v$FF1_5229_out0;
assign v$HALT$PREV_10386_out0 = v$FF10_7890_out0;
assign v$HALT$PREV_10387_out0 = v$FF10_7891_out0;
assign v$R3_10746_out0 = v$REG3_11001_out0;
assign v$R3_10747_out0 = v$REG3_11002_out0;
assign v$Q1_10923_out0 = v$FF1_1178_out0;
assign v$Q1_10924_out0 = v$FF1_1179_out0;
assign v$PHALT0_11638_out0 = v$REG13_296_out0;
assign v$ISINTERRUPTED_11856_out0 = v$FF1_13095_out0;
assign v$ISINTERRUPTED_11857_out0 = v$FF1_13096_out0;
assign v$G21_11874_out0 = ((v$FF5_16338_out0 && !v$FF6_15324_out0) || (!v$FF5_16338_out0) && v$FF6_15324_out0);
assign v$G21_11875_out0 = ((v$FF5_16339_out0 && !v$FF6_15325_out0) || (!v$FF5_16339_out0) && v$FF6_15325_out0);
assign v$INT2_11881_out0 = v$C3_18130_out0;
assign v$G24_12087_out0 = ! v$FF3_15030_out0;
assign v$G24_12088_out0 = ! v$FF3_15031_out0;
assign v$LASTQ_12098_out0 = v$FF2_13039_out0;
assign v$LASTQ_12099_out0 = v$FF2_13040_out0;
assign v$LASTQ_12100_out0 = v$FF2_13041_out0;
assign v$LASTQ_12101_out0 = v$FF2_13042_out0;
assign v$LASTQ_12102_out0 = v$FF2_13043_out0;
assign v$LASTQ_12103_out0 = v$FF2_13044_out0;
assign v$LASTQ_12104_out0 = v$FF2_13045_out0;
assign v$LASTQ_12105_out0 = v$FF2_13046_out0;
assign v$LASTQ_12106_out0 = v$FF2_13047_out0;
assign v$LASTQ_12107_out0 = v$FF2_13048_out0;
assign v$LASTQ_12108_out0 = v$FF2_13049_out0;
assign v$LASTQ_12109_out0 = v$FF2_13050_out0;
assign v$LASTQ_12110_out0 = v$FF2_13051_out0;
assign v$LASTQ_12111_out0 = v$FF2_13052_out0;
assign v$LASTQ_12112_out0 = v$FF2_13053_out0;
assign v$LASTQ_12113_out0 = v$FF2_13054_out0;
assign v$LASTQ_12114_out0 = v$FF2_13055_out0;
assign v$LASTQ_12115_out0 = v$FF2_13056_out0;
assign v$LASTQ_12116_out0 = v$FF2_13057_out0;
assign v$LASTQ_12117_out0 = v$FF2_13058_out0;
assign v$LASTQ_12118_out0 = v$FF2_13059_out0;
assign v$LASTQ_12119_out0 = v$FF2_13060_out0;
assign v$PCHALT_12746_out0 = v$REG1_8824_out0;
assign v$LEFT$SHIFT_12832_out0 = v$C11_3632_out0;
assign v$LEFT$SHIFT_12833_out0 = v$C2_17020_out0;
assign v$LEFT$SHIFT_12834_out0 = v$C3_1362_out0;
assign v$LEFT$SHIFT_12835_out0 = v$C3_18128_out0;
assign v$LEFT$SHIFT_12836_out0 = v$C3_18129_out0;
assign v$LEFT$SHIFT_12837_out0 = v$C11_3633_out0;
assign v$LEFT$SHIFT_12838_out0 = v$C2_17021_out0;
assign v$LEFT$SHIFT_12839_out0 = v$C3_1363_out0;
assign v$RMORIGINAL_12978_out0 = v$REG1_14099_out0;
assign v$RMORIGINAL_12979_out0 = v$REG1_14100_out0;
assign v$G1_13147_out0 = ! v$FF0_5007_out0;
assign v$G1_13148_out0 = ! v$FF0_5008_out0;
assign v$VALID$PREV_13429_out0 = v$FF14_10906_out0;
assign v$VALID$PREV_13430_out0 = v$FF14_10907_out0;
assign v$CARRY_13442_out0 = v$FF1_10306_out0;
assign v$CARRY_13443_out0 = v$FF1_10307_out0;
assign v$Q0_13703_out0 = v$FF0_655_out0;
assign v$Q0_13704_out0 = v$FF0_656_out0;
assign v$R1_13766_out0 = v$REG1_4894_out0;
assign v$R1_13767_out0 = v$REG1_4895_out0;
assign v$B$SHIFTED_13792_out0 = v$REG1_12089_out0;
assign v$Q1_14326_out0 = v$FF1_2525_out0;
assign v$Q1_14327_out0 = v$FF1_2526_out0;
assign v$G1_14473_out0 = ! v$FF1_6026_out0;
assign v$G1_14474_out0 = ! v$FF1_6027_out0;
assign v$ADDRESS_14580_out0 = v$REG2_657_out0;
assign v$ADDRESS_14581_out0 = v$REG2_658_out0;
assign v$G5_14653_out0 = ((v$FF8_16727_out0 && !v$FF4_8252_out0) || (!v$FF8_16727_out0) && v$FF4_8252_out0);
assign v$G5_14654_out0 = ((v$FF8_16728_out0 && !v$FF4_8253_out0) || (!v$FF8_16728_out0) && v$FF4_8253_out0);
assign v$_14774_out0 = { v$FF1_9422_out0,v$FF2_2951_out0 };
assign v$_14775_out0 = { v$FF1_9423_out0,v$FF2_2952_out0 };
assign {v$A2_14825_out1,v$A2_14825_out0 } = v$REG2_657_out0 + v$C6_8046_out0 + v$C4_6367_out0;
assign {v$A2_14826_out1,v$A2_14826_out0 } = v$REG2_658_out0 + v$C6_8047_out0 + v$C4_6368_out0;
assign v$_14895_out0 = { v$FF1_16187_out0,v$FF2_1572_out0 };
assign v$_14896_out0 = { v$FF1_16188_out0,v$FF2_1573_out0 };
assign v$CIN_15050_out0 = v$C6_12551_out0;
assign v$CIN_15052_out0 = v$C5_16095_out0;
assign v$CIN_15053_out0 = v$C6_12552_out0;
assign v$G71_15274_out0 = ! v$FF4_8055_out0;
assign v$G71_15275_out0 = ! v$FF4_8056_out0;
assign v$LSBS_15316_out0 = v$REG1_8890_out0;
assign v$LSBS_15317_out0 = v$REG1_8891_out0;
assign v$EQ1_15322_out0 = v$REG1_14834_out0 == 6'h1e;
assign v$EQ1_15323_out0 = v$REG1_14835_out0 == 6'h1e;
assign v$SAVED_15383_out0 = v$REG3_6998_out0;
assign v$G3_15837_out0 = ((v$FF1_16187_out0 && !v$FF2_1572_out0) || (!v$FF1_16187_out0) && v$FF2_1572_out0);
assign v$G3_15838_out0 = ((v$FF1_16188_out0 && !v$FF2_1573_out0) || (!v$FF1_16188_out0) && v$FF2_1573_out0);
assign v$G52_15938_out0 = ! v$FF4_7017_out0;
assign v$G52_15939_out0 = ! v$FF4_7018_out0;
assign v$_15954_out0 = { v$FF5_16338_out0,v$FF6_15324_out0 };
assign v$_15955_out0 = { v$FF5_16339_out0,v$FF6_15325_out0 };
assign v$STATE_16013_out0 = v$FF1_5226_out0;
assign v$STATE_16014_out0 = v$FF1_5227_out0;
assign v$STATE_16015_out0 = v$FF1_5228_out0;
assign v$STATE_16016_out0 = v$FF1_5229_out0;
assign v$STATE_16017_out0 = v$REG1_7074_out0;
assign v$IR2_16559_out0 = v$REG4_6650_out0;
assign v$IR2_16560_out0 = v$REG4_6651_out0;
assign v$G24_17018_out0 = ((v$FF3_262_out0 && !v$FF4_2347_out0) || (!v$FF3_262_out0) && v$FF4_2347_out0);
assign v$G24_17019_out0 = ((v$FF3_263_out0 && !v$FF4_2348_out0) || (!v$FF3_263_out0) && v$FF4_2348_out0);
assign v$A_17045_out0 = v$REG1_13592_out0;
assign v$A_17046_out0 = v$REG1_13593_out0;
assign v$Q2_17486_out0 = v$FF2_4345_out0;
assign v$Q2_17487_out0 = v$FF2_4346_out0;
assign v$RD$OUT_17889_out0 = v$REG4_10777_out0;
assign v$B_17974_out0 = v$REG2_16345_out0;
assign v$B_17975_out0 = v$REG2_16346_out0;
assign v$HALT$PREV$PREV_18074_out0 = v$FF12_16427_out0;
assign v$HALT$PREV$PREV_18075_out0 = v$FF12_16428_out0;
assign v$INT3_18126_out0 = v$C2_18320_out0;
assign v$INT3_18127_out0 = v$C2_18321_out0;
assign v$SOUT_18193_out0 = v$FF1_9422_out0;
assign v$SOUT_18194_out0 = v$FF1_9423_out0;
assign v$AUTODISABLE_18213_out0 = v$FF3_18116_out0;
assign v$AUTODISABLE_18214_out0 = v$FF3_18117_out0;
assign v$Q3_18289_out0 = v$FF3_15956_out0;
assign v$Q3_18290_out0 = v$FF3_15957_out0;
assign v$EPARITY_18309_out0 = v$FF9_16021_out0;
assign v$EPARITY_18310_out0 = v$FF9_16022_out0;
assign v$Q0_18318_out0 = v$FF0_4326_out0;
assign v$Q0_18319_out0 = v$FF0_4327_out0;
assign v$_18410_out0 = { v$FF5_18473_out0,v$FF3_1296_out0 };
assign v$_18411_out0 = { v$FF5_18474_out0,v$FF3_1297_out0 };
assign v$Q3_18425_out0 = v$FF3_10915_out0;
assign v$Q3_18426_out0 = v$FF3_10916_out0;
assign v$_18459_out0 = v$REG1_4043_out0[3:0];
assign v$_18459_out1 = v$REG1_4043_out0[7:4];
assign v$_18460_out0 = v$REG1_4044_out0[3:0];
assign v$_18460_out1 = v$REG1_4044_out0[7:4];
assign v$OUTPUT_18477_out0 = v$REG1_7074_out0;
assign v$G1_33_out0 = v$Wordlength_5140_out0 || v$G2_65_out0;
assign v$G1_34_out0 = v$Wordlength_5141_out0 || v$G2_66_out0;
assign v$SIN_91_out0 = v$SOUT1_1918_out0;
assign v$SIN_92_out0 = v$SOUT1_1921_out0;
assign v$SIN_93_out0 = v$SOUT1_1922_out0;
assign v$SIN_95_out0 = v$SOUT1_1920_out0;
assign v$SIN_96_out0 = v$SOUT1_1917_out0;
assign v$SIN_97_out0 = v$SOUT1_1924_out0;
assign v$SIN_98_out0 = v$SOUT1_1927_out0;
assign v$SIN_99_out0 = v$SOUT1_1928_out0;
assign v$SIN_101_out0 = v$SOUT1_1926_out0;
assign v$SIN_102_out0 = v$SOUT1_1923_out0;
assign v$CALCULATING_1493_out0 = v$OUTPUT_10339_out0;
assign v$_1528_out0 = v$A_17045_out0[7:0];
assign v$_1528_out1 = v$A_17045_out0[15:8];
assign v$_1529_out0 = v$A_17046_out0[7:0];
assign v$_1529_out1 = v$A_17046_out0[15:8];
assign v$G1_1592_out0 = ! v$Q0_18318_out0;
assign v$G1_1593_out0 = ! v$Q0_18319_out0;
assign v$IR2_1750_out0 = v$IR2_16559_out0;
assign v$IR2_1751_out0 = v$IR2_16560_out0;
assign v$_1829_out0 = { v$Q0_18318_out0,v$Q1_4450_out0 };
assign v$_1830_out0 = { v$Q0_18319_out0,v$Q1_4451_out0 };
assign v$G8_2267_out0 = ! v$Q1_14326_out0;
assign v$G8_2268_out0 = ! v$Q1_14327_out0;
assign v$I1P_2514_out0 = v$I1P_6440_out0;
assign v$I1P_2515_out0 = v$I1P_6441_out0;
assign v$IR2_2933_out0 = v$IR2_16559_out0;
assign v$IR2_2934_out0 = v$IR2_16560_out0;
assign {v$A1_2938_out1,v$A1_2938_out0 } = v$D_5727_out0 + v$C1_5239_out0 + v$C2_10701_out0;
assign v$G18_2988_out0 = ! v$ISINTERRUPTED_11856_out0;
assign v$G18_2989_out0 = ! v$ISINTERRUPTED_11857_out0;
assign v$END4_3267_out0 = v$LASTQ_12108_out0;
assign v$END4_3268_out0 = v$LASTQ_12119_out0;
assign v$G6_3357_out0 = ((v$Q0_75_out0 && !v$Q1_14326_out0) || (!v$Q0_75_out0) && v$Q1_14326_out0);
assign v$G6_3358_out0 = ((v$Q0_76_out0 && !v$Q1_14327_out0) || (!v$Q0_76_out0) && v$Q1_14327_out0);
assign v$INTERRUPT3_3508_out0 = v$INT3_18126_out0;
assign v$INTERRUPT3_3509_out0 = v$INT3_18127_out0;
assign v$INTERRUPT2_3854_out0 = v$INT2_11881_out0;
assign v$B$SAVED_3884_out0 = v$B$SAVED_4748_out0;
assign v$B$SAVED_3885_out0 = v$B$SAVED_4749_out0;
assign v$CIN_3887_out0 = v$CIN$EXEC1_1591_out0;
assign v$_3985_out0 = v$B2_8415_out0[11:0];
assign v$_3985_out1 = v$B2_8415_out0[23:12];
assign v$_3988_out0 = v$B2_8418_out0[11:0];
assign v$_3988_out1 = v$B2_8418_out0[23:12];
assign v$OFF_4039_out0 = v$EQ1_6932_out0;
assign v$OFF_4040_out0 = v$EQ1_6933_out0;
assign v$G22_4313_out0 = ((v$Q1_10923_out0 && !v$Q0_13703_out0) || (!v$Q1_10923_out0) && v$Q0_13703_out0);
assign v$G22_4314_out0 = ((v$Q1_10924_out0 && !v$Q0_13704_out0) || (!v$Q1_10924_out0) && v$Q0_13704_out0);
assign v$G35_4315_out0 = v$Q1_4450_out0 && v$Q0_18318_out0;
assign v$G35_4316_out0 = v$Q1_4451_out0 && v$Q0_18319_out0;
assign v$I0P_4347_out0 = v$I0P_10308_out0;
assign v$I0P_4348_out0 = v$I0P_10309_out0;
assign v$B$SAVED_4358_out0 = v$B$SAVED_4748_out0;
assign v$B$SAVED_4359_out0 = v$B$SAVED_4749_out0;
assign v$G48_4876_out0 = ! v$STALL$PREV$CYCLE_5772_out0;
assign v$G48_4877_out0 = ! v$STALL$PREV$CYCLE_5773_out0;
assign v$G87_5144_out0 = ! v$PHALT0_11638_out0;
assign v$_5474_out0 = { v$_14774_out0,v$_7734_out0 };
assign v$_5475_out0 = { v$_14775_out0,v$_7735_out0 };
assign v$_5517_out0 = { v$_18410_out0,v$_14895_out0 };
assign v$_5518_out0 = { v$_18411_out0,v$_14896_out0 };
assign v$SERIALIN_5728_out0 = v$SOUT_18193_out0;
assign v$SERIALIN_5729_out0 = v$SOUT_18194_out0;
assign v$SEL6_5757_out0 = v$SAVED_15383_out0[35:12];
assign v$PIPELINE$RESTART_6071_out0 = v$PIPELINERESTART_2418_out0;
assign v$PIPELINE$RESTART_6072_out0 = v$PIPELINERESTART_2419_out0;
assign v$RECIEVEDPARITY_6224_out0 = v$RecievedParity_9538_out0;
assign v$RECIEVEDPARITY_6225_out0 = v$RecievedParity_9539_out0;
assign v$G64_6395_out0 = v$HALT$PREV_10386_out0 && v$STALL$PREV$PREV_5809_out0;
assign v$G64_6396_out0 = v$HALT$PREV_10387_out0 && v$STALL$PREV$PREV_5810_out0;
assign v$END1_6960_out0 = v$LASTQ_12107_out0;
assign v$END1_6961_out0 = v$LASTQ_12118_out0;
assign v$END1_6986_out0 = v$A2_14825_out1;
assign v$END1_6987_out0 = v$A2_14826_out1;
assign v$_7023_out0 = { v$_15954_out0,v$_2264_out0 };
assign v$_7024_out0 = { v$_15955_out0,v$_2265_out0 };
assign v$G22_7267_out0 = ((v$G21_11874_out0 && !v$G20_7402_out0) || (!v$G21_11874_out0) && v$G20_7402_out0);
assign v$G22_7268_out0 = ((v$G21_11875_out0 && !v$G20_7403_out0) || (!v$G21_11875_out0) && v$G20_7403_out0);
assign v$I2P_7492_out0 = v$I2P_2258_out0;
assign v$I2P_7493_out0 = v$I2P_2259_out0;
assign v$R3TEST_7537_out0 = v$R3_10746_out0;
assign v$R3TEST_7538_out0 = v$R3_10747_out0;
assign v$END6_7544_out0 = v$LASTQ_12102_out0;
assign v$END6_7545_out0 = v$LASTQ_12113_out0;
assign v$G2_7562_out0 = ! v$OUTPUT_18477_out0;
assign v$CALCULATING_7798_out0 = v$OUTPUT_10340_out0;
assign v$G7_7846_out0 = ! v$Q3_18289_out0;
assign v$G7_7847_out0 = ! v$Q3_18290_out0;
assign v$DM1_7858_out0 = v$SELOUT_1720_out0 ? 16'h0 : v$RAM1_12913_out0;
assign v$DM1_7858_out1 = v$SELOUT_1720_out0 ? v$RAM1_12913_out0 : 16'h0;
assign v$RXDISABLE_7888_out0 = v$_4896_out1;
assign v$RXDISABLE_7889_out0 = v$_4897_out1;
assign v$G3_8040_out0 = v$FF1_191_out0 || v$G2_65_out0;
assign v$G3_8041_out0 = v$FF1_192_out0 || v$G2_66_out0;
assign v$END_8096_out0 = v$A1_4011_out1;
assign v$END_8097_out0 = v$A1_4012_out1;
assign v$_8101_out0 = { v$_1273_out0,v$Q2_3149_out0 };
assign v$_8102_out0 = { v$_1274_out0,v$Q2_3150_out0 };
assign v$END4_8128_out0 = v$LASTQ_12099_out0;
assign v$END4_8129_out0 = v$LASTQ_12110_out0;
assign v$R0TEST_8236_out0 = v$R0_3278_out0;
assign v$R0TEST_8237_out0 = v$R0_3279_out0;
assign v$LEFT$SHIFT_8798_out0 = v$LEFT$SHIFT_12832_out0;
assign v$LEFT$SHIFT_8799_out0 = v$LEFT$SHIFT_12833_out0;
assign v$LEFT$SHIFT_8800_out0 = v$LEFT$SHIFT_12834_out0;
assign v$LEFT$SHIFT_8801_out0 = v$LEFT$SHIFT_12835_out0;
assign v$LEFT$SHIFT_8802_out0 = v$LEFT$SHIFT_12836_out0;
assign v$LEFT$SHIFT_8803_out0 = v$LEFT$SHIFT_12837_out0;
assign v$LEFT$SHIFT_8804_out0 = v$LEFT$SHIFT_12838_out0;
assign v$LEFT$SHIFT_8805_out0 = v$LEFT$SHIFT_12839_out0;
assign v$_8976_out0 = v$B_17974_out0[7:0];
assign v$_8976_out1 = v$B_17974_out0[15:8];
assign v$_8977_out0 = v$B_17975_out0[7:0];
assign v$_8977_out1 = v$B_17975_out0[15:8];
assign v$G6_9076_out0 = ! v$Q2_5457_out0;
assign v$G6_9077_out0 = ! v$Q2_5458_out0;
assign v$MODE_9126_out0 = v$_4896_out0;
assign v$MODE_9127_out0 = v$_4897_out0;
assign v$A$SAVED_9967_out0 = v$A$SAVED_3698_out0;
assign v$A$SAVED_9968_out0 = v$A$SAVED_3699_out0;
assign v$G38_10252_out0 = v$Q0_18318_out0 || v$Q1_4450_out0;
assign v$G38_10253_out0 = v$Q0_18319_out0 || v$Q1_4451_out0;
assign v$INIT_10752_out0 = v$G2_65_out0;
assign v$INIT_10753_out0 = v$G2_66_out0;
assign v$_10810_out0 = v$_18459_out0[1:0];
assign v$_10810_out1 = v$_18459_out0[3:2];
assign v$_10811_out0 = v$_18460_out0[1:0];
assign v$_10811_out1 = v$_18460_out0[3:2];
assign v$I3P_10827_out0 = v$I3P_8969_out0;
assign v$I3P_10828_out0 = v$I3P_8970_out0;
assign v$CARRY_10908_out0 = v$CARRY_13442_out0;
assign v$CARRY_10909_out0 = v$CARRY_13443_out0;
assign v$TXLast_11385_out0 = v$LASTQ_12104_out0;
assign v$TXLast_11386_out0 = v$LASTQ_12115_out0;
assign v$G57_11652_out0 = ! v$HALT$PREV_10386_out0;
assign v$G57_11653_out0 = ! v$HALT$PREV_10387_out0;
assign v$G27_11706_out0 = v$Q0_13703_out0 && v$Q1_10923_out0;
assign v$G27_11707_out0 = v$Q0_13704_out0 && v$Q1_10924_out0;
assign v$_11816_out0 = v$_18459_out1[1:0];
assign v$_11816_out1 = v$_18459_out1[3:2];
assign v$_11817_out0 = v$_18460_out1[1:0];
assign v$_11817_out1 = v$_18460_out1[3:2];
assign v$HALTED_11827_out0 = v$OUTPUT_10341_out0;
assign v$HALTED_11828_out0 = v$OUTPUT_10342_out0;
assign v$INSTR$READ1_11970_out0 = v$OUT_5260_out0;
assign v$SEL8_12749_out0 = v$SAVED_15383_out0[11:0];
assign v$RXlast_12821_out0 = v$LASTQ_12105_out0;
assign v$RXlast_12822_out0 = v$LASTQ_12116_out0;
assign v$RD$FPU_12947_out0 = v$RD$OUT_17889_out0;
assign v$G6_13009_out0 = ((v$G2_1288_out0 && !v$G3_15837_out0) || (!v$G2_1288_out0) && v$G3_15837_out0);
assign v$G6_13010_out0 = ((v$G2_1289_out0 && !v$G3_15838_out0) || (!v$G2_1289_out0) && v$G3_15838_out0);
assign v$_13410_out0 = { v$Q2_17486_out0,v$Q3_18425_out0 };
assign v$_13411_out0 = { v$Q2_17487_out0,v$Q3_18426_out0 };
assign v$G7_13431_out0 = ((v$G4_2889_out0 && !v$G5_14653_out0) || (!v$G4_2889_out0) && v$G5_14653_out0);
assign v$G7_13432_out0 = ((v$G4_2890_out0 && !v$G5_14654_out0) || (!v$G4_2890_out0) && v$G5_14654_out0);
assign v$G86_13527_out0 = ! v$PHALT1_8934_out0;
assign v$EVENPARITY_13588_out0 = v$EPARITY_18309_out0;
assign v$EVENPARITY_13589_out0 = v$EPARITY_18310_out0;
assign v$G4_13999_out0 = ! v$Q0_13703_out0;
assign v$G4_14000_out0 = ! v$Q0_13704_out0;
assign v$G51_14015_out0 = ! v$HALT$PREV_10386_out0;
assign v$G51_14016_out0 = ! v$HALT$PREV_10387_out0;
assign v$G25_14030_out0 = ((v$Q0_18318_out0 && !v$Q1_4450_out0) || (!v$Q0_18318_out0) && v$Q1_4450_out0);
assign v$G25_14031_out0 = ((v$Q0_18319_out0 && !v$Q1_4451_out0) || (!v$Q0_18319_out0) && v$Q1_4451_out0);
assign v$INSTR$READ0_14172_out0 = v$OUT_5259_out0;
assign v$G7_14311_out0 = ! v$Q2_3149_out0;
assign v$G7_14312_out0 = ! v$Q2_3150_out0;
assign v$A$SAVED_14631_out0 = v$A$SAVED_3698_out0;
assign v$A$SAVED_14632_out0 = v$A$SAVED_3699_out0;
assign v$PHALT_15137_out0 = v$PHALT_1636_out0;
assign v$R1TEST_15146_out0 = v$R1_13766_out0;
assign v$R1TEST_15147_out0 = v$R1_13767_out0;
assign v$R2TEST_15718_out0 = v$R2_7958_out0;
assign v$R2TEST_15719_out0 = v$R2_7959_out0;
assign v$G2_15761_out0 = ! v$Q1_4450_out0;
assign v$G2_15762_out0 = ! v$Q1_4451_out0;
assign v$G25_16104_out0 = ((v$G23_9360_out0 && !v$G24_17018_out0) || (!v$G23_9360_out0) && v$G24_17018_out0);
assign v$G25_16105_out0 = ((v$G23_9361_out0 && !v$G24_17019_out0) || (!v$G23_9361_out0) && v$G24_17019_out0);
assign v$_16127_out0 = { v$_3785_out0,v$_9436_out0 };
assign v$_16128_out0 = { v$_3786_out0,v$_9437_out0 };
assign v$G5_16154_out0 = ! v$Q1_10923_out0;
assign v$G5_16155_out0 = ! v$Q1_10924_out0;
v$AROM1_16158 I16158 (v$AROM1_16158_out0, v$ADDRESS_14580_out0);
v$AROM1_16159 I16159 (v$AROM1_16159_out0, v$ADDRESS_14581_out0);
assign v$G61_16446_out0 = ! v$HALT$PREV_10386_out0;
assign v$G61_16447_out0 = ! v$HALT$PREV_10387_out0;
assign v$G9_16494_out0 = ! v$Q0_75_out0;
assign v$G9_16495_out0 = ! v$Q0_76_out0;
assign v$PCHALT_16563_out0 = v$PCHALT_12746_out0;
assign v$CLK4_16733_out0 = v$G3_20_out0;
assign v$CLK4_16734_out0 = v$G3_21_out0;
assign v$END_17049_out0 = v$LASTQ_12106_out0;
assign v$END_17050_out0 = v$LASTQ_12117_out0;
assign v$CIN_17342_out0 = v$CIN_15050_out0;
assign v$CIN_17344_out0 = v$CIN_15052_out0;
assign v$CIN_17345_out0 = v$CIN_15053_out0;
assign v$G4_17586_out0 = ! v$Q3_18425_out0;
assign v$G4_17587_out0 = ! v$Q3_18426_out0;
assign v$increment_17844_out0 = v$EQ1_15322_out0;
assign v$increment_17845_out0 = v$EQ1_15323_out0;
assign v$G55_18199_out0 = ! v$HALT$PREV_10386_out0;
assign v$G55_18200_out0 = ! v$HALT$PREV_10387_out0;
assign v$_18326_out0 = { v$Q2_5457_out0,v$Q3_18289_out0 };
assign v$_18327_out0 = { v$Q2_5458_out0,v$Q3_18290_out0 };
assign v$G3_18414_out0 = ! v$Q2_17486_out0;
assign v$G3_18415_out0 = ! v$Q2_17487_out0;
assign v$G41_18479_out0 = v$Q0_18318_out0 && v$Q1_4450_out0;
assign v$G41_18480_out0 = v$Q0_18319_out0 && v$Q1_4451_out0;
assign v$_18518_out0 = { v$Q0_13703_out0,v$Q1_10923_out0 };
assign v$_18519_out0 = { v$Q0_13704_out0,v$Q1_10924_out0 };
assign v$NQ1_254_out0 = v$G5_16154_out0;
assign v$NQ1_255_out0 = v$G5_16155_out0;
assign v$SEL5_644_out0 = v$IR2_1750_out0[11:10];
assign v$SEL5_645_out0 = v$IR2_1751_out0[11:10];
assign v$G1_1195_out0 = ! v$OFF_4039_out0;
assign v$G1_1196_out0 = ! v$OFF_4040_out0;
assign v$_1218_out0 = v$_3985_out1[5:0];
assign v$_1218_out1 = v$_3985_out1[11:6];
assign v$_1221_out0 = v$_3988_out1[5:0];
assign v$_1221_out1 = v$_3988_out1[11:6];
assign v$NQ3_1491_out0 = v$G7_7846_out0;
assign v$NQ3_1492_out0 = v$G7_7847_out0;
assign v$_1523_out0 = v$_3985_out0[5:0];
assign v$_1523_out1 = v$_3985_out0[11:6];
assign v$_1526_out0 = v$_3988_out0[5:0];
assign v$_1526_out1 = v$_3988_out0[11:6];
assign v$MODE_1617_out0 = v$MODE_9126_out0;
assign v$MODE_1618_out0 = v$MODE_9127_out0;
assign v$IR2_2217_out0 = v$IR2_2933_out0;
assign v$IR2_2218_out0 = v$IR2_2934_out0;
assign v$_2345_out0 = v$_8976_out0[3:0];
assign v$_2345_out1 = v$_8976_out0[7:4];
assign v$_2346_out0 = v$_8977_out0[3:0];
assign v$_2346_out1 = v$_8977_out0[7:4];
assign v$G58_2518_out0 = v$FF11_2449_out0 && v$G57_11652_out0;
assign v$G58_2519_out0 = v$FF11_2450_out0 && v$G57_11653_out0;
assign v$_2897_out0 = v$_8976_out1[3:0];
assign v$_2897_out1 = v$_8976_out1[7:4];
assign v$_2898_out0 = v$_8977_out1[3:0];
assign v$_2898_out1 = v$_8977_out1[7:4];
assign v$NQ2_2980_out0 = v$G6_9076_out0;
assign v$NQ2_2981_out0 = v$G6_9077_out0;
assign v$NQ3_2998_out0 = v$G4_17586_out0;
assign v$NQ3_2999_out0 = v$G4_17587_out0;
assign v$LEFT$SHIT_3041_out0 = v$LEFT$SHIFT_8798_out0;
assign v$LEFT$SHIT_3042_out0 = v$LEFT$SHIFT_8798_out0;
assign v$LEFT$SHIT_3043_out0 = v$LEFT$SHIFT_8798_out0;
assign v$LEFT$SHIT_3044_out0 = v$LEFT$SHIFT_8798_out0;
assign v$LEFT$SHIT_3045_out0 = v$LEFT$SHIFT_8798_out0;
assign v$LEFT$SHIT_3046_out0 = v$LEFT$SHIFT_8799_out0;
assign v$LEFT$SHIT_3047_out0 = v$LEFT$SHIFT_8799_out0;
assign v$LEFT$SHIT_3048_out0 = v$LEFT$SHIFT_8799_out0;
assign v$LEFT$SHIT_3049_out0 = v$LEFT$SHIFT_8799_out0;
assign v$LEFT$SHIT_3050_out0 = v$LEFT$SHIFT_8799_out0;
assign v$LEFT$SHIT_3051_out0 = v$LEFT$SHIFT_8800_out0;
assign v$LEFT$SHIT_3052_out0 = v$LEFT$SHIFT_8800_out0;
assign v$LEFT$SHIT_3053_out0 = v$LEFT$SHIFT_8800_out0;
assign v$LEFT$SHIT_3054_out0 = v$LEFT$SHIFT_8800_out0;
assign v$LEFT$SHIT_3055_out0 = v$LEFT$SHIFT_8800_out0;
assign v$LEFT$SHIT_3061_out0 = v$LEFT$SHIFT_8801_out0;
assign v$LEFT$SHIT_3062_out0 = v$LEFT$SHIFT_8801_out0;
assign v$LEFT$SHIT_3063_out0 = v$LEFT$SHIFT_8801_out0;
assign v$LEFT$SHIT_3064_out0 = v$LEFT$SHIFT_8801_out0;
assign v$LEFT$SHIT_3065_out0 = v$LEFT$SHIFT_8801_out0;
assign v$LEFT$SHIT_3072_out0 = v$LEFT$SHIFT_8802_out0;
assign v$LEFT$SHIT_3073_out0 = v$LEFT$SHIFT_8802_out0;
assign v$LEFT$SHIT_3074_out0 = v$LEFT$SHIFT_8802_out0;
assign v$LEFT$SHIT_3075_out0 = v$LEFT$SHIFT_8802_out0;
assign v$LEFT$SHIT_3076_out0 = v$LEFT$SHIFT_8802_out0;
assign v$LEFT$SHIT_3089_out0 = v$LEFT$SHIFT_8803_out0;
assign v$LEFT$SHIT_3090_out0 = v$LEFT$SHIFT_8803_out0;
assign v$LEFT$SHIT_3091_out0 = v$LEFT$SHIFT_8803_out0;
assign v$LEFT$SHIT_3092_out0 = v$LEFT$SHIFT_8803_out0;
assign v$LEFT$SHIT_3093_out0 = v$LEFT$SHIFT_8803_out0;
assign v$LEFT$SHIT_3094_out0 = v$LEFT$SHIFT_8804_out0;
assign v$LEFT$SHIT_3095_out0 = v$LEFT$SHIFT_8804_out0;
assign v$LEFT$SHIT_3096_out0 = v$LEFT$SHIFT_8804_out0;
assign v$LEFT$SHIT_3097_out0 = v$LEFT$SHIFT_8804_out0;
assign v$LEFT$SHIT_3098_out0 = v$LEFT$SHIFT_8804_out0;
assign v$LEFT$SHIT_3099_out0 = v$LEFT$SHIFT_8805_out0;
assign v$LEFT$SHIT_3100_out0 = v$LEFT$SHIFT_8805_out0;
assign v$LEFT$SHIT_3101_out0 = v$LEFT$SHIFT_8805_out0;
assign v$LEFT$SHIT_3102_out0 = v$LEFT$SHIFT_8805_out0;
assign v$LEFT$SHIT_3103_out0 = v$LEFT$SHIFT_8805_out0;
assign v$_3109_out0 = v$_11816_out1[0:0];
assign v$_3109_out1 = v$_11816_out1[1:1];
assign v$_3110_out0 = v$_11817_out1[0:0];
assign v$_3110_out1 = v$_11817_out1[1:1];
assign v$_3685_out0 = v$_10810_out1[0:0];
assign v$_3685_out1 = v$_10810_out1[1:1];
assign v$_3686_out0 = v$_10811_out1[0:0];
assign v$_3686_out1 = v$_10811_out1[1:1];
assign v$XOR1_3954_out0 = v$A1_2938_out0 ^ v$C3_7014_out0;
assign v$SEL13_4841_out0 = v$IR2_1750_out0[9:8];
assign v$SEL13_4842_out0 = v$IR2_1751_out0[9:8];
assign v$CARRY_5003_out0 = v$CARRY_10908_out0;
assign v$CARRY_5004_out0 = v$CARRY_10909_out0;
assign v$_5074_out0 = v$_11816_out0[0:0];
assign v$_5074_out1 = v$_11816_out0[1:1];
assign v$_5075_out0 = v$_11817_out0[0:0];
assign v$_5075_out1 = v$_11817_out0[1:1];
assign v$_6461_out0 = v$_1528_out1[3:0];
assign v$_6461_out1 = v$_1528_out1[7:4];
assign v$_6462_out0 = v$_1529_out1[3:0];
assign v$_6462_out1 = v$_1529_out1[7:4];
assign v$_6982_out0 = v$_10810_out0[0:0];
assign v$_6982_out1 = v$_10810_out0[1:1];
assign v$_6983_out0 = v$_10811_out0[0:0];
assign v$_6983_out1 = v$_10811_out0[1:1];
assign v$EDGE2_7000_out0 = v$INTERRUPT2_3854_out0;
assign v$SEL4_7053_out0 = v$IR2_1750_out0[15:15];
assign v$SEL4_7054_out0 = v$IR2_1751_out0[15:15];
assign v$CLK4_7060_out0 = v$CLK4_16733_out0;
assign v$CLK4_7061_out0 = v$CLK4_16734_out0;
assign v$INSTR$READ_7221_out0 = v$INSTR$READ0_14172_out0;
assign v$INSTR$READ_7222_out0 = v$INSTR$READ1_11970_out0;
assign v$SEL10_7279_out0 = v$IR2_1750_out0[9:9];
assign v$SEL10_7280_out0 = v$IR2_1751_out0[9:9];
assign v$NQ0_7796_out0 = v$G4_13999_out0;
assign v$NQ0_7797_out0 = v$G4_14000_out0;
assign v$RAMDOUT1_8315_out0 = v$DM1_7858_out1;
assign v$SEL11_8352_out0 = v$IR2_1750_out0[8:8];
assign v$SEL11_8353_out0 = v$IR2_1751_out0[8:8];
assign v$_8408_out0 = v$_1528_out0[3:0];
assign v$_8408_out1 = v$_1528_out0[7:4];
assign v$_8409_out0 = v$_1529_out0[3:0];
assign v$_8409_out1 = v$_1529_out0[7:4];
assign v$G65_8809_out0 = ! v$PHALT_15137_out0;
assign v$_8935_out0 = { v$_18518_out0,v$_18326_out0 };
assign v$_8936_out0 = { v$_18519_out0,v$_18327_out0 };
assign v$RAMDOUT0_9099_out0 = v$DM1_7858_out0;
assign v$G3_9434_out0 = ! v$RXDISABLE_7888_out0;
assign v$G3_9435_out0 = ! v$RXDISABLE_7889_out0;
assign v$_9931_out0 = v$AROM1_16158_out0[27:0];
assign v$_9931_out1 = v$AROM1_16158_out0[43:16];
assign v$_9932_out0 = v$AROM1_16159_out0[27:0];
assign v$_9932_out1 = v$AROM1_16159_out0[43:16];
assign v$_10250_out0 = { v$_1829_out0,v$_13410_out0 };
assign v$_10251_out0 = { v$_1830_out0,v$_13411_out0 };
assign v$G25_10273_out0 = ! v$CALCULATING_7798_out0;
assign v$Mode_10976_out0 = v$MODE_9126_out0;
assign v$Mode_10977_out0 = v$MODE_9127_out0;
assign v$G3_10988_out0 = ! v$OFF_4039_out0;
assign v$G3_10989_out0 = ! v$OFF_4040_out0;
assign v$NQ1_11038_out0 = v$G2_15761_out0;
assign v$NQ1_11039_out0 = v$G2_15762_out0;
assign v$G8_12296_out0 = ((v$G6_13009_out0 && !v$G7_13431_out0) || (!v$G6_13009_out0) && v$G7_13431_out0);
assign v$G8_12297_out0 = ((v$G6_13010_out0 && !v$G7_13432_out0) || (!v$G6_13010_out0) && v$G7_13432_out0);
assign v$SEL12_12802_out0 = v$IR2_1750_out0[15:12];
assign v$SEL12_12803_out0 = v$IR2_1751_out0[15:12];
assign v$Mode_13197_out0 = v$MODE_9126_out0;
assign v$Mode_13198_out0 = v$MODE_9127_out0;
assign v$EQ1_13353_out0 = v$_8101_out0 == 3'h0;
assign v$EQ1_13354_out0 = v$_8102_out0 == 3'h0;
assign v$COUT_13515_out0 = v$A1_2938_out1;
assign v$G67_13755_out0 = ! v$PHALT_15137_out0;
assign v$G70_14028_out0 = v$PCHALT_16563_out0 && v$PHALT_15137_out0;
assign v$G67_14107_out0 = v$HALTED_11827_out0 && v$VALID$PREV_13429_out0;
assign v$G67_14108_out0 = v$HALTED_11828_out0 && v$VALID$PREV_13430_out0;
assign v$G4_14214_out0 = v$SOUT1_1919_out0 || v$INIT_10752_out0;
assign v$G4_14215_out0 = v$SOUT1_1925_out0 || v$INIT_10753_out0;
assign v$_14651_out0 = { v$_5474_out0,v$_7023_out0 };
assign v$_14652_out0 = { v$_5475_out0,v$_7024_out0 };
assign v$HALTSEL_14742_out0 = v$G2_7562_out0;
assign v$NQ0_15381_out0 = v$G9_16494_out0;
assign v$NQ0_15382_out0 = v$G9_16495_out0;
assign v$NQ0_15621_out0 = v$G1_1592_out0;
assign v$NQ0_15622_out0 = v$G1_1593_out0;
assign v$_15670_out0 = { v$_5517_out0,v$_16127_out0 };
assign v$_15671_out0 = { v$_5518_out0,v$_16128_out0 };
assign v$G69_15812_out0 = v$PCHALT_16563_out0 && v$PHALT_15137_out0;
assign v$G26_16019_out0 = ((v$G25_16104_out0 && !v$G22_7267_out0) || (!v$G25_16104_out0) && v$G22_7267_out0);
assign v$G26_16020_out0 = ((v$G25_16105_out0 && !v$G22_7268_out0) || (!v$G25_16105_out0) && v$G22_7268_out0);
assign v$CIN_16106_out0 = v$CIN_17342_out0;
assign v$CIN_16108_out0 = v$CIN_17344_out0;
assign v$CIN_16109_out0 = v$CIN_17345_out0;
assign v$NQ2_16698_out0 = v$G7_14311_out0;
assign v$NQ2_16699_out0 = v$G7_14312_out0;
assign v$NQ1_16729_out0 = v$G8_2267_out0;
assign v$NQ1_16730_out0 = v$G8_2268_out0;
assign v$CIN_16813_out0 = v$CIN_3887_out0;
assign v$PHALT_17485_out0 = v$G2_7562_out0;
assign v$CLEAR_18404_out0 = v$G1_33_out0;
assign v$CLEAR_18405_out0 = v$G1_34_out0;
assign v$RceivedParity_18539_out0 = v$RECIEVEDPARITY_6224_out0;
assign v$RceivedParity_18540_out0 = v$RECIEVEDPARITY_6225_out0;
assign v$NQ2_18563_out0 = v$G3_18414_out0;
assign v$NQ2_18564_out0 = v$G3_18415_out0;
assign v$PIPELINE$RESTART_18625_out0 = v$PIPELINE$RESTART_6071_out0;
assign v$PIPELINE$RESTART_18626_out0 = v$PIPELINE$RESTART_6072_out0;
assign v$_212_out0 = v$_8408_out1[1:0];
assign v$_212_out1 = v$_8408_out1[3:2];
assign v$_213_out0 = v$_8409_out1[1:0];
assign v$_213_out1 = v$_8409_out1[3:2];
assign v$G43_390_out0 = v$NQ2_18563_out0 && v$Q3_18425_out0;
assign v$G43_391_out0 = v$NQ2_18564_out0 && v$Q3_18426_out0;
assign v$G37_685_out0 = v$NQ0_7796_out0 || v$NQ1_254_out0;
assign v$G37_686_out0 = v$NQ0_7797_out0 || v$NQ1_255_out0;
assign v$S_1226_out0 = v$PHALT_17485_out0;
assign v$RXCLK_1240_out0 = v$EQ1_13353_out0;
assign v$RXCLK_1241_out0 = v$EQ1_13354_out0;
assign v$EQ12_1539_out0 = v$SEL12_12802_out0 == 4'h0;
assign v$EQ12_1540_out0 = v$SEL12_12803_out0 == 4'h0;
assign v$_1604_out0 = v$_6461_out1[1:0];
assign v$_1604_out1 = v$_6461_out1[3:2];
assign v$_1605_out0 = v$_6462_out1[1:0];
assign v$_1605_out1 = v$_6462_out1[3:2];
assign v$INTERRUPT2_1664_out0 = v$EDGE2_7000_out0;
assign v$_1671_out0 = v$_9931_out1[7:0];
assign v$_1671_out1 = v$_9931_out1[15:8];
assign v$_1672_out0 = v$_9932_out1[7:0];
assign v$_1672_out1 = v$_9932_out1[15:8];
assign v$G54_1901_out0 = v$NQ1_254_out0 && v$NQ0_7796_out0;
assign v$G54_1902_out0 = v$NQ1_255_out0 && v$NQ0_7797_out0;
assign v$G23_2277_out0 = v$NQ3_1491_out0 || v$NQ2_2980_out0;
assign v$G23_2278_out0 = v$NQ3_1492_out0 || v$NQ2_2981_out0;
assign v$_2289_out0 = v$_2345_out0[1:0];
assign v$_2289_out1 = v$_2345_out0[3:2];
assign v$_2290_out0 = v$_2346_out0[1:0];
assign v$_2290_out1 = v$_2346_out0[3:2];
assign v$G19_2412_out0 = v$NQ1_254_out0 && v$NQ2_2980_out0;
assign v$G19_2413_out0 = v$NQ1_255_out0 && v$NQ2_2981_out0;
assign v$G51_2863_out0 = v$Q3_18289_out0 && v$NQ2_2980_out0;
assign v$G51_2864_out0 = v$Q3_18290_out0 && v$NQ2_2981_out0;
assign v$G16_3022_out0 = v$NQ1_16729_out0 && v$Q2_3149_out0;
assign v$G16_3023_out0 = v$NQ1_16730_out0 && v$Q2_3150_out0;
assign v$G56_3143_out0 = v$NQ3_1491_out0 && v$Q0_13703_out0;
assign v$G56_3144_out0 = v$NQ3_1492_out0 && v$Q0_13704_out0;
assign v$Write_3255_out0 = v$CLEAR_18404_out0;
assign v$Write_3256_out0 = v$CLEAR_18404_out0;
assign v$Write_3257_out0 = v$CLEAR_18404_out0;
assign v$Write_3258_out0 = v$CLEAR_18404_out0;
assign v$Write_3259_out0 = v$CLEAR_18404_out0;
assign v$Write_3260_out0 = v$CLEAR_18404_out0;
assign v$Write_3261_out0 = v$CLEAR_18405_out0;
assign v$Write_3262_out0 = v$CLEAR_18405_out0;
assign v$Write_3263_out0 = v$CLEAR_18405_out0;
assign v$Write_3264_out0 = v$CLEAR_18405_out0;
assign v$Write_3265_out0 = v$CLEAR_18405_out0;
assign v$Write_3266_out0 = v$CLEAR_18405_out0;
assign v$F1_3488_out0 = v$_5074_out1;
assign v$F1_3489_out0 = v$_5075_out1;
assign v$C_3641_out0 = v$CARRY_5003_out0;
assign v$C_3642_out0 = v$CARRY_5004_out0;
assign v$CLK4_3694_out0 = v$CLK4_7060_out0;
assign v$CLK4_3695_out0 = v$CLK4_7061_out0;
assign v$RXENABLE_3716_out0 = v$G3_9434_out0;
assign v$RXENABLE_3717_out0 = v$G3_9435_out0;
assign v$G59_3843_out0 = v$Q2_17486_out0 && v$NQ3_2998_out0;
assign v$G59_3844_out0 = v$Q2_17487_out0 && v$NQ3_2999_out0;
assign v$R2_3845_out0 = v$_3685_out0;
assign v$R2_3846_out0 = v$_3686_out0;
assign v$IR2_3948_out0 = v$IR2_2217_out0;
assign v$IR2_3949_out0 = v$IR2_2218_out0;
assign v$G26_4097_out0 = v$G27_11706_out0 && v$NQ2_2980_out0;
assign v$G26_4098_out0 = v$G27_11707_out0 && v$NQ2_2981_out0;
assign v$G15_4205_out0 = v$NQ0_15621_out0 && v$Q1_4450_out0;
assign v$G15_4206_out0 = v$NQ0_15622_out0 && v$Q1_4451_out0;
assign v$G11_4865_out0 = v$NQ2_2980_out0 && v$NQ1_254_out0;
assign v$G11_4866_out0 = v$NQ2_2981_out0 && v$NQ1_255_out0;
assign v$_5142_out0 = v$_2345_out1[1:0];
assign v$_5142_out1 = v$_2345_out1[3:2];
assign v$_5143_out0 = v$_2346_out1[1:0];
assign v$_5143_out1 = v$_2346_out1[3:2];
assign v$EQ13_5251_out0 = v$SEL12_12802_out0 == 4'h1;
assign v$EQ13_5252_out0 = v$SEL12_12803_out0 == 4'h1;
assign v$_6075_out0 = v$Mode_10976_out0[0:0];
assign v$_6075_out1 = v$Mode_10976_out0[2:2];
assign v$_6076_out0 = v$Mode_10977_out0[0:0];
assign v$_6076_out1 = v$Mode_10977_out0[2:2];
assign v$Q_6153_out0 = v$_10250_out0;
assign v$Q_6154_out0 = v$_10251_out0;
assign v$IR2$REG$IMMEDIATE_6195_out0 = v$SEL10_7279_out0;
assign v$IR2$REG$IMMEDIATE_6196_out0 = v$SEL10_7280_out0;
assign v$G16_6407_out0 = v$NQ3_1491_out0 && v$Q2_5457_out0;
assign v$G16_6408_out0 = v$NQ3_1492_out0 && v$Q2_5458_out0;
assign v$_7374_out0 = v$_2897_out0[1:0];
assign v$_7374_out1 = v$_2897_out0[3:2];
assign v$_7375_out0 = v$_2898_out0[1:0];
assign v$_7375_out1 = v$_2898_out0[3:2];
assign v$G29_7465_out0 = v$NQ1_254_out0 || v$NQ0_7796_out0;
assign v$G29_7466_out0 = v$NQ1_255_out0 || v$NQ0_7797_out0;
assign v$IR2$FPU$OP_7546_out0 = v$SEL13_4841_out0;
assign v$IR2$FPU$OP_7547_out0 = v$SEL13_4842_out0;
assign v$_8208_out0 = v$_8408_out0[1:0];
assign v$_8208_out1 = v$_8408_out0[3:2];
assign v$_8209_out0 = v$_8409_out0[1:0];
assign v$_8209_out1 = v$_8409_out0[3:2];
assign v$G11_8230_out0 = v$NQ1_16729_out0 && v$NQ0_15381_out0;
assign v$G11_8231_out0 = v$NQ1_16730_out0 && v$NQ0_15382_out0;
assign v$F3_8247_out0 = v$_3109_out1;
assign v$F3_8248_out0 = v$_3110_out1;
assign v$CINA_8468_out0 = v$CIN_16106_out0;
assign v$CINA_8550_out0 = v$CIN_16108_out0;
assign v$CINA_8591_out0 = v$CIN_16109_out0;
assign v$G66_8931_out0 = v$PCHALT_16563_out0 && v$G65_8809_out0;
assign v$G32_9114_out0 = v$NQ1_11038_out0 || v$NQ0_15621_out0;
assign v$G32_9115_out0 = v$NQ1_11039_out0 || v$NQ0_15622_out0;
assign v$_9420_out0 = v$_2897_out1[1:0];
assign v$_9420_out1 = v$_2897_out1[3:2];
assign v$_9421_out0 = v$_2898_out1[1:0];
assign v$_9421_out1 = v$_2898_out1[3:2];
assign v$G42_9578_out0 = v$Q2_17486_out0 && v$NQ3_2998_out0;
assign v$G42_9579_out0 = v$Q2_17487_out0 && v$NQ3_2999_out0;
assign v$MUX1_9915_out0 = v$CLEAR_18404_out0 ? v$C3_13163_out0 : v$A1_4011_out0;
assign v$MUX1_9916_out0 = v$CLEAR_18405_out0 ? v$C3_13164_out0 : v$A1_4012_out0;
assign v$_9933_out0 = v$_1218_out1[2:0];
assign v$_9933_out1 = v$_1218_out1[5:3];
assign v$_9936_out0 = v$_1221_out1[2:0];
assign v$_9936_out1 = v$_1221_out1[5:3];
assign v$IS$IR2$DATA$PROCESSING_9944_out0 = v$SEL4_7053_out0;
assign v$IS$IR2$DATA$PROCESSING_9945_out0 = v$SEL4_7054_out0;
assign v$G49_10451_out0 = v$NQ3_1491_out0 && v$Q1_10923_out0;
assign v$G49_10452_out0 = v$NQ3_1492_out0 && v$Q1_10924_out0;
assign v$G5_10690_out0 = v$NQ2_16698_out0 && v$G6_3357_out0;
assign v$G5_10691_out0 = v$NQ2_16699_out0 && v$G6_3358_out0;
assign v$G36_10864_out0 = v$NQ2_2980_out0 && v$Q3_18289_out0;
assign v$G36_10865_out0 = v$NQ2_2981_out0 && v$Q3_18290_out0;
assign v$G17_11683_out0 = v$NQ2_2980_out0 && v$Q1_10923_out0;
assign v$G17_11684_out0 = v$NQ2_2981_out0 && v$Q1_10924_out0;
assign v$F2_12096_out0 = v$_3109_out0;
assign v$F2_12097_out0 = v$_3110_out0;
assign v$DATA$OUT0_12300_out0 = v$RAMDOUT0_9099_out0;
assign v$Q_12980_out0 = v$_8935_out0;
assign v$Q_12981_out0 = v$_8936_out0;
assign v$_12987_out0 = v$_1523_out1[2:0];
assign v$_12987_out1 = v$_1523_out1[5:3];
assign v$_12990_out0 = v$_1526_out1[2:0];
assign v$_12990_out1 = v$_1526_out1[5:3];
assign v$G50_13210_out0 = v$NQ3_1491_out0 && v$Q2_5457_out0;
assign v$G50_13211_out0 = v$NQ3_1492_out0 && v$Q2_5458_out0;
assign v$_13283_out0 = v$_6461_out0[1:0];
assign v$_13283_out1 = v$_6461_out0[3:2];
assign v$_13284_out0 = v$_6462_out0[1:0];
assign v$_13284_out1 = v$_6462_out0[3:2];
assign v$_13289_out0 = v$Mode_13197_out0[0:0];
assign v$_13289_out1 = v$Mode_13197_out0[2:2];
assign v$_13290_out0 = v$Mode_13198_out0[0:0];
assign v$_13290_out1 = v$Mode_13198_out0[2:2];
assign v$G9_13446_out0 = v$NQ2_18563_out0 && v$NQ1_11038_out0;
assign v$G9_13447_out0 = v$NQ2_18564_out0 && v$NQ1_11039_out0;
assign v$MUX6_13557_out0 = v$PIPELINE$RESTART_18625_out0 ? v$C2_13509_out0 : v$FF9_10664_out0;
assign v$MUX6_13558_out0 = v$PIPELINE$RESTART_18626_out0 ? v$C2_13510_out0 : v$FF9_10665_out0;
assign v$POut_13688_out0 = v$_15670_out0;
assign v$POut_13689_out0 = v$_15671_out0;
assign v$_13741_out0 = v$_1523_out0[2:0];
assign v$_13741_out1 = v$_1523_out0[5:3];
assign v$_13744_out0 = v$_1526_out0[2:0];
assign v$_13744_out1 = v$_1526_out0[5:3];
assign v$G68_14822_out0 = v$PCHALT_16563_out0 && v$G67_13755_out0;
assign v$INSTR$READ_14891_out0 = v$INSTR$READ_7221_out0;
assign v$INSTR$READ_14892_out0 = v$INSTR$READ_7222_out0;
assign v$G62_14987_out0 = v$Q3_18425_out0 && v$NQ2_18563_out0;
assign v$G62_14988_out0 = v$Q3_18426_out0 && v$NQ2_18564_out0;
assign v$R1_15011_out0 = v$_6982_out1;
assign v$R1_15012_out0 = v$_6983_out1;
assign v$R0_15192_out0 = v$_6982_out0;
assign v$R0_15193_out0 = v$_6983_out0;
assign v$R3_15314_out0 = v$_3685_out1;
assign v$R3_15315_out0 = v$_3686_out1;
assign v$DATA$OUT1_15602_out0 = v$RAMDOUT1_8315_out0;
assign v$F0_15834_out0 = v$_5074_out0;
assign v$F0_15835_out0 = v$_5075_out0;
assign v$G3_16089_out0 = ! v$PHALT_17485_out0;
assign v$IR2$RD_16358_out0 = v$SEL5_644_out0;
assign v$IR2$RD_16359_out0 = v$SEL5_645_out0;
assign v$_16367_out0 = v$_9931_out0[11:0];
assign v$_16367_out1 = v$_9931_out0[27:16];
assign v$_16368_out0 = v$_9932_out0[11:0];
assign v$_16368_out1 = v$_9932_out0[27:16];
assign v$G50_17323_out0 = v$Q2_17486_out0 && v$NQ3_2998_out0;
assign v$G50_17324_out0 = v$Q2_17487_out0 && v$NQ3_2999_out0;
assign v$EQ1_17399_out0 = v$XOR1_3954_out0 == 5'h0;
assign v$IR2$S$WB_17436_out0 = v$SEL11_8352_out0;
assign v$IR2$S$WB_17437_out0 = v$SEL11_8353_out0;
assign v$_17478_out0 = { v$G1_1195_out0,v$C2_18012_out0 };
assign v$_17479_out0 = { v$G1_1196_out0,v$C2_18013_out0 };
assign v$_17732_out0 = v$_1218_out0[2:0];
assign v$_17732_out1 = v$_1218_out0[5:3];
assign v$_17735_out0 = v$_1221_out0[2:0];
assign v$_17735_out1 = v$_1221_out0[5:3];
assign v$CLK4_17983_out0 = v$CLK4_7060_out0;
assign v$CLK4_17984_out0 = v$CLK4_7061_out0;
assign v$G68_18108_out0 = v$HALT$PREV$PREV_18074_out0 || v$G67_14107_out0;
assign v$G68_18109_out0 = v$HALT$PREV$PREV_18075_out0 || v$G67_14108_out0;
assign v$TX_18258_out0 = v$G4_14214_out0;
assign v$TX_18259_out0 = v$G4_14215_out0;
assign v$_18297_out0 = v$MODE_1617_out0[0:0];
assign v$_18297_out1 = v$MODE_1617_out0[2:2];
assign v$_18298_out0 = v$MODE_1618_out0[0:0];
assign v$_18298_out1 = v$MODE_1618_out0[2:2];
assign v$G14_18435_out0 = v$NQ0_15381_out0 && v$NQ2_16698_out0;
assign v$G14_18436_out0 = v$NQ0_15382_out0 && v$NQ2_16699_out0;
assign v$G42_18475_out0 = v$Q0_13703_out0 && v$NQ3_1491_out0;
assign v$G42_18476_out0 = v$Q0_13704_out0 && v$NQ3_1492_out0;
assign v$G60_18758_out0 = v$NQ3_2998_out0 && v$Q1_4450_out0;
assign v$G60_18759_out0 = v$NQ3_2999_out0 && v$Q1_4451_out0;
assign v$R_59_out0 = v$INSTR$READ_14891_out0;
assign v$R_60_out0 = v$INSTR$READ_14892_out0;
assign v$EQ7_231_out0 = v$Q_6153_out0 == 4'hc;
assign v$EQ7_232_out0 = v$Q_6154_out0 == 4'hc;
assign v$END_388_out0 = v$_13289_out1;
assign v$END_389_out0 = v$_13290_out1;
assign v$8_1193_out0 = v$IR2_3948_out0[11:10];
assign v$8_1194_out0 = v$IR2_3949_out0[11:10];
assign v$SEL12_1351_out0 = v$IR2_3948_out0[6:6];
assign v$SEL12_1352_out0 = v$IR2_3949_out0[6:6];
assign v$EQ6_1566_out0 = v$Q_6153_out0 == 4'hb;
assign v$EQ6_1567_out0 = v$Q_6154_out0 == 4'hb;
assign v$6_1948_out0 = v$IR2_3948_out0[15:15];
assign v$6_1949_out0 = v$IR2_3949_out0[15:15];
assign v$G48_2281_out0 = v$G51_2863_out0 && v$G54_1901_out0;
assign v$G48_2282_out0 = v$G51_2864_out0 && v$G54_1902_out0;
assign v$EQ3_2613_out0 = v$Q_6153_out0 == 4'hb;
assign v$EQ3_2614_out0 = v$Q_6154_out0 == 4'hb;
assign v$EQ4_2617_out0 = v$Q_12980_out0 == 4'h9;
assign v$EQ4_2618_out0 = v$Q_12981_out0 == 4'h9;
assign v$_2922_out0 = v$_13741_out0[0:0];
assign v$_2922_out1 = v$_13741_out0[2:2];
assign v$_2925_out0 = v$_13744_out0[0:0];
assign v$_2925_out1 = v$_13744_out0[2:2];
assign v$IR2_3286_out0 = v$IR2_3948_out0;
assign v$IR2_3287_out0 = v$IR2_3949_out0;
assign v$_3787_out0 = v$_7374_out0[0:0];
assign v$_3787_out1 = v$_7374_out0[1:1];
assign v$_3788_out0 = v$_7375_out0[0:0];
assign v$_3788_out1 = v$_7375_out0[1:1];
assign v$_3992_out0 = v$_6075_out1[0:0];
assign v$_3992_out1 = v$_6075_out1[1:1];
assign v$_3993_out0 = v$_6076_out1[0:0];
assign v$_3993_out1 = v$_6076_out1[1:1];
assign v$_4015_out0 = v$_8208_out0[0:0];
assign v$_4015_out1 = v$_8208_out0[1:1];
assign v$_4016_out0 = v$_8209_out0[0:0];
assign v$_4016_out1 = v$_8209_out0[1:1];
assign v$SEL10_4152_out0 = v$IR2_3948_out0[5:5];
assign v$SEL10_4153_out0 = v$IR2_3949_out0[5:5];
assign v$EQ3_4203_out0 = v$Q_12980_out0 == 4'hb;
assign v$EQ3_4204_out0 = v$Q_12981_out0 == 4'hb;
assign v$IR2$IS$LDST_4395_out0 = v$EQ12_1539_out0;
assign v$IR2$IS$LDST_4396_out0 = v$EQ12_1540_out0;
assign v$_4774_out0 = v$_212_out1[0:0];
assign v$_4774_out1 = v$_212_out1[1:1];
assign v$_4775_out0 = v$_213_out1[0:0];
assign v$_4775_out1 = v$_213_out1[1:1];
assign v$G47_5419_out0 = v$G49_10451_out0 || v$G50_13210_out0;
assign v$G47_5420_out0 = v$G49_10452_out0 || v$G50_13211_out0;
assign v$EQ14_5487_out0 = v$IR2$FPU$OP_7546_out0 == 2'h3;
assign v$EQ14_5488_out0 = v$IR2$FPU$OP_7547_out0 == 2'h3;
assign v$_5786_out0 = v$_212_out0[0:0];
assign v$_5786_out1 = v$_212_out0[1:1];
assign v$_5787_out0 = v$_213_out0[0:0];
assign v$_5787_out1 = v$_213_out0[1:1];
assign v$RX_6186_out0 = v$TX_18258_out0;
assign v$RX_6187_out0 = v$TX_18259_out0;
assign v$PIN_6636_out0 = v$_1671_out1;
assign v$PIN_6639_out0 = v$_1671_out0;
assign v$PIN_6642_out0 = v$_1672_out1;
assign v$PIN_6645_out0 = v$_1672_out0;
assign v$G21_7037_out0 = ! v$INTERRUPT2_1664_out0;
assign v$G58_7047_out0 = v$G60_18758_out0 || v$G59_3843_out0;
assign v$G58_7048_out0 = v$G60_18759_out0 || v$G59_3844_out0;
assign v$IR2$IS$FPU_7049_out0 = v$EQ13_5251_out0;
assign v$IR2$IS$FPU_7050_out0 = v$EQ13_5252_out0;
assign v$_7287_out0 = v$_13283_out1[0:0];
assign v$_7287_out1 = v$_13283_out1[1:1];
assign v$_7288_out0 = v$_13284_out1[0:0];
assign v$_7288_out1 = v$_13284_out1[1:1];
assign v$EQ1_7437_out0 = v$Q_6153_out0 == 4'h9;
assign v$EQ1_7438_out0 = v$Q_6154_out0 == 4'h9;
assign v$5_7508_out0 = v$IR2_3948_out0[1:0];
assign v$5_7509_out0 = v$IR2_3949_out0[1:0];
assign v$STP$SAVED_7560_out0 = v$MUX6_13557_out0;
assign v$STP$SAVED_7561_out0 = v$MUX6_13558_out0;
assign v$DATA$OUT_7608_out0 = v$DATA$OUT0_12300_out0;
assign v$DATA$OUT_7609_out0 = v$DATA$OUT1_15602_out0;
assign v$_7768_out0 = v$_17732_out0[0:0];
assign v$_7768_out1 = v$_17732_out0[2:2];
assign v$_7771_out0 = v$_17735_out0[0:0];
assign v$_7771_out1 = v$_17735_out0[2:2];
assign v$_7981_out0 = v$_2289_out1[0:0];
assign v$_7981_out1 = v$_2289_out1[1:1];
assign v$_7982_out0 = v$_2290_out1[0:0];
assign v$_7982_out1 = v$_2290_out1[1:1];
assign v$S_8021_out0 = v$S_1226_out0;
assign v$G61_8281_out0 = v$G62_14987_out0 && v$NQ1_11038_out0;
assign v$G61_8282_out0 = v$G62_14988_out0 && v$NQ1_11039_out0;
assign v$P_8310_out0 = v$_13289_out0;
assign v$P_8311_out0 = v$_13290_out0;
assign v$_8776_out0 = v$_1604_out0[0:0];
assign v$_8776_out1 = v$_1604_out0[1:1];
assign v$_8777_out0 = v$_1605_out0[0:0];
assign v$_8777_out1 = v$_1605_out0[1:1];
assign v$_8812_out0 = v$_5142_out1[0:0];
assign v$_8812_out1 = v$_5142_out1[1:1];
assign v$_8813_out0 = v$_5143_out1[0:0];
assign v$_8813_out1 = v$_5143_out1[1:1];
assign v$_9062_out0 = v$_9933_out1[0:0];
assign v$_9062_out1 = v$_9933_out1[2:2];
assign v$_9065_out0 = v$_9936_out1[0:0];
assign v$_9065_out1 = v$_9936_out1[2:2];
assign v$EQ5_9106_out0 = v$Q_6153_out0 == 4'ha;
assign v$EQ5_9107_out0 = v$Q_6154_out0 == 4'ha;
assign v$SEL4_9443_out0 = v$IR2_3948_out0[9:8];
assign v$SEL4_9444_out0 = v$IR2_3949_out0[9:8];
assign v$G60_9467_out0 = v$G61_16446_out0 && v$G68_18108_out0;
assign v$G60_9468_out0 = v$G61_16447_out0 && v$G68_18109_out0;
assign v$_9482_out0 = v$_9420_out0[0:0];
assign v$_9482_out1 = v$_9420_out0[1:1];
assign v$_9483_out0 = v$_9421_out0[0:0];
assign v$_9483_out1 = v$_9421_out0[1:1];
assign v$EQ4_9625_out0 = v$Q_6153_out0 == 4'hc;
assign v$EQ4_9626_out0 = v$Q_6154_out0 == 4'hc;
assign v$RXBYTE_9628_out0 = v$POut_13688_out0;
assign v$RXBYTE_9629_out0 = v$POut_13689_out0;
assign v$_10772_out0 = v$_12987_out1[0:0];
assign v$_10772_out1 = v$_12987_out1[2:2];
assign v$_10775_out0 = v$_12990_out1[0:0];
assign v$_10775_out1 = v$_12990_out1[2:2];
assign v$EQ2_11605_out0 = v$Q_12980_out0 == 4'ha;
assign v$EQ2_11606_out0 = v$Q_12981_out0 == 4'ha;
assign v$G28_11939_out0 = v$Q2_5457_out0 && v$G29_7465_out0;
assign v$G28_11940_out0 = v$Q2_5458_out0 && v$G29_7466_out0;
assign v$PARITY_12073_out0 = v$_18297_out0;
assign v$PARITY_12074_out0 = v$_18298_out0;
assign v$_12077_out0 = v$_8208_out1[0:0];
assign v$_12077_out1 = v$_8208_out1[1:1];
assign v$_12078_out0 = v$_8209_out1[0:0];
assign v$_12078_out1 = v$_8209_out1[1:1];
assign v$G35_12635_out0 = v$G36_10864_out0 && v$G37_685_out0;
assign v$G35_12636_out0 = v$G36_10865_out0 && v$G37_686_out0;
assign v$_12902_out0 = v$_16367_out0[3:0];
assign v$_12902_out1 = v$_16367_out0[11:8];
assign v$_12903_out0 = v$_16368_out0[3:0];
assign v$_12903_out1 = v$_16368_out0[11:8];
assign v$G40_13678_out0 = v$G41_18479_out0 && v$G42_9578_out0;
assign v$G40_13679_out0 = v$G41_18480_out0 && v$G42_9579_out0;
assign {v$A1_13701_out1,v$A1_13701_out0 } = v$REG1_13592_out0 + v$_17478_out0 + v$C1_6457_out0;
assign {v$A1_13702_out1,v$A1_13702_out0 } = v$REG1_13593_out0 + v$_17479_out0 + v$C1_6458_out0;
assign v$_13842_out0 = v$_7374_out1[0:0];
assign v$_13842_out1 = v$_7374_out1[1:1];
assign v$_13843_out0 = v$_7375_out1[0:0];
assign v$_13843_out1 = v$_7375_out1[1:1];
assign v$9_14162_out0 = v$IR2_3948_out0[14:12];
assign v$9_14163_out0 = v$IR2_3949_out0[14:12];
assign v$_14247_out0 = v$_1604_out1[0:0];
assign v$_14247_out1 = v$_1604_out1[1:1];
assign v$_14248_out0 = v$_1605_out1[0:0];
assign v$_14248_out1 = v$_1605_out1[1:1];
assign v$EQ1_14322_out0 = v$Q_12980_out0 == 4'h1;
assign v$EQ1_14323_out0 = v$Q_12981_out0 == 4'h1;
assign v$_14509_out0 = v$_2289_out0[0:0];
assign v$_14509_out1 = v$_2289_out0[1:1];
assign v$_14510_out0 = v$_2290_out0[0:0];
assign v$_14510_out1 = v$_2290_out0[1:1];
assign v$G25_14579_out0 = v$INTERRUPT2_1664_out0 && v$G24_12088_out0;
assign v$G2_15033_out0 = ! v$Write_3255_out0;
assign v$G2_15034_out0 = ! v$Write_3256_out0;
assign v$G2_15035_out0 = ! v$Write_3257_out0;
assign v$G2_15036_out0 = ! v$Write_3258_out0;
assign v$G2_15037_out0 = ! v$Write_3259_out0;
assign v$G2_15038_out0 = ! v$Write_3260_out0;
assign v$G2_15039_out0 = ! v$Write_3261_out0;
assign v$G2_15040_out0 = ! v$Write_3262_out0;
assign v$G2_15041_out0 = ! v$Write_3263_out0;
assign v$G2_15042_out0 = ! v$Write_3264_out0;
assign v$G2_15043_out0 = ! v$Write_3265_out0;
assign v$G2_15044_out0 = ! v$Write_3266_out0;
assign v$_15148_out0 = v$_9933_out0[0:0];
assign v$_15148_out1 = v$_9933_out0[2:2];
assign v$_15151_out0 = v$_9936_out0[0:0];
assign v$_15151_out1 = v$_9936_out0[2:2];
assign v$_15186_out0 = v$_13283_out0[0:0];
assign v$_15186_out1 = v$_13283_out0[1:1];
assign v$_15187_out0 = v$_13284_out0[0:0];
assign v$_15187_out1 = v$_13284_out0[1:1];
assign v$7_15358_out0 = v$IR2_3948_out0[8:8];
assign v$7_15359_out0 = v$IR2_3949_out0[8:8];
assign v$ParityEN_15784_out0 = v$_6075_out0;
assign v$ParityEN_15785_out0 = v$_6076_out0;
assign v$_15839_out0 = v$_9420_out1[0:0];
assign v$_15839_out1 = v$_9420_out1[1:1];
assign v$_15840_out0 = v$_9421_out1[0:0];
assign v$_15840_out1 = v$_9421_out1[1:1];
assign v$RXCLK_15844_out0 = v$RXCLK_1240_out0;
assign v$RXCLK_15845_out0 = v$RXCLK_1241_out0;
assign v$SEL11_15890_out0 = v$IR2_3948_out0[7:7];
assign v$SEL11_15891_out0 = v$IR2_3949_out0[7:7];
assign v$C_15895_out0 = v$C_3641_out0;
assign v$C_15896_out0 = v$C_3642_out0;
assign v$_16265_out0 = v$_17732_out1[0:0];
assign v$_16265_out1 = v$_17732_out1[2:2];
assign v$_16268_out0 = v$_17735_out1[0:0];
assign v$_16268_out1 = v$_17735_out1[2:2];
assign v$_16740_out0 = v$_13741_out1[0:0];
assign v$_16740_out1 = v$_13741_out1[2:2];
assign v$_16743_out0 = v$_13744_out1[0:0];
assign v$_16743_out1 = v$_13744_out1[2:2];
assign v$R_16745_out0 = v$G3_16089_out0;
assign v$_16760_out0 = v$_16367_out1[7:0];
assign v$_16760_out1 = v$_16367_out1[15:8];
assign v$_16761_out0 = v$_16368_out1[7:0];
assign v$_16761_out1 = v$_16368_out1[15:8];
assign v$G39_16890_out0 = v$Q2_5457_out0 && v$G42_18475_out0;
assign v$G39_16891_out0 = v$Q2_5458_out0 && v$G42_18476_out0;
assign v$_16980_out0 = v$_5142_out0[0:0];
assign v$_16980_out1 = v$_5142_out0[1:1];
assign v$_16981_out0 = v$_5143_out0[0:0];
assign v$_16981_out1 = v$_5143_out0[1:1];
assign v$G21_17674_out0 = v$G23_2277_out0 && v$G22_4313_out0;
assign v$G21_17675_out0 = v$G23_2278_out0 && v$G22_4314_out0;
assign v$_17981_out0 = v$_18297_out1[0:0];
assign v$_17981_out1 = v$_18297_out1[1:1];
assign v$_17982_out0 = v$_18298_out1[0:0];
assign v$_17982_out1 = v$_18298_out1[1:1];
assign v$_18188_out0 = v$_12987_out0[0:0];
assign v$_18188_out1 = v$_12987_out0[2:2];
assign v$_18191_out0 = v$_12990_out0[0:0];
assign v$_18191_out1 = v$_12990_out0[2:2];
assign v$MUX1_18598_out0 = v$EQ1_17399_out0 ? v$C4_14657_out0 : v$A1_2938_out0;
assign v$G31_18635_out0 = v$G32_9114_out0 && v$NQ3_2998_out0;
assign v$G31_18636_out0 = v$G32_9115_out0 && v$NQ3_2999_out0;
assign v$EQ2_18657_out0 = v$Q_6153_out0 == 4'h0;
assign v$EQ2_18658_out0 = v$Q_6154_out0 == 4'h0;
assign v$G56_648_out0 = v$EQ3_2613_out0 || v$EQ4_9625_out0;
assign v$G56_649_out0 = v$EQ3_2614_out0 || v$EQ4_9626_out0;
assign v$IR2$S_1169_out0 = v$7_15358_out0;
assign v$IR2$S_1170_out0 = v$7_15359_out0;
assign v$G9_1184_out0 = ((v$_7287_out1 && !v$_13842_out1) || (!v$_7287_out1) && v$_13842_out1);
assign v$G9_1185_out0 = ((v$_7288_out1 && !v$_13843_out1) || (!v$_7288_out1) && v$_13843_out1);
assign v$DATA$OUT_1307_out0 = v$DATA$OUT_7608_out0;
assign v$DATA$OUT_1308_out0 = v$DATA$OUT_7609_out0;
assign v$G4_1329_out0 = ((v$_12077_out1 && !v$_7981_out1) || (!v$_12077_out1) && v$_7981_out1);
assign v$G4_1330_out0 = ((v$_12078_out1 && !v$_7982_out1) || (!v$_12078_out1) && v$_7982_out1);
assign v$G47_1531_out0 = v$PARITY_12073_out0 && v$EQ1_7437_out0;
assign v$G47_1532_out0 = v$PARITY_12074_out0 && v$EQ1_7438_out0;
assign v$R_1590_out0 = v$R_16745_out0;
assign v$_1669_out0 = { v$C8_7281_out0,v$_12902_out0 };
assign v$_1670_out0 = { v$C8_7282_out0,v$_12903_out0 };
assign v$IR2$FPU$OP_1687_out0 = v$SEL4_9443_out0;
assign v$IR2$FPU$OP_1688_out0 = v$SEL4_9444_out0;
assign v$G12_1820_out0 = ((v$_8776_out1 && !v$_9482_out1) || (!v$_8776_out1) && v$_9482_out1);
assign v$G12_1821_out0 = ((v$_8777_out1 && !v$_9483_out1) || (!v$_8777_out1) && v$_9483_out1);
assign v$G15_1868_out0 = ((v$_8776_out0 && !v$_9482_out0) || (!v$_8776_out0) && v$_9482_out0);
assign v$G15_1869_out0 = ((v$_8777_out0 && !v$_9483_out0) || (!v$_8777_out0) && v$_9483_out0);
assign v$B12_1950_out0 = v$_7768_out0;
assign v$B12_1953_out0 = v$_7771_out0;
assign v$G10_1998_out0 = ((v$_14247_out1 && !v$_15839_out1) || (!v$_14247_out1) && v$_15839_out1);
assign v$G10_1999_out0 = ((v$_14248_out1 && !v$_15840_out1) || (!v$_14248_out1) && v$_15840_out1);
assign v$G25_2464_out0 = v$IR2$IS$LDST_4395_out0 && v$IR2$S$WB_17436_out0;
assign v$G25_2465_out0 = v$IR2$IS$LDST_4396_out0 && v$IR2$S$WB_17437_out0;
assign v$G30_2466_out0 = v$G31_18635_out0 && v$Q2_17486_out0;
assign v$G30_2467_out0 = v$G31_18636_out0 && v$Q2_17487_out0;
assign v$B0_3200_out0 = v$_2922_out0;
assign v$B0_3203_out0 = v$_2925_out0;
assign v$2StopBits_3484_out0 = v$_3992_out1;
assign v$2StopBits_3485_out0 = v$_3993_out1;
assign v$G16_3520_out0 = ((v$_7287_out0 && !v$_13842_out0) || (!v$_7287_out0) && v$_13842_out0);
assign v$G16_3521_out0 = ((v$_7288_out0 && !v$_13843_out0) || (!v$_7288_out0) && v$_13843_out0);
assign v$S_4025_out0 = v$_17981_out1;
assign v$S_4026_out0 = v$_17982_out1;
assign v$B9_4065_out0 = v$_10772_out0;
assign v$B9_4068_out0 = v$_10775_out0;
assign v$IR2$FPU$LOAD_4231_out0 = v$SEL11_15890_out0;
assign v$IR2$FPU$LOAD_4232_out0 = v$SEL11_15891_out0;
assign v$G8_4819_out0 = ((v$_4774_out1 && !v$_8812_out1) || (!v$_4774_out1) && v$_8812_out1);
assign v$G8_4820_out0 = ((v$_4775_out1 && !v$_8813_out1) || (!v$_4775_out1) && v$_8813_out1);
assign v$_4997_out0 = v$IR2_3286_out0[14:12];
assign v$_4998_out0 = v$IR2_3287_out0[14:12];
assign v$OUT_5002_out0 = v$MUX1_18598_out0;
assign v$G55_5049_out0 = v$G56_3143_out0 || v$G48_2281_out0;
assign v$G55_5050_out0 = v$G56_3144_out0 || v$G48_2282_out0;
assign v$G2_5429_out0 = ((v$_4015_out1 && !v$_14509_out1) || (!v$_4015_out1) && v$_14509_out1);
assign v$G2_5430_out0 = ((v$_4016_out1 && !v$_14510_out1) || (!v$_4016_out1) && v$_14510_out1);
assign v$G22_5463_out0 = v$G25_14579_out0 && v$R2_3846_out0;
assign v$G39_6045_out0 = v$G40_13678_out0 || v$G43_390_out0;
assign v$G39_6046_out0 = v$G40_13679_out0 || v$G43_391_out0;
assign v$G6_6163_out0 = ((v$_5786_out1 && !v$_16980_out1) || (!v$_5786_out1) && v$_16980_out1);
assign v$G6_6164_out0 = ((v$_5787_out1 && !v$_16981_out1) || (!v$_5787_out1) && v$_16981_out1);
assign v$PIN_6634_out0 = v$_16760_out1;
assign v$PIN_6635_out0 = v$_16760_out0;
assign v$PIN_6638_out0 = v$_12902_out1;
assign v$PIN_6640_out0 = v$_16761_out1;
assign v$PIN_6641_out0 = v$_16761_out0;
assign v$PIN_6644_out0 = v$_12903_out1;
assign v$_6898_out0 = v$_18188_out1[0:0];
assign v$_6898_out1 = v$_18188_out1[1:1];
assign v$_6901_out0 = v$_18191_out1[0:0];
assign v$_6901_out1 = v$_18191_out1[1:1];
assign v$_6977_out0 = v$_16740_out1[0:0];
assign v$_6977_out1 = v$_16740_out1[1:1];
assign v$_6980_out0 = v$_16743_out1[0:0];
assign v$_6980_out1 = v$_16743_out1[1:1];
assign v$_6990_out0 = v$IR2_3286_out0[7:4];
assign v$_6991_out0 = v$IR2_3287_out0[7:4];
assign v$_7273_out0 = v$IR2_3286_out0[4:0];
assign v$_7274_out0 = v$IR2_3287_out0[4:0];
assign v$IR2$15_7435_out0 = v$6_1948_out0;
assign v$IR2$15_7436_out0 = v$6_1949_out0;
assign v$IR2_7773_out0 = v$IR2_3286_out0;
assign v$IR2_7774_out0 = v$IR2_3287_out0;
assign v$G64_7783_out0 = v$EQ3_4203_out0 && v$G63_10019_out0;
assign v$G64_7784_out0 = v$EQ3_4204_out0 && v$G63_10020_out0;
assign v$G11_8263_out0 = ((v$_15186_out1 && !v$_3787_out1) || (!v$_15186_out1) && v$_3787_out1);
assign v$G11_8264_out0 = ((v$_15187_out1 && !v$_3788_out1) || (!v$_15187_out1) && v$_3788_out1);
assign v$CLK4_8834_out0 = v$RXCLK_15844_out0;
assign v$CLK4_8835_out0 = v$RXCLK_15845_out0;
assign v$RXBIT_8913_out0 = v$RX_6186_out0;
assign v$RXBIT_8914_out0 = v$RX_6187_out0;
assign v$G57_8978_out0 = v$EQ2_11605_out0 && v$G58_168_out0;
assign v$G57_8979_out0 = v$EQ2_11606_out0 && v$G58_169_out0;
assign v$_9381_out0 = v$_9062_out1[0:0];
assign v$_9381_out1 = v$_9062_out1[1:1];
assign v$_9384_out0 = v$_9065_out1[0:0];
assign v$_9384_out1 = v$_9065_out1[1:1];
assign v$B3_9471_out0 = v$_16740_out0;
assign v$B3_9474_out0 = v$_16743_out0;
assign v$_9497_out0 = v$_10772_out1[0:0];
assign v$_9497_out1 = v$_10772_out1[1:1];
assign v$_9500_out0 = v$_10775_out1[0:0];
assign v$_9500_out1 = v$_10775_out1[1:1];
assign v$G23_9602_out0 = v$FF3_15031_out0 && v$G21_7037_out0;
assign v$B15_10021_out0 = v$_16265_out0;
assign v$B15_10024_out0 = v$_16268_out0;
assign v$G1_10317_out0 = ((v$_4015_out0 && !v$_14509_out0) || (!v$_4015_out0) && v$_14509_out0);
assign v$G1_10318_out0 = ((v$_4016_out0 && !v$_14510_out0) || (!v$_4016_out0) && v$_14510_out0);
assign v$OddParity_10686_out0 = v$_3992_out0;
assign v$OddParity_10687_out0 = v$_3993_out0;
assign v$B18_10867_out0 = v$_15148_out0;
assign v$B18_10870_out0 = v$_15151_out0;
assign v$Q1P_11007_out0 = v$G21_17674_out0;
assign v$Q1P_11008_out0 = v$G21_17675_out0;
assign v$_11022_out0 = v$_2922_out1[0:0];
assign v$_11022_out1 = v$_2922_out1[1:1];
assign v$_11025_out0 = v$_2925_out1[0:0];
assign v$_11025_out1 = v$_2925_out1[1:1];
assign v$_11391_out0 = v$IR2_3286_out0[9:9];
assign v$_11392_out0 = v$IR2_3287_out0[9:9];
assign v$G61_11603_out0 = v$EQ4_2617_out0 && v$P_8310_out0;
assign v$G61_11604_out0 = v$EQ4_2618_out0 && v$P_8311_out0;
assign v$IR2$FPU$32BIT_11800_out0 = v$SEL10_4152_out0;
assign v$IR2$FPU$32BIT_11801_out0 = v$SEL10_4153_out0;
assign v$G14_12046_out0 = ((v$_14247_out0 && !v$_15839_out0) || (!v$_14247_out0) && v$_15839_out0);
assign v$G14_12047_out0 = ((v$_14248_out0 && !v$_15840_out0) || (!v$_14248_out0) && v$_15840_out0);
assign v$G7_12647_out0 = ((v$_4774_out0 && !v$_8812_out0) || (!v$_4774_out0) && v$_8812_out0);
assign v$G7_12648_out0 = ((v$_4775_out0 && !v$_8813_out0) || (!v$_4775_out0) && v$_8813_out0);
assign v$G53_12714_out0 = v$EQ1_14322_out0 && v$G52_15938_out0;
assign v$G53_12715_out0 = v$EQ1_14323_out0 && v$G52_15939_out0;
assign v$_12862_out0 = v$PIN_6636_out0[3:0];
assign v$_12862_out1 = v$PIN_6636_out0[7:4];
assign v$_12865_out0 = v$PIN_6639_out0[3:0];
assign v$_12865_out1 = v$PIN_6639_out0[7:4];
assign v$_12868_out0 = v$PIN_6642_out0[3:0];
assign v$_12868_out1 = v$PIN_6642_out0[7:4];
assign v$_12871_out0 = v$PIN_6645_out0[3:0];
assign v$_12871_out1 = v$PIN_6645_out0[7:4];
assign v$IR2$M_12993_out0 = v$5_7508_out0;
assign v$IR2$M_12994_out0 = v$5_7509_out0;
assign v$_13180_out0 = v$_16265_out1[0:0];
assign v$_13180_out1 = v$_16265_out1[1:1];
assign v$_13183_out0 = v$_16268_out1[0:0];
assign v$_13183_out1 = v$_16268_out1[1:1];
assign v$B6_13298_out0 = v$_18188_out0;
assign v$B6_13301_out0 = v$_18191_out0;
assign v$G13_13444_out0 = ((v$_15186_out0 && !v$_3787_out0) || (!v$_15186_out0) && v$_3787_out0);
assign v$G13_13445_out0 = ((v$_15187_out0 && !v$_3788_out0) || (!v$_15187_out0) && v$_3788_out0);
assign v$G57_13452_out0 = v$G61_8281_out0 || v$G58_7047_out0;
assign v$G57_13453_out0 = v$G61_8282_out0 || v$G58_7048_out0;
assign v$G18_13513_out0 = ! v$C_15895_out0;
assign v$G18_13514_out0 = ! v$C_15896_out0;
assign v$IR2$D_14491_out0 = v$8_1193_out0;
assign v$IR2$D_14492_out0 = v$8_1194_out0;
assign v$G28_14668_out0 = v$IR2$IS$FPU_7049_out0 && v$EQ14_5487_out0;
assign v$G28_14669_out0 = v$IR2$IS$FPU_7050_out0 && v$EQ14_5488_out0;
assign v$G59_15123_out0 = v$G58_2518_out0 || v$G60_9467_out0;
assign v$G59_15124_out0 = v$G58_2519_out0 || v$G60_9468_out0;
assign v$G40_15130_out0 = v$Q1_10923_out0 && v$G39_16890_out0;
assign v$G40_15131_out0 = v$Q1_10924_out0 && v$G39_16891_out0;
assign v$G5_15232_out0 = ((v$_5786_out0 && !v$_16980_out0) || (!v$_5786_out0) && v$_16980_out0);
assign v$G5_15233_out0 = ((v$_5787_out0 && !v$_16981_out0) || (!v$_5787_out0) && v$_16981_out0);
assign v$IR2$FPU$LOADA_15268_out0 = v$SEL12_1351_out0;
assign v$IR2$FPU$LOADA_15269_out0 = v$SEL12_1352_out0;
assign v$G22_15342_out0 = ! v$C_15895_out0;
assign v$G22_15343_out0 = ! v$C_15896_out0;
assign v$G28_15633_out0 = v$STALL$PREV$CYCLE_5772_out0 || v$STP$SAVED_7560_out0;
assign v$G28_15634_out0 = v$STALL$PREV$CYCLE_5773_out0 || v$STP$SAVED_7561_out0;
assign v$END_15738_out0 = v$A1_13701_out1;
assign v$END_15739_out0 = v$A1_13702_out1;
assign v$ODDPARITY_15928_out0 = v$_17981_out0;
assign v$ODDPARITY_15929_out0 = v$_17982_out0;
assign v$_16589_out0 = v$_15148_out1[0:0];
assign v$_16589_out1 = v$_15148_out1[1:1];
assign v$_16592_out0 = v$_15151_out1[0:0];
assign v$_16592_out1 = v$_15151_out1[1:1];
assign v$SEL3_16650_out0 = v$IR2_3286_out0[15:12];
assign v$SEL3_16651_out0 = v$IR2_3287_out0[15:12];
assign v$_16737_out0 = v$IR2_3286_out0[3:2];
assign v$_16738_out0 = v$IR2_3287_out0[3:2];
assign v$G45_16900_out0 = ! v$P_8310_out0;
assign v$G45_16901_out0 = ! v$P_8311_out0;
assign v$_17325_out0 = v$_7768_out1[0:0];
assign v$_17325_out1 = v$_7768_out1[1:1];
assign v$_17328_out0 = v$_7771_out1[0:0];
assign v$_17328_out1 = v$_7771_out1[1:1];
assign v$G3_17452_out0 = ((v$_12077_out0 && !v$_7981_out0) || (!v$_12077_out0) && v$_7981_out0);
assign v$G3_17453_out0 = ((v$_12078_out0 && !v$_7982_out0) || (!v$_12078_out0) && v$_7982_out0);
assign v$_18018_out0 = v$IR2_3286_out0[8:8];
assign v$_18019_out0 = v$IR2_3287_out0[8:8];
assign v$IR2$OP_18020_out0 = v$9_14162_out0;
assign v$IR2$OP_18021_out0 = v$9_14163_out0;
assign v$B21_18082_out0 = v$_9062_out0;
assign v$B21_18085_out0 = v$_9065_out0;
assign v$G25_18095_out0 = v$G26_4097_out0 || v$G28_11939_out0;
assign v$G25_18096_out0 = v$G26_4098_out0 || v$G28_11940_out0;
assign v$R_18353_out0 = v$R_59_out0;
assign v$R_18354_out0 = v$R_60_out0;
assign v$G35_18495_out0 = ! v$IR2$IS$LDST_4395_out0;
assign v$G35_18496_out0 = ! v$IR2$IS$LDST_4396_out0;
assign v$G33_18616_out0 = v$IR2$IS$LDST_4395_out0 && v$IR2$S$WB_17436_out0;
assign v$G33_18617_out0 = v$IR2$IS$LDST_4396_out0 && v$IR2$S$WB_17437_out0;
assign v$EQ7_18631_out0 = v$IR2_3286_out0 == 16'h7000;
assign v$EQ7_18632_out0 = v$IR2_3287_out0 == 16'h7000;
assign v$G2_18697_out0 = v$RXENABLE_3716_out0 && v$RXCLK_15844_out0;
assign v$G2_18698_out0 = v$RXENABLE_3717_out0 && v$RXCLK_15845_out0;
assign v$RX_43_out0 = v$RXBIT_8913_out0;
assign v$RX_44_out0 = v$RXBIT_8914_out0;
assign v$G27_260_out0 = v$G1_10317_out0 || v$G2_5429_out0;
assign v$G27_261_out0 = v$G1_10318_out0 || v$G2_5430_out0;
assign v$K_301_out0 = v$_7273_out0;
assign v$K_302_out0 = v$_7274_out0;
assign v$G17_362_out0 = v$S_4025_out0 && v$NQ2_18563_out0;
assign v$G17_363_out0 = v$S_4026_out0 && v$NQ2_18564_out0;
assign v$B23_1283_out0 = v$_9381_out1;
assign v$B23_1286_out0 = v$_9384_out1;
assign v$G25_1309_out0 = v$G5_15232_out0 || v$G6_6163_out0;
assign v$G25_1310_out0 = v$G5_15233_out0 || v$G6_6164_out0;
assign v$OP_1872_out0 = v$IR2$OP_18020_out0;
assign v$OP_1873_out0 = v$IR2$OP_18021_out0;
assign v$B_2696_out0 = v$B6_13298_out0;
assign v$B_2697_out0 = v$B3_9471_out0;
assign v$B_2698_out0 = v$B21_18082_out0;
assign v$B_2699_out0 = v$B9_4065_out0;
assign v$B_2700_out0 = v$B15_10021_out0;
assign v$B_2704_out0 = v$B12_1950_out0;
assign v$B_2708_out0 = v$B0_3200_out0;
assign v$B_2713_out0 = v$B18_10867_out0;
assign v$B_2768_out0 = v$B6_13301_out0;
assign v$B_2769_out0 = v$B3_9474_out0;
assign v$B_2770_out0 = v$B21_18085_out0;
assign v$B_2771_out0 = v$B9_4068_out0;
assign v$B_2772_out0 = v$B15_10024_out0;
assign v$B_2776_out0 = v$B12_1953_out0;
assign v$B_2780_out0 = v$B0_3203_out0;
assign v$B_2785_out0 = v$B18_10870_out0;
assign v$RX_2966_out0 = v$RXBIT_8913_out0;
assign v$RX_2967_out0 = v$RXBIT_8914_out0;
assign v$G52_2971_out0 = v$S_4025_out0 || v$NQ0_15621_out0;
assign v$G52_2972_out0 = v$S_4026_out0 || v$NQ0_15622_out0;
assign v$B2_3113_out0 = v$_11022_out1;
assign v$B2_3116_out0 = v$_11025_out1;
assign v$C_3198_out0 = v$_11391_out0;
assign v$C_3199_out0 = v$_11392_out0;
assign v$G12_3615_out0 = ! v$IR2$FPU$LOADA_15268_out0;
assign v$G12_3616_out0 = ! v$IR2$FPU$LOADA_15269_out0;
assign v$B20_3943_out0 = v$_16589_out1;
assign v$B20_3946_out0 = v$_16592_out1;
assign v$B14_4002_out0 = v$_17325_out1;
assign v$B14_4005_out0 = v$_17328_out1;
assign v$IR1_4156_out0 = v$R_18353_out0;
assign v$IR1_4157_out0 = v$R_18354_out0;
assign v$IR2$VALID_4217_out0 = v$G59_15123_out0;
assign v$IR2$VALID_4218_out0 = v$G59_15124_out0;
assign v$RX_4808_out0 = v$RXBIT_8913_out0;
assign v$RX_4809_out0 = v$RXBIT_8914_out0;
assign v$G34_4880_out0 = v$G33_18616_out0 || v$G35_18495_out0;
assign v$G34_4881_out0 = v$G33_18617_out0 || v$G35_18496_out0;
assign v$LOADA_5145_out0 = v$IR2$FPU$LOADA_15268_out0;
assign v$LOADA_5146_out0 = v$IR2$FPU$LOADA_15269_out0;
assign v$S_5733_out0 = v$_18018_out0;
assign v$S_5734_out0 = v$_18019_out0;
assign v$G9_6337_out0 = ((v$G8_12296_out0 && !v$OddParity_10686_out0) || (!v$G8_12296_out0) && v$OddParity_10686_out0);
assign v$G9_6338_out0 = ((v$G8_12297_out0 && !v$OddParity_10687_out0) || (!v$G8_12297_out0) && v$OddParity_10687_out0);
assign v$PIN_6637_out0 = v$_1669_out0;
assign v$PIN_6643_out0 = v$_1670_out0;
assign v$NP_7258_out0 = v$G45_16900_out0;
assign v$NP_7259_out0 = v$G45_16901_out0;
assign v$EQ1_7789_out0 = v$OUT_5002_out0 == 5'h0;
assign v$OPCODE_7892_out0 = v$_4997_out0;
assign v$OPCODE_7893_out0 = v$_4998_out0;
assign v$SHIFT_8028_out0 = v$_16737_out0;
assign v$SHIFT_8029_out0 = v$_16738_out0;
assign v$B1_8123_out0 = v$_11022_out0;
assign v$B1_8126_out0 = v$_11025_out0;
assign v$_8454_out0 = v$_12862_out1[1:0];
assign v$_8454_out1 = v$_12862_out1[3:2];
assign v$_8457_out0 = v$_12865_out1[1:0];
assign v$_8457_out1 = v$_12865_out1[3:2];
assign v$_8460_out0 = v$_12868_out1[1:0];
assign v$_8460_out1 = v$_12868_out1[3:2];
assign v$_8463_out0 = v$_12871_out1[1:0];
assign v$_8463_out1 = v$_12871_out1[3:2];
assign v$B13_8675_out0 = v$_17325_out0;
assign v$B13_8678_out0 = v$_17328_out0;
assign v$G17_8830_out0 = v$G13_13444_out0 || v$G11_8263_out0;
assign v$G17_8831_out0 = v$G13_13445_out0 || v$G11_8264_out0;
assign v$RXFlagSet_9108_out0 = v$G53_12714_out0;
assign v$RXFlagSet_9109_out0 = v$G53_12715_out0;
assign v$B11_9116_out0 = v$_9497_out1;
assign v$B11_9119_out0 = v$_9500_out1;
assign v$G24_9618_out0 = v$NQ3_1491_out0 && v$G25_18095_out0;
assign v$G24_9619_out0 = v$NQ3_1492_out0 && v$G25_18096_out0;
assign v$EQ10_9866_out0 = v$IR2$FPU$OP_1687_out0 == 2'h3;
assign v$EQ10_9867_out0 = v$IR2$FPU$OP_1688_out0 == 2'h3;
assign v$B10_9877_out0 = v$_9497_out0;
assign v$B10_9880_out0 = v$_9500_out0;
assign v$G27_10235_out0 = v$S_4025_out0 && v$NQ2_18563_out0;
assign v$G27_10236_out0 = v$S_4026_out0 && v$NQ2_18564_out0;
assign v$G18_10254_out0 = v$G16_3520_out0 || v$G9_1184_out0;
assign v$G18_10255_out0 = v$G16_3521_out0 || v$G9_1185_out0;
assign v$G70_10280_out0 = v$S_4025_out0 && v$EQ6_1566_out0;
assign v$G70_10281_out0 = v$S_4026_out0 && v$EQ6_1567_out0;
assign v$G24_10343_out0 = v$G7_12647_out0 || v$G8_4819_out0;
assign v$G24_10344_out0 = v$G7_12648_out0 || v$G8_4820_out0;
assign v$IR15_10688_out0 = v$IR2$15_7435_out0;
assign v$IR15_10689_out0 = v$IR2$15_7436_out0;
assign v$B22_10805_out0 = v$_9381_out0;
assign v$B22_10808_out0 = v$_9384_out0;
assign v$G46_10902_out0 = ! v$S_4025_out0;
assign v$G46_10903_out0 = ! v$S_4026_out0;
assign v$LOAD_11702_out0 = v$IR2$FPU$LOAD_4231_out0;
assign v$LOAD_11703_out0 = v$IR2$FPU$LOAD_4232_out0;
assign v$G20_11711_out0 = v$G23_9602_out0 && v$F2_12097_out0;
assign v$IR2$FULL$OP$CODE_11820_out0 = v$SEL3_16650_out0;
assign v$IR2$FULL$OP$CODE_11821_out0 = v$SEL3_16651_out0;
assign v$CLK4_12213_out0 = v$G2_18697_out0;
assign v$CLK4_12214_out0 = v$G2_18698_out0;
assign v$G20_12740_out0 = v$G15_1868_out0 || v$G12_1820_out0;
assign v$G20_12741_out0 = v$G15_1869_out0 || v$G12_1821_out0;
assign v$SHIFTEN_12766_out0 = v$G57_13452_out0;
assign v$SHIFTEN_12767_out0 = v$G57_13453_out0;
assign v$_12842_out0 = v$_12862_out0[1:0];
assign v$_12842_out1 = v$_12862_out0[3:2];
assign v$_12845_out0 = v$_12865_out0[1:0];
assign v$_12845_out1 = v$_12865_out0[3:2];
assign v$_12848_out0 = v$_12868_out0[1:0];
assign v$_12848_out1 = v$_12868_out0[3:2];
assign v$_12851_out0 = v$_12871_out0[1:0];
assign v$_12851_out1 = v$_12871_out0[3:2];
assign v$_12860_out0 = v$PIN_6634_out0[3:0];
assign v$_12860_out1 = v$PIN_6634_out0[7:4];
assign v$_12861_out0 = v$PIN_6635_out0[3:0];
assign v$_12861_out1 = v$PIN_6635_out0[7:4];
assign v$_12864_out0 = v$PIN_6638_out0[3:0];
assign v$_12864_out1 = v$PIN_6638_out0[7:4];
assign v$_12866_out0 = v$PIN_6640_out0[3:0];
assign v$_12866_out1 = v$PIN_6640_out0[7:4];
assign v$_12867_out0 = v$PIN_6641_out0[3:0];
assign v$_12867_out1 = v$PIN_6641_out0[7:4];
assign v$_12870_out0 = v$PIN_6644_out0[3:0];
assign v$_12870_out1 = v$PIN_6644_out0[7:4];
assign v$B8_13138_out0 = v$_6898_out1;
assign v$B8_13141_out0 = v$_6901_out1;
assign v$B_13212_out0 = v$_6990_out0;
assign v$B_13213_out0 = v$_6991_out0;
assign v$G54_14197_out0 = v$G28_15633_out0 || v$HALT$PREV_10386_out0;
assign v$G54_14198_out0 = v$G28_15634_out0 || v$HALT$PREV_10387_out0;
assign v$G21_14245_out0 = v$G14_12046_out0 || v$G10_1998_out0;
assign v$G21_14246_out0 = v$G14_12047_out0 || v$G10_1999_out0;
assign v$B4_14663_out0 = v$_6977_out0;
assign v$B4_14666_out0 = v$_6980_out0;
assign v$G26_14899_out0 = v$G3_17452_out0 || v$G4_1329_out0;
assign v$G26_14900_out0 = v$G3_17453_out0 || v$G4_1330_out0;
assign v$G66_15270_out0 = ((v$ODDPARITY_15928_out0 && !v$EVENPARITY_13588_out0) || (!v$ODDPARITY_15928_out0) && v$EVENPARITY_13588_out0);
assign v$G66_15271_out0 = ((v$ODDPARITY_15929_out0 && !v$EVENPARITY_13589_out0) || (!v$ODDPARITY_15929_out0) && v$EVENPARITY_13589_out0);
assign v$B17_15535_out0 = v$_13180_out1;
assign v$B17_15538_out0 = v$_13183_out1;
assign v$G46_16116_out0 = v$G55_5049_out0 || v$G47_5419_out0;
assign v$G46_16117_out0 = v$G55_5050_out0 || v$G47_5420_out0;
assign v$ParityCheck_16120_out0 = v$G57_8978_out0;
assign v$ParityCheck_16121_out0 = v$G57_8979_out0;
assign v$G32_16334_out0 = v$G35_12635_out0 || v$G40_15130_out0;
assign v$G32_16335_out0 = v$G35_12636_out0 || v$G40_15131_out0;
assign v$B16_16414_out0 = v$_13180_out0;
assign v$B16_16417_out0 = v$_13183_out0;
assign v$RXReset_16530_out0 = v$G64_7783_out0;
assign v$RXReset_16531_out0 = v$G64_7784_out0;
assign v$G55_16658_out0 = v$EQ2_18657_out0 || v$G56_648_out0;
assign v$G55_16659_out0 = v$EQ2_18658_out0 || v$G56_649_out0;
assign v$RAMDOUT_16779_out0 = v$DATA$OUT_1307_out0;
assign v$RAMDOUT_16780_out0 = v$DATA$OUT_1308_out0;
assign v$B19_16789_out0 = v$_16589_out0;
assign v$B19_16792_out0 = v$_16592_out0;
assign v$G63_16810_out0 = v$G57_13452_out0 && v$SERIALIN_5728_out0;
assign v$G63_16811_out0 = v$G57_13453_out0 && v$SERIALIN_5729_out0;
assign v$B7_17040_out0 = v$_6898_out0;
assign v$B7_17043_out0 = v$_6901_out0;
assign v$MUX4_17084_out0 = v$G47_1531_out0 ? v$C4_2920_out0 : v$G39_6045_out0;
assign v$MUX4_17085_out0 = v$G47_1532_out0 ? v$C4_2921_out0 : v$G39_6046_out0;
assign v$G3_17694_out0 = ! v$R_1590_out0;
assign v$G9_17710_out0 = ! v$EQ7_18631_out0;
assign v$G9_17711_out0 = ! v$EQ7_18632_out0;
assign v$IR2_17953_out0 = v$IR2_7773_out0;
assign v$IR2_17954_out0 = v$IR2_7774_out0;
assign v$B5_18374_out0 = v$_6977_out1;
assign v$B5_18377_out0 = v$_6980_out1;
assign v$CHECKPARITY_1327_out0 = v$ParityCheck_16120_out0;
assign v$CHECKPARITY_1328_out0 = v$ParityCheck_16121_out0;
assign v$1_1533_out0 = v$IR2_17953_out0[8:8];
assign v$1_1534_out0 = v$IR2_17954_out0[8:8];
assign v$_1641_out0 = v$_12842_out1[0:0];
assign v$_1641_out1 = v$_12842_out1[1:1];
assign v$_1644_out0 = v$_12845_out1[0:0];
assign v$_1644_out1 = v$_12845_out1[1:1];
assign v$_1647_out0 = v$_12848_out1[0:0];
assign v$_1647_out1 = v$_12848_out1[1:1];
assign v$_1650_out0 = v$_12851_out1[0:0];
assign v$_1650_out1 = v$_12851_out1[1:1];
assign v$G65_2460_out0 = v$EQ5_9106_out0 && v$G66_15270_out0;
assign v$G65_2461_out0 = v$EQ5_9107_out0 && v$G66_15271_out0;
assign v$CLK4_2531_out0 = v$CLK4_12213_out0;
assign v$CLK4_2532_out0 = v$CLK4_12214_out0;
assign v$B_2701_out0 = v$B7_17040_out0;
assign v$B_2702_out0 = v$B1_8123_out0;
assign v$B_2703_out0 = v$B14_4002_out0;
assign v$B_2705_out0 = v$B8_13138_out0;
assign v$B_2706_out0 = v$B17_15535_out0;
assign v$B_2707_out0 = v$B23_1283_out0;
assign v$B_2709_out0 = v$B13_8675_out0;
assign v$B_2710_out0 = v$B4_14663_out0;
assign v$B_2711_out0 = v$B19_16789_out0;
assign v$B_2712_out0 = v$B22_10805_out0;
assign v$B_2714_out0 = v$B10_9877_out0;
assign v$B_2715_out0 = v$B20_3943_out0;
assign v$B_2716_out0 = v$B2_3113_out0;
assign v$B_2717_out0 = v$B11_9116_out0;
assign v$B_2718_out0 = v$B5_18374_out0;
assign v$B_2719_out0 = v$B16_16414_out0;
assign v$B_2773_out0 = v$B7_17043_out0;
assign v$B_2774_out0 = v$B1_8126_out0;
assign v$B_2775_out0 = v$B14_4005_out0;
assign v$B_2777_out0 = v$B8_13141_out0;
assign v$B_2778_out0 = v$B17_15538_out0;
assign v$B_2779_out0 = v$B23_1286_out0;
assign v$B_2781_out0 = v$B13_8678_out0;
assign v$B_2782_out0 = v$B4_14666_out0;
assign v$B_2783_out0 = v$B19_16792_out0;
assign v$B_2784_out0 = v$B22_10808_out0;
assign v$B_2786_out0 = v$B10_9880_out0;
assign v$B_2787_out0 = v$B20_3946_out0;
assign v$B_2788_out0 = v$B2_3116_out0;
assign v$B_2789_out0 = v$B11_9119_out0;
assign v$B_2790_out0 = v$B5_18377_out0;
assign v$B_2791_out0 = v$B16_16417_out0;
assign v$G10_2906_out0 = ((v$G9_6337_out0 && !v$RceivedParity_18539_out0) || (!v$G9_6337_out0) && v$RceivedParity_18539_out0);
assign v$G10_2907_out0 = ((v$G9_6338_out0 && !v$RceivedParity_18540_out0) || (!v$G9_6338_out0) && v$RceivedParity_18540_out0);
assign v$SEL6_3008_out0 = v$IR1_4156_out0[1:0];
assign v$SEL6_3009_out0 = v$IR1_4157_out0[1:0];
assign v$G11_3251_out0 = v$IR2$FPU$LOAD_4231_out0 && v$G12_3615_out0;
assign v$G11_3252_out0 = v$IR2$FPU$LOAD_4232_out0 && v$G12_3616_out0;
assign v$SEL2_3714_out0 = v$IR1_4156_out0[8:8];
assign v$SEL2_3715_out0 = v$IR1_4157_out0[8:8];
assign v$Q2P_4160_out0 = v$G24_9618_out0;
assign v$Q2P_4161_out0 = v$G24_9619_out0;
assign v$S_4239_out0 = v$S_5733_out0;
assign v$S_4240_out0 = v$S_5734_out0;
assign v$LOADA_5076_out0 = v$LOADA_5145_out0;
assign v$LOADA_5077_out0 = v$LOADA_5146_out0;
assign v$C_6062_out0 = v$C_3198_out0;
assign v$C_6063_out0 = v$C_3199_out0;
assign v$LOAD_6190_out0 = v$LOAD_11702_out0;
assign v$LOAD_6191_out0 = v$LOAD_11703_out0;
assign v$EQ6_6411_out0 = v$IR2$FULL$OP$CODE_11820_out0 == 4'h7;
assign v$EQ6_6412_out0 = v$IR2$FULL$OP$CODE_11821_out0 == 4'h7;
assign v$SHIFT_7019_out0 = v$SHIFT_8028_out0;
assign v$SHIFT_7020_out0 = v$SHIFT_8029_out0;
assign v$_7658_out0 = v$_12842_out0[0:0];
assign v$_7658_out1 = v$_12842_out0[1:1];
assign v$_7661_out0 = v$_12845_out0[0:0];
assign v$_7661_out1 = v$_12845_out0[1:1];
assign v$_7664_out0 = v$_12848_out0[0:0];
assign v$_7664_out1 = v$_12848_out0[1:1];
assign v$_7667_out0 = v$_12851_out0[0:0];
assign v$_7667_out1 = v$_12851_out0[1:1];
assign v$SEL9_7983_out0 = v$IR1_4156_out0[11:10];
assign v$SEL9_7984_out0 = v$IR1_4157_out0[11:10];
assign v$G54_8133_out0 = v$G55_16658_out0 || v$G63_16810_out0;
assign v$G54_8134_out0 = v$G55_16659_out0 || v$G63_16811_out0;
assign v$_8452_out0 = v$_12860_out1[1:0];
assign v$_8452_out1 = v$_12860_out1[3:2];
assign v$_8453_out0 = v$_12861_out1[1:0];
assign v$_8453_out1 = v$_12861_out1[3:2];
assign v$_8456_out0 = v$_12864_out1[1:0];
assign v$_8456_out1 = v$_12864_out1[3:2];
assign v$_8458_out0 = v$_12866_out1[1:0];
assign v$_8458_out1 = v$_12866_out1[3:2];
assign v$_8459_out0 = v$_12867_out1[1:0];
assign v$_8459_out1 = v$_12867_out1[3:2];
assign v$_8462_out0 = v$_12870_out1[1:0];
assign v$_8462_out1 = v$_12870_out1[3:2];
assign v$R_8778_out0 = v$RX_4808_out0;
assign v$R_8779_out0 = v$RX_4809_out0;
assign v$SEL1_8796_out0 = v$IR1_4156_out0[15:12];
assign v$SEL1_8797_out0 = v$IR1_4157_out0[15:12];
assign v$6_9868_out0 = v$IR2_17953_out0[7:7];
assign v$6_9869_out0 = v$IR2_17954_out0[7:7];
assign v$SHIFTEN_10282_out0 = v$SHIFTEN_12766_out0;
assign v$SHIFTEN_10283_out0 = v$SHIFTEN_12767_out0;
assign v$G26_10320_out0 = v$G22_5463_out0 || v$G20_11711_out0;
assign v$G28_10803_out0 = v$G27_260_out0 || v$G26_14899_out0;
assign v$G28_10804_out0 = v$G27_261_out0 || v$G26_14900_out0;
assign v$FINISHED_10861_out0 = v$EQ1_7789_out0;
assign v$IR15_10986_out0 = v$IR15_10688_out0;
assign v$IR15_10987_out0 = v$IR15_10689_out0;
assign v$G18_11028_out0 = v$IR2$FPU$LOAD_4231_out0 && v$EQ10_9866_out0;
assign v$G18_11029_out0 = v$IR2$FPU$LOAD_4232_out0 && v$EQ10_9867_out0;
assign v$Q3P_11672_out0 = v$MUX4_17084_out0;
assign v$Q3P_11673_out0 = v$MUX4_17085_out0;
assign v$IR2$VALID_11794_out0 = v$IR2$VALID_4217_out0;
assign v$IR2$VALID_11795_out0 = v$IR2$VALID_4218_out0;
assign v$G11_11845_out0 = v$Q3_18425_out0 && v$G52_2971_out0;
assign v$G11_11846_out0 = v$Q3_18426_out0 && v$G52_2972_out0;
assign v$_11860_out0 = v$_8454_out1[0:0];
assign v$_11860_out1 = v$_8454_out1[1:1];
assign v$_11863_out0 = v$_8457_out1[0:0];
assign v$_11863_out1 = v$_8457_out1[1:1];
assign v$_11866_out0 = v$_8460_out1[0:0];
assign v$_11866_out1 = v$_8460_out1[1:1];
assign v$_11869_out0 = v$_8463_out1[0:0];
assign v$_11869_out1 = v$_8463_out1[1:1];
assign v$EQ11_11882_out0 = v$IR2$FULL$OP$CODE_11820_out0 == 4'h1;
assign v$EQ11_11883_out0 = v$IR2$FULL$OP$CODE_11821_out0 == 4'h1;
assign v$SEL11_12201_out0 = v$IR2_17953_out0[7:7];
assign v$SEL11_12202_out0 = v$IR2_17954_out0[7:7];
assign v$_12228_out0 = { v$K_301_out0,v$C1_15804_out0 };
assign v$_12229_out0 = { v$K_302_out0,v$C1_15805_out0 };
assign v$5_12290_out0 = v$IR2_17953_out0[9:9];
assign v$5_12291_out0 = v$IR2_17954_out0[9:9];
assign v$EQ4_12725_out0 = v$IR2_17953_out0 == 16'h7000;
assign v$EQ4_12726_out0 = v$IR2_17954_out0 == 16'h7000;
assign v$2_12738_out0 = v$IR2_17953_out0[11:10];
assign v$2_12739_out0 = v$IR2_17954_out0[11:10];
assign v$SEL10_12823_out0 = v$IR2_17953_out0[9:8];
assign v$SEL10_12824_out0 = v$IR2_17954_out0[9:8];
assign v$_12840_out0 = v$_12860_out0[1:0];
assign v$_12840_out1 = v$_12860_out0[3:2];
assign v$_12841_out0 = v$_12861_out0[1:0];
assign v$_12841_out1 = v$_12861_out0[3:2];
assign v$_12844_out0 = v$_12864_out0[1:0];
assign v$_12844_out1 = v$_12864_out0[3:2];
assign v$_12846_out0 = v$_12866_out0[1:0];
assign v$_12846_out1 = v$_12866_out0[3:2];
assign v$_12847_out0 = v$_12867_out0[1:0];
assign v$_12847_out1 = v$_12867_out0[3:2];
assign v$_12850_out0 = v$_12870_out0[1:0];
assign v$_12850_out1 = v$_12870_out0[3:2];
assign v$_12863_out0 = v$PIN_6637_out0[3:0];
assign v$_12863_out1 = v$PIN_6637_out0[7:4];
assign v$_12869_out0 = v$PIN_6643_out0[3:0];
assign v$_12869_out1 = v$PIN_6643_out0[7:4];
assign v$G1_12986_out0 = v$STATE_16017_out0 && v$G3_17694_out0;
assign v$EQ12_13260_out0 = v$IR2$FULL$OP$CODE_11820_out0 == 4'h1;
assign v$EQ12_13261_out0 = v$IR2$FULL$OP$CODE_11821_out0 == 4'h1;
assign v$3_13396_out0 = v$IR2_17953_out0[5:2];
assign v$3_13397_out0 = v$IR2_17954_out0[5:2];
assign v$Q3P_13809_out0 = v$G32_16334_out0;
assign v$Q3P_13810_out0 = v$G32_16335_out0;
assign v$G29_13993_out0 = v$G25_1309_out0 || v$G24_10343_out0;
assign v$G29_13994_out0 = v$G25_1310_out0 || v$G24_10344_out0;
assign v$7_14010_out0 = v$IR2_17953_out0[1:0];
assign v$7_14011_out0 = v$IR2_17954_out0[1:0];
assign v$9_14315_out0 = v$IR2_17953_out0[15:12];
assign v$9_14316_out0 = v$IR2_17954_out0[15:12];
assign v$G2_14499_out0 = ((v$RX_43_out0 && !v$FF3_7331_out0) || (!v$RX_43_out0) && v$FF3_7331_out0);
assign v$G2_14500_out0 = ((v$RX_44_out0 && !v$FF3_7332_out0) || (!v$RX_44_out0) && v$FF3_7332_out0);
assign v$_14513_out0 = v$_8454_out0[0:0];
assign v$_14513_out1 = v$_8454_out0[1:1];
assign v$_14516_out0 = v$_8457_out0[0:0];
assign v$_14516_out1 = v$_8457_out0[1:1];
assign v$_14519_out0 = v$_8460_out0[0:0];
assign v$_14519_out1 = v$_8460_out0[1:1];
assign v$_14522_out0 = v$_8463_out0[0:0];
assign v$_14522_out1 = v$_8463_out0[1:1];
assign v$B_14623_out0 = v$B_13212_out0;
assign v$B_14624_out0 = v$B_13213_out0;
assign v$RXSET_14687_out0 = v$RXFlagSet_9108_out0;
assign v$RXSET_14688_out0 = v$RXFlagSet_9109_out0;
assign v$RXINTERRUPT_14845_out0 = v$RXReset_16530_out0;
assign v$RXINTERRUPT_14846_out0 = v$RXReset_16531_out0;
assign v$SEL8_15116_out0 = v$IR1_4156_out0[9:8];
assign v$SEL8_15117_out0 = v$IR1_4157_out0[9:8];
assign v$4_15164_out0 = v$IR2_17953_out0[6:6];
assign v$4_15165_out0 = v$IR2_17954_out0[6:6];
assign v$MUX1_15262_out0 = v$G54_14197_out0 ? v$REG3_2822_out0 : v$R_18353_out0;
assign v$MUX1_15263_out0 = v$G54_14198_out0 ? v$REG3_2823_out0 : v$R_18354_out0;
assign v$8_15540_out0 = v$IR2_17953_out0[15:15];
assign v$8_15541_out0 = v$IR2_17954_out0[15:15];
assign v$SEL7_15615_out0 = v$IR1_4156_out0[9:9];
assign v$SEL7_15616_out0 = v$IR1_4157_out0[9:9];
assign v$G53_15830_out0 = v$G17_362_out0 || v$NQ3_2998_out0;
assign v$G53_15831_out0 = v$G17_363_out0 || v$NQ3_2999_out0;
assign v$G22_15852_out0 = v$G20_12740_out0 || v$G21_14245_out0;
assign v$G22_15853_out0 = v$G20_12741_out0 || v$G21_14246_out0;
assign v$G19_15948_out0 = v$G17_8830_out0 || v$G18_10254_out0;
assign v$G19_15949_out0 = v$G17_8831_out0 || v$G18_10255_out0;
assign v$G26_16025_out0 = v$NQ3_2998_out0 || v$G27_10235_out0;
assign v$G26_16026_out0 = v$NQ3_2999_out0 || v$G27_10236_out0;
assign v$EQ1_16122_out0 = v$OPCODE_7892_out0 == 3'h4;
assign v$EQ1_16123_out0 = v$OPCODE_7893_out0 == 3'h4;
assign v$ShiftOut_16343_out0 = v$G46_16116_out0;
assign v$ShiftOut_16344_out0 = v$G46_16117_out0;
assign v$OP_17642_out0 = v$OP_1872_out0;
assign v$OP_17643_out0 = v$OP_1873_out0;
assign v$G10_18186_out0 = v$NP_7258_out0 && v$G11_4865_out0;
assign v$G10_18187_out0 = v$NP_7259_out0 && v$G11_4866_out0;
assign v$NS_18201_out0 = v$G46_10902_out0;
assign v$NS_18202_out0 = v$G46_10903_out0;
assign v$EQ9_18283_out0 = v$IR2$FULL$OP$CODE_11820_out0 == 4'h1;
assign v$EQ9_18284_out0 = v$IR2$FULL$OP$CODE_11821_out0 == 4'h1;
assign v$EQ1_18594_out0 = v$IR2$FULL$OP$CODE_11820_out0 == 4'h1;
assign v$EQ1_18595_out0 = v$IR2$FULL$OP$CODE_11821_out0 == 4'h1;
assign v$IR1$S$WB_322_out0 = v$SEL2_3714_out0;
assign v$IR1$S$WB_323_out0 = v$SEL2_3715_out0;
assign v$RXSHIFT_674_out0 = v$ShiftOut_16343_out0;
assign v$RXSHIFT_675_out0 = v$ShiftOut_16344_out0;
assign v$G69_1206_out0 = ! v$R_8778_out0;
assign v$G69_1207_out0 = ! v$R_8779_out0;
assign v$R_1487_out0 = v$FINISHED_10861_out0;
assign v$_1639_out0 = v$_12840_out1[0:0];
assign v$_1639_out1 = v$_12840_out1[1:1];
assign v$_1640_out0 = v$_12841_out1[0:0];
assign v$_1640_out1 = v$_12841_out1[1:1];
assign v$_1643_out0 = v$_12844_out1[0:0];
assign v$_1643_out1 = v$_12844_out1[1:1];
assign v$_1645_out0 = v$_12846_out1[0:0];
assign v$_1645_out1 = v$_12846_out1[1:1];
assign v$_1646_out0 = v$_12847_out1[0:0];
assign v$_1646_out1 = v$_12847_out1[1:1];
assign v$_1649_out0 = v$_12850_out1[0:0];
assign v$_1649_out1 = v$_12850_out1[1:1];
assign v$EQ1_2516_out0 = v$OP_17642_out0 == 3'h4;
assign v$EQ1_2517_out0 = v$OP_17643_out0 == 3'h4;
assign v$IR2$OPCODE_2569_out0 = v$9_14315_out0;
assign v$IR2$OPCODE_2570_out0 = v$9_14316_out0;
assign v$MUX1_2584_out0 = v$G2_15035_out0 ? v$SIN_93_out0 : v$_7658_out0;
assign v$MUX1_2587_out0 = v$G2_15038_out0 ? v$SIN_96_out0 : v$_7661_out0;
assign v$MUX1_2590_out0 = v$G2_15041_out0 ? v$SIN_99_out0 : v$_7664_out0;
assign v$MUX1_2593_out0 = v$G2_15044_out0 ? v$SIN_102_out0 : v$_7667_out0;
assign v$_2652_out0 = v$OP_17642_out0[0:0];
assign v$_2653_out0 = v$OP_17643_out0[0:0];
assign v$IR2$FPU$OP_2881_out0 = v$SEL10_12823_out0;
assign v$IR2$FPU$OP_2882_out0 = v$SEL10_12824_out0;
assign v$IR2$IS$FPU_2929_out0 = v$EQ12_13260_out0;
assign v$IR2$IS$FPU_2930_out0 = v$EQ12_13261_out0;
assign v$_2982_out0 = v$OP_17642_out0[2:2];
assign v$_2983_out0 = v$OP_17643_out0[2:2];
assign v$IR2$N_2984_out0 = v$3_13396_out0;
assign v$IR2$N_2985_out0 = v$3_13397_out0;
assign v$MUX8_3605_out0 = v$G2_15035_out0 ? v$FF2_14784_out0 : v$_14513_out0;
assign v$MUX8_3608_out0 = v$G2_15038_out0 ? v$FF2_14787_out0 : v$_14516_out0;
assign v$MUX8_3611_out0 = v$G2_15041_out0 ? v$FF2_14790_out0 : v$_14519_out0;
assign v$MUX8_3614_out0 = v$G2_15044_out0 ? v$FF2_14793_out0 : v$_14522_out0;
assign v$B_3704_out0 = v$B_14623_out0;
assign v$B_3705_out0 = v$B_14624_out0;
assign v$G23_4385_out0 = v$G19_15948_out0 || v$G22_15852_out0;
assign v$G23_4386_out0 = v$G19_15949_out0 || v$G22_15853_out0;
assign v$IR2$D_4898_out0 = v$2_12738_out0;
assign v$IR2$D_4899_out0 = v$2_12739_out0;
assign v$RXset_5101_out0 = v$RXSET_14687_out0;
assign v$RXset_5102_out0 = v$RXSET_14688_out0;
assign v$MUX1_5137_out0 = v$FINISHED_10861_out0 ? v$C1_15678_out0 : v$OUT_5002_out0;
assign v$EQ4_5414_out0 = v$SEL8_15116_out0 == 2'h2;
assign v$EQ4_5415_out0 = v$SEL8_15117_out0 == 2'h2;
assign v$IR1$RD_5489_out0 = v$SEL9_7983_out0;
assign v$IR1$RD_5490_out0 = v$SEL9_7984_out0;
assign v$IR2$U_5904_out0 = v$4_15164_out0;
assign v$IR2$U_5905_out0 = v$4_15165_out0;
assign v$G14_6127_out0 = v$G15_4205_out0 && v$G53_15830_out0;
assign v$G14_6128_out0 = v$G15_4206_out0 && v$G53_15831_out0;
assign v$ISMOV_6670_out0 = v$EQ1_16122_out0;
assign v$ISMOV_6671_out0 = v$EQ1_16123_out0;
assign v$FINISHED_7003_out0 = v$FINISHED_10861_out0;
assign v$SHIFTEN_7092_out0 = v$SHIFTEN_10282_out0;
assign v$SHIFTEN_7093_out0 = v$SHIFTEN_10283_out0;
assign v$G2_7578_out0 = v$G1_12986_out0 || v$S_8021_out0;
assign v$_7656_out0 = v$_12840_out0[0:0];
assign v$_7656_out1 = v$_12840_out0[1:1];
assign v$_7657_out0 = v$_12841_out0[0:0];
assign v$_7657_out1 = v$_12841_out0[1:1];
assign v$_7660_out0 = v$_12844_out0[0:0];
assign v$_7660_out1 = v$_12844_out0[1:1];
assign v$_7662_out0 = v$_12846_out0[0:0];
assign v$_7662_out1 = v$_12846_out0[1:1];
assign v$_7663_out0 = v$_12847_out0[0:0];
assign v$_7663_out1 = v$_12847_out0[1:1];
assign v$_7666_out0 = v$_12850_out0[0:0];
assign v$_7666_out1 = v$_12850_out0[1:1];
assign v$EQ2_7952_out0 = v$OP_17642_out0 == 3'h5;
assign v$EQ2_7953_out0 = v$OP_17643_out0 == 3'h5;
assign v$S_8167_out0 = v$S_4239_out0;
assign v$S_8168_out0 = v$S_4240_out0;
assign v$G69_8210_out0 = v$EQ7_231_out0 && v$NS_18201_out0;
assign v$G69_8211_out0 = v$EQ7_232_out0 && v$NS_18202_out0;
assign v$_8232_out0 = v$OP_17642_out0[1:1];
assign v$_8233_out0 = v$OP_17643_out0[1:1];
assign v$STOP$2_8234_out0 = v$EQ4_12725_out0;
assign v$STOP$2_8235_out0 = v$EQ4_12726_out0;
assign v$_8455_out0 = v$_12863_out1[1:0];
assign v$_8455_out1 = v$_12863_out1[3:2];
assign v$_8461_out0 = v$_12869_out1[1:0];
assign v$_8461_out1 = v$_12869_out1[3:2];
assign v$IR2$M_8832_out0 = v$7_14010_out0;
assign v$IR2$M_8833_out0 = v$7_14011_out0;
assign v$G8_9504_out0 = v$G9_13446_out0 && v$G11_11845_out0;
assign v$G8_9505_out0 = v$G9_13447_out0 && v$G11_11846_out0;
assign v$MUX5_9526_out0 = v$G2_15035_out0 ? v$FF5_1756_out0 : v$_7658_out1;
assign v$MUX5_9529_out0 = v$G2_15038_out0 ? v$FF5_1759_out0 : v$_7661_out1;
assign v$MUX5_9532_out0 = v$G2_15041_out0 ? v$FF5_1762_out0 : v$_7664_out1;
assign v$MUX5_9535_out0 = v$G2_15044_out0 ? v$FF5_1765_out0 : v$_7667_out1;
assign v$IR1$OPCODE_9564_out0 = v$SEL1_8796_out0;
assign v$IR1$OPCODE_9565_out0 = v$SEL1_8797_out0;
assign v$_9580_out0 = v$OP_17642_out0[2:2];
assign v$_9581_out0 = v$OP_17643_out0[2:2];
assign v$C_9609_out0 = v$C_6062_out0;
assign v$C_9610_out0 = v$C_6063_out0;
assign v$MUX3_9952_out0 = v$G2_15035_out0 ? v$FF7_8300_out0 : v$_14513_out1;
assign v$MUX3_9955_out0 = v$G2_15038_out0 ? v$FF7_8303_out0 : v$_14516_out1;
assign v$MUX3_9958_out0 = v$G2_15041_out0 ? v$FF7_8306_out0 : v$_14519_out1;
assign v$MUX3_9961_out0 = v$G2_15044_out0 ? v$FF7_8309_out0 : v$_14522_out1;
assign v$IR1$C$L_10053_out0 = v$SEL7_15615_out0;
assign v$IR1$C$L_10054_out0 = v$SEL7_15616_out0;
assign v$G10_10271_out0 = v$EQ6_6411_out0 && v$G9_17710_out0;
assign v$G10_10272_out0 = v$EQ6_6412_out0 && v$G9_17711_out0;
assign v$_10278_out0 = v$OP_17642_out0[1:1];
assign v$_10279_out0 = v$OP_17643_out0[1:1];
assign v$MUX6_10390_out0 = v$G2_15035_out0 ? v$FF1_16076_out0 : v$_1641_out1;
assign v$MUX6_10393_out0 = v$G2_15038_out0 ? v$FF1_16079_out0 : v$_1644_out1;
assign v$MUX6_10396_out0 = v$G2_15041_out0 ? v$FF1_16082_out0 : v$_1647_out1;
assign v$MUX6_10399_out0 = v$G2_15044_out0 ? v$FF1_16085_out0 : v$_1650_out1;
assign v$IR2$FPU$L_10744_out0 = v$SEL11_12201_out0;
assign v$IR2$FPU$L_10745_out0 = v$SEL11_12202_out0;
assign v$G62_11755_out0 = v$G61_11603_out0 && v$CLK4_2531_out0;
assign v$G62_11756_out0 = v$G61_11604_out0 && v$CLK4_2532_out0;
assign v$_11858_out0 = v$_8452_out1[0:0];
assign v$_11858_out1 = v$_8452_out1[1:1];
assign v$_11859_out0 = v$_8453_out1[0:0];
assign v$_11859_out1 = v$_8453_out1[1:1];
assign v$_11862_out0 = v$_8456_out1[0:0];
assign v$_11862_out1 = v$_8456_out1[1:1];
assign v$_11864_out0 = v$_8458_out1[0:0];
assign v$_11864_out1 = v$_8458_out1[1:1];
assign v$_11865_out0 = v$_8459_out1[0:0];
assign v$_11865_out1 = v$_8459_out1[1:1];
assign v$_11868_out0 = v$_8462_out1[0:0];
assign v$_11868_out1 = v$_8462_out1[1:1];
assign v$G1_12223_out0 = v$FINISHED_10861_out0 || v$CALCULATING_1493_out0;
assign v$G20_12292_out0 = ! v$LOAD_6190_out0;
assign v$G20_12293_out0 = ! v$LOAD_6191_out0;
assign v$IR2$L_12464_out0 = v$5_12290_out0;
assign v$IR2$L_12465_out0 = v$5_12291_out0;
assign v$_12843_out0 = v$_12863_out0[1:0];
assign v$_12843_out1 = v$_12863_out0[3:2];
assign v$_12849_out0 = v$_12869_out0[1:0];
assign v$_12849_out1 = v$_12869_out0[3:2];
assign v$_13065_out0 = { v$Q2P_4160_out0,v$Q3P_13809_out0 };
assign v$_13066_out0 = { v$Q2P_4161_out0,v$Q3P_13810_out0 };
assign v$G11_13406_out0 = ! v$LOAD_6190_out0;
assign v$G11_13407_out0 = ! v$LOAD_6191_out0;
assign v$_13691_out0 = v$OP_17642_out0[0:0];
assign v$_13692_out0 = v$OP_17643_out0[0:0];
assign v$MUX2_13821_out0 = v$G2_15035_out0 ? v$FF8_14462_out0 : v$_11860_out1;
assign v$MUX2_13824_out0 = v$G2_15038_out0 ? v$FF8_14465_out0 : v$_11863_out1;
assign v$MUX2_13827_out0 = v$G2_15041_out0 ? v$FF8_14468_out0 : v$_11866_out1;
assign v$MUX2_13830_out0 = v$G2_15044_out0 ? v$FF8_14471_out0 : v$_11869_out1;
assign v$B$IS$RD_14084_out0 = v$G11_3251_out0;
assign v$B$IS$RD_14085_out0 = v$G11_3252_out0;
assign v$_14511_out0 = v$_8452_out0[0:0];
assign v$_14511_out1 = v$_8452_out0[1:1];
assign v$_14512_out0 = v$_8453_out0[0:0];
assign v$_14512_out1 = v$_8453_out0[1:1];
assign v$_14515_out0 = v$_8456_out0[0:0];
assign v$_14515_out1 = v$_8456_out0[1:1];
assign v$_14517_out0 = v$_8458_out0[0:0];
assign v$_14517_out1 = v$_8458_out0[1:1];
assign v$_14518_out0 = v$_8459_out0[0:0];
assign v$_14518_out1 = v$_8459_out0[1:1];
assign v$_14521_out0 = v$_8462_out0[0:0];
assign v$_14521_out1 = v$_8462_out0[1:1];
assign v$G10_14588_out0 = ! v$LOADA_5076_out0;
assign v$G10_14589_out0 = ! v$LOADA_5077_out0;
assign v$IR2$W_15109_out0 = v$1_1533_out0;
assign v$IR2$W_15110_out0 = v$1_1534_out0;
assign v$G64_15260_out0 = v$G54_8133_out0 || v$G65_2460_out0;
assign v$G64_15261_out0 = v$G54_8134_out0 || v$G65_2461_out0;
assign v$RXINTERRUPT_15347_out0 = v$RXINTERRUPT_14845_out0;
assign v$RXINTERRUPT_15348_out0 = v$RXINTERRUPT_14846_out0;
assign v$EQ3_15504_out0 = v$OP_17642_out0 == 3'h7;
assign v$EQ3_15505_out0 = v$OP_17643_out0 == 3'h7;
assign v$IR2$LS_15832_out0 = v$8_15540_out0;
assign v$IR2$LS_15833_out0 = v$8_15541_out0;
assign v$G19_16043_out0 = v$EQ9_18283_out0 && v$G18_11028_out0;
assign v$G19_16044_out0 = v$EQ9_18284_out0 && v$G18_11029_out0;
assign v$G12_16252_out0 = ! v$R_8778_out0;
assign v$G12_16253_out0 = ! v$R_8779_out0;
assign v$IR1_16680_out0 = v$MUX1_15262_out0;
assign v$IR1_16681_out0 = v$MUX1_15263_out0;
assign v$MUX4_16849_out0 = v$G2_15035_out0 ? v$FF6_2623_out0 : v$_11860_out0;
assign v$MUX4_16852_out0 = v$G2_15038_out0 ? v$FF6_2626_out0 : v$_11863_out0;
assign v$MUX4_16855_out0 = v$G2_15041_out0 ? v$FF6_2629_out0 : v$_11866_out0;
assign v$MUX4_16858_out0 = v$G2_15044_out0 ? v$FF6_2632_out0 : v$_11869_out0;
assign v$IR2$P_17316_out0 = v$6_9868_out0;
assign v$IR2$P_17317_out0 = v$6_9869_out0;
assign v$E_17351_out0 = v$G2_14499_out0;
assign v$E_17352_out0 = v$G2_14500_out0;
assign v$MUX7_17905_out0 = v$G2_15035_out0 ? v$FF3_9973_out0 : v$_1641_out0;
assign v$MUX7_17908_out0 = v$G2_15038_out0 ? v$FF3_9976_out0 : v$_1644_out0;
assign v$MUX7_17911_out0 = v$G2_15041_out0 ? v$FF3_9979_out0 : v$_1647_out0;
assign v$MUX7_17914_out0 = v$G2_15044_out0 ? v$FF3_9982_out0 : v$_1650_out0;
assign v$EDGE2_18119_out0 = v$G26_10320_out0;
assign v$IR1$RM_18301_out0 = v$SEL6_3008_out0;
assign v$IR1$RM_18302_out0 = v$SEL6_3009_out0;
assign v$IR1$FPU$OP$CODE_18316_out0 = v$SEL8_15116_out0;
assign v$IR1$FPU$OP$CODE_18317_out0 = v$SEL8_15117_out0;
assign v$G24_18388_out0 = v$G25_14030_out0 && v$G26_16025_out0;
assign v$G24_18389_out0 = v$G25_14031_out0 && v$G26_16026_out0;
assign v$G37_18464_out0 = v$Q3_18425_out0 && v$NS_18201_out0;
assign v$G37_18465_out0 = v$Q3_18426_out0 && v$NS_18202_out0;
assign v$G30_18605_out0 = v$G28_10803_out0 || v$G29_13993_out0;
assign v$G30_18606_out0 = v$G28_10804_out0 || v$G29_13994_out0;
assign v$CheckParity_18678_out0 = v$CHECKPARITY_1327_out0;
assign v$CheckParity_18679_out0 = v$CHECKPARITY_1328_out0;
assign v$IR2$VALID_18756_out0 = v$IR2$VALID_11794_out0;
assign v$IR2$VALID_18757_out0 = v$IR2$VALID_11795_out0;
assign v$_304_out0 = v$IR1_16680_out0[15:12];
assign v$_305_out0 = v$IR1_16681_out0[15:12];
assign v$S_901_out0 = v$S_8167_out0;
assign v$S_902_out0 = v$S_8168_out0;
assign v$TX_1298_out0 = v$G64_15260_out0;
assign v$TX_1299_out0 = v$G64_15261_out0;
assign v$EQ16_1582_out0 = v$IR1$FPU$OP$CODE_18316_out0 == 2'h3;
assign v$EQ16_1583_out0 = v$IR1$FPU$OP$CODE_18317_out0 == 2'h3;
assign v$R_1586_out0 = v$R_1487_out0;
assign v$_1642_out0 = v$_12843_out1[0:0];
assign v$_1642_out1 = v$_12843_out1[1:1];
assign v$_1648_out0 = v$_12849_out1[0:0];
assign v$_1648_out1 = v$_12849_out1[1:1];
assign v$RXset_1701_out0 = v$RXset_5101_out0;
assign v$RXset_1702_out0 = v$RXset_5102_out0;
assign v$S_2443_out0 = v$S_8167_out0;
assign v$S_2444_out0 = v$S_8168_out0;
assign v$MUX1_2582_out0 = v$G2_15033_out0 ? v$SIN_91_out0 : v$_7656_out0;
assign v$MUX1_2583_out0 = v$G2_15034_out0 ? v$SIN_92_out0 : v$_7657_out0;
assign v$MUX1_2586_out0 = v$G2_15037_out0 ? v$SIN_95_out0 : v$_7660_out0;
assign v$MUX1_2588_out0 = v$G2_15039_out0 ? v$SIN_97_out0 : v$_7662_out0;
assign v$MUX1_2589_out0 = v$G2_15040_out0 ? v$SIN_98_out0 : v$_7663_out0;
assign v$MUX1_2592_out0 = v$G2_15043_out0 ? v$SIN_101_out0 : v$_7666_out0;
assign v$G6_3163_out0 = v$G8_9504_out0 || v$G14_6127_out0;
assign v$G6_3164_out0 = v$G8_9505_out0 || v$G14_6128_out0;
assign v$EQ7_3506_out0 = v$IR2$OPCODE_2569_out0 == 4'h1;
assign v$EQ7_3507_out0 = v$IR2$OPCODE_2570_out0 == 4'h1;
assign v$MUX8_3603_out0 = v$G2_15033_out0 ? v$FF2_14782_out0 : v$_14511_out0;
assign v$MUX8_3604_out0 = v$G2_15034_out0 ? v$FF2_14783_out0 : v$_14512_out0;
assign v$MUX8_3607_out0 = v$G2_15037_out0 ? v$FF2_14786_out0 : v$_14515_out0;
assign v$MUX8_3609_out0 = v$G2_15039_out0 ? v$FF2_14788_out0 : v$_14517_out0;
assign v$MUX8_3610_out0 = v$G2_15040_out0 ? v$FF2_14789_out0 : v$_14518_out0;
assign v$MUX8_3613_out0 = v$G2_15043_out0 ? v$FF2_14792_out0 : v$_14521_out0;
assign v$XOR3_4037_out0 = v$IR2$RD_16358_out0 ^ v$IR1$RM_18301_out0;
assign v$XOR3_4038_out0 = v$IR2$RD_16359_out0 ^ v$IR1$RM_18302_out0;
assign v$G20_5451_out0 = ! v$G19_16043_out0;
assign v$G20_5452_out0 = ! v$G19_16044_out0;
assign v$ShiftEN_5827_out0 = v$RXSHIFT_674_out0;
assign v$ShiftEN_5828_out0 = v$RXSHIFT_675_out0;
assign v$G6_5944_out0 = v$_9580_out0 && v$_8232_out0;
assign v$G6_5945_out0 = v$_9581_out0 && v$_8233_out0;
assign v$G9_6226_out0 = v$EQ2_7952_out0 || v$EQ3_15504_out0;
assign v$G9_6227_out0 = v$EQ2_7953_out0 || v$EQ3_15505_out0;
assign v$MUX2_6685_out0 = v$G47_1531_out0 ? v$C2_16240_out0 : v$G24_18388_out0;
assign v$MUX2_6686_out0 = v$G47_1532_out0 ? v$C2_16241_out0 : v$G24_18389_out0;
assign v$IR2$VALID_7421_out0 = v$IR2$VALID_18756_out0;
assign v$IR2$VALID_7422_out0 = v$IR2$VALID_18757_out0;
assign v$_7659_out0 = v$_12843_out0[0:0];
assign v$_7659_out1 = v$_12843_out0[1:1];
assign v$_7665_out0 = v$_12849_out0[0:0];
assign v$_7665_out1 = v$_12849_out0[1:1];
assign v$_7720_out0 = v$IR1_16680_out0[11:0];
assign v$_7721_out0 = v$IR1_16681_out0[11:0];
assign v$EQ9_7979_out0 = v$IR1_16680_out0 == 16'h7000;
assign v$EQ9_7980_out0 = v$IR1_16681_out0 == 16'h7000;
assign v$G19_8261_out0 = v$SHIFTEN_7092_out0 && v$CLK4_3694_out0;
assign v$G19_8262_out0 = v$SHIFTEN_7093_out0 && v$CLK4_3695_out0;
assign v$B_8316_out0 = v$B_3704_out0;
assign v$B_8317_out0 = v$B_3705_out0;
assign v$XOR1_8327_out0 = v$IR1$RM_18301_out0 ^ v$IR2$RD_16358_out0;
assign v$XOR1_8328_out0 = v$IR1$RM_18302_out0 ^ v$IR2$RD_16359_out0;
assign v$MUX1_8336_out0 = v$C_9609_out0 ? v$C1_14253_out0 : v$SHIFT_7019_out0;
assign v$MUX1_8337_out0 = v$C_9610_out0 ? v$C1_14254_out0 : v$SHIFT_7020_out0;
assign v$S_9424_out0 = v$S_8167_out0;
assign v$S_9425_out0 = v$S_8168_out0;
assign v$MUX5_9524_out0 = v$G2_15033_out0 ? v$FF5_1754_out0 : v$_7656_out1;
assign v$MUX5_9525_out0 = v$G2_15034_out0 ? v$FF5_1755_out0 : v$_7657_out1;
assign v$MUX5_9528_out0 = v$G2_15037_out0 ? v$FF5_1758_out0 : v$_7660_out1;
assign v$MUX5_9530_out0 = v$G2_15039_out0 ? v$FF5_1760_out0 : v$_7662_out1;
assign v$MUX5_9531_out0 = v$G2_15040_out0 ? v$FF5_1761_out0 : v$_7663_out1;
assign v$MUX5_9534_out0 = v$G2_15043_out0 ? v$FF5_1764_out0 : v$_7666_out1;
assign v$MUX3_9950_out0 = v$G2_15033_out0 ? v$FF7_8298_out0 : v$_14511_out1;
assign v$MUX3_9951_out0 = v$G2_15034_out0 ? v$FF7_8299_out0 : v$_14512_out1;
assign v$MUX3_9954_out0 = v$G2_15037_out0 ? v$FF7_8302_out0 : v$_14515_out1;
assign v$MUX3_9956_out0 = v$G2_15039_out0 ? v$FF7_8304_out0 : v$_14517_out1;
assign v$MUX3_9957_out0 = v$G2_15040_out0 ? v$FF7_8305_out0 : v$_14518_out1;
assign v$MUX3_9960_out0 = v$G2_15043_out0 ? v$FF7_8308_out0 : v$_14521_out1;
assign v$G3_10233_out0 = ! v$E_17351_out0;
assign v$G3_10234_out0 = ! v$E_17352_out0;
assign v$MUX6_10388_out0 = v$G2_15033_out0 ? v$FF1_16074_out0 : v$_1639_out1;
assign v$MUX6_10389_out0 = v$G2_15034_out0 ? v$FF1_16075_out0 : v$_1640_out1;
assign v$MUX6_10392_out0 = v$G2_15037_out0 ? v$FF1_16078_out0 : v$_1643_out1;
assign v$MUX6_10394_out0 = v$G2_15039_out0 ? v$FF1_16080_out0 : v$_1645_out1;
assign v$MUX6_10395_out0 = v$G2_15040_out0 ? v$FF1_16081_out0 : v$_1646_out1;
assign v$MUX6_10398_out0 = v$G2_15043_out0 ? v$FF1_16084_out0 : v$_1649_out1;
assign v$IR2$IS$FPU_11843_out0 = v$IR2$IS$FPU_2929_out0;
assign v$IR2$IS$FPU_11844_out0 = v$IR2$IS$FPU_2930_out0;
assign v$_11861_out0 = v$_8455_out1[0:0];
assign v$_11861_out1 = v$_8455_out1[1:1];
assign v$_11867_out0 = v$_8461_out1[0:0];
assign v$_11867_out1 = v$_8461_out1[1:1];
assign v$G32_11884_out0 = !(v$G30_18605_out0 || v$G23_4385_out0);
assign v$G32_11885_out0 = !(v$G30_18606_out0 || v$G23_4386_out0);
assign v$MUX5_11943_out0 = v$STP$SAVED_7560_out0 ? v$IR1_16680_out0 : v$R_18353_out0;
assign v$MUX5_11944_out0 = v$STP$SAVED_7561_out0 ? v$IR1_16681_out0 : v$R_18354_out0;
assign v$G4_11988_out0 = ! v$_2982_out0;
assign v$G4_11989_out0 = ! v$_2983_out0;
assign v$MUX2_12234_out0 = v$_10278_out0 ? v$FF1_10306_out0 : v$_13691_out0;
assign v$MUX2_12235_out0 = v$_10279_out0 ? v$FF1_10307_out0 : v$_13692_out0;
assign v$RXINT_12545_out0 = v$RXINTERRUPT_15347_out0;
assign v$RXINT_12546_out0 = v$RXINTERRUPT_15348_out0;
assign v$ISMOV_12630_out0 = v$ISMOV_6670_out0;
assign v$ISMOV_12631_out0 = v$ISMOV_6671_out0;
assign v$S_12819_out0 = v$S_8167_out0;
assign v$S_12820_out0 = v$S_8168_out0;
assign v$EQ2_12874_out0 = v$IR1$OPCODE_9564_out0 == 4'h1;
assign v$EQ2_12875_out0 = v$IR1$OPCODE_9565_out0 == 4'h1;
assign v$EQ1_12945_out0 = v$IR1$OPCODE_9564_out0 == 4'h0;
assign v$EQ1_12946_out0 = v$IR1$OPCODE_9565_out0 == 4'h0;
assign v$IR1_13389_out0 = v$IR1_16680_out0;
assign v$IR1_13390_out0 = v$IR1_16681_out0;
assign v$NEXTSTATE_13539_out0 = v$G2_7578_out0;
assign v$MUX2_13819_out0 = v$G2_15033_out0 ? v$FF8_14460_out0 : v$_11858_out1;
assign v$MUX2_13820_out0 = v$G2_15034_out0 ? v$FF8_14461_out0 : v$_11859_out1;
assign v$MUX2_13823_out0 = v$G2_15037_out0 ? v$FF8_14464_out0 : v$_11862_out1;
assign v$MUX2_13825_out0 = v$G2_15039_out0 ? v$FF8_14466_out0 : v$_11864_out1;
assign v$MUX2_13826_out0 = v$G2_15040_out0 ? v$FF8_14467_out0 : v$_11865_out1;
assign v$MUX2_13829_out0 = v$G2_15043_out0 ? v$FF8_14470_out0 : v$_11868_out1;
assign v$G36_14103_out0 = v$G37_18464_out0 && v$G38_10252_out0;
assign v$G36_14104_out0 = v$G37_18465_out0 && v$G38_10253_out0;
assign v$_14514_out0 = v$_8455_out0[0:0];
assign v$_14514_out1 = v$_8455_out0[1:1];
assign v$_14520_out0 = v$_8461_out0[0:0];
assign v$_14520_out1 = v$_8461_out0[1:1];
assign v$G68_15184_out0 = v$G69_8210_out0 || v$G70_10280_out0;
assign v$G68_15185_out0 = v$G69_8211_out0 || v$G70_10281_out0;
assign v$EQ6_15876_out0 = v$IR2$FPU$OP_2881_out0 == 2'h3;
assign v$EQ6_15877_out0 = v$IR2$FPU$OP_2882_out0 == 2'h3;
assign v$G9_16037_out0 = ! v$IR1$C$L_10053_out0;
assign v$G9_16038_out0 = ! v$IR1$C$L_10054_out0;
assign v$G10_16500_out0 = v$E_17351_out0 && v$NQ2_16698_out0;
assign v$G10_16501_out0 = v$E_17352_out0 && v$NQ2_16699_out0;
assign v$NR_16656_out0 = v$G12_16252_out0;
assign v$NR_16657_out0 = v$G12_16253_out0;
assign v$MUX4_16847_out0 = v$G2_15033_out0 ? v$FF6_2621_out0 : v$_11858_out0;
assign v$MUX4_16848_out0 = v$G2_15034_out0 ? v$FF6_2622_out0 : v$_11859_out0;
assign v$MUX4_16851_out0 = v$G2_15037_out0 ? v$FF6_2625_out0 : v$_11862_out0;
assign v$MUX4_16853_out0 = v$G2_15039_out0 ? v$FF6_2627_out0 : v$_11864_out0;
assign v$MUX4_16854_out0 = v$G2_15040_out0 ? v$FF6_2628_out0 : v$_11865_out0;
assign v$MUX4_16857_out0 = v$G2_15043_out0 ? v$FF6_2631_out0 : v$_11868_out0;
assign v$EQ15_17047_out0 = v$IR1$OPCODE_9564_out0 == 4'h1;
assign v$EQ15_17048_out0 = v$IR1$OPCODE_9565_out0 == 4'h1;
assign v$G2_17663_out0 = ! v$C_9609_out0;
assign v$G2_17664_out0 = ! v$C_9610_out0;
assign v$MUX1_17728_out0 = v$_2652_out0 ? v$C2_10009_out0 : v$C1_16322_out0;
assign v$MUX1_17729_out0 = v$_2653_out0 ? v$C2_10010_out0 : v$C1_16323_out0;
assign v$MUX7_17903_out0 = v$G2_15033_out0 ? v$FF3_9971_out0 : v$_1639_out0;
assign v$MUX7_17904_out0 = v$G2_15034_out0 ? v$FF3_9972_out0 : v$_1640_out0;
assign v$MUX7_17907_out0 = v$G2_15037_out0 ? v$FF3_9975_out0 : v$_1643_out0;
assign v$MUX7_17909_out0 = v$G2_15039_out0 ? v$FF3_9977_out0 : v$_1645_out0;
assign v$MUX7_17910_out0 = v$G2_15040_out0 ? v$FF3_9978_out0 : v$_1646_out0;
assign v$MUX7_17913_out0 = v$G2_15043_out0 ? v$FF3_9981_out0 : v$_1649_out0;
assign v$G11_18016_out0 = v$G10_2906_out0 && v$CheckParity_18678_out0;
assign v$G11_18017_out0 = v$G10_2907_out0 && v$CheckParity_18679_out0;
assign v$XOR2_18493_out0 = v$IR1$RD_5489_out0 ^ v$IR2$RD_16358_out0;
assign v$XOR2_18494_out0 = v$IR1$RD_5490_out0 ^ v$IR2$RD_16359_out0;
assign v$FINISHED_18669_out0 = v$FINISHED_7003_out0;
assign v$IR1_22_out0 = v$IR1_13389_out0;
assign v$IR1_23_out0 = v$IR1_13390_out0;
assign v$G29_681_out0 = ! v$EQ16_1582_out0;
assign v$G29_682_out0 = ! v$EQ16_1583_out0;
assign v$_893_out0 = v$B_8316_out0[2:2];
assign v$_894_out0 = v$B_8317_out0[2:2];
assign v$G34_1570_out0 = v$G35_4315_out0 || v$G36_14103_out0;
assign v$G34_1571_out0 = v$G35_4316_out0 || v$G36_14104_out0;
assign v$FINISHED_2255_out0 = v$FINISHED_18669_out0;
assign v$G8_2414_out0 = ! v$G9_6226_out0;
assign v$G8_2415_out0 = ! v$G9_6227_out0;
assign v$MUX1_2585_out0 = v$G2_15036_out0 ? v$SIN_94_out0 : v$_7659_out0;
assign v$MUX1_2591_out0 = v$G2_15042_out0 ? v$SIN_100_out0 : v$_7665_out0;
assign v$NE_3429_out0 = v$G3_10233_out0;
assign v$NE_3430_out0 = v$G3_10234_out0;
assign v$RXErrorSet_3480_out0 = v$G11_18016_out0;
assign v$RXErrorSet_3481_out0 = v$G11_18017_out0;
assign v$MUX8_3606_out0 = v$G2_15036_out0 ? v$FF2_14785_out0 : v$_14514_out0;
assign v$MUX8_3612_out0 = v$G2_15042_out0 ? v$FF2_14791_out0 : v$_14520_out0;
assign v$EQ6_3957_out0 = v$XOR2_18493_out0 == 2'h0;
assign v$EQ6_3958_out0 = v$XOR2_18494_out0 == 2'h0;
assign v$ISMOV_4078_out0 = v$ISMOV_12630_out0;
assign v$ISMOV_4079_out0 = v$ISMOV_12631_out0;
assign v$EQ5_4856_out0 = v$XOR3_4037_out0 == 2'h0;
assign v$EQ5_4857_out0 = v$XOR3_4038_out0 == 2'h0;
assign v$G1_5421_out0 = v$G10_16500_out0 && v$G11_8230_out0;
assign v$G1_5422_out0 = v$G10_16501_out0 && v$G11_8231_out0;
assign v$Q1P_5742_out0 = v$MUX2_6685_out0;
assign v$Q1P_5743_out0 = v$MUX2_6686_out0;
assign v$G21_7484_out0 = v$EQ6_15876_out0 && v$IR2$FPU$L_10744_out0;
assign v$G21_7485_out0 = v$EQ6_15877_out0 && v$IR2$FPU$L_10745_out0;
assign v$INTERRUPT1_8284_out0 = v$RXINT_12545_out0;
assign v$INTERRUPT1_8285_out0 = v$RXINT_12546_out0;
assign v$ISMOV_8767_out0 = v$ISMOV_12630_out0;
assign v$ISMOV_8768_out0 = v$ISMOV_12631_out0;
assign v$MUX5_9527_out0 = v$G2_15036_out0 ? v$FF5_1757_out0 : v$_7659_out1;
assign v$MUX5_9533_out0 = v$G2_15042_out0 ? v$FF5_1763_out0 : v$_7665_out1;
assign v$SR_9927_out0 = v$MUX1_8336_out0;
assign v$SR_9928_out0 = v$MUX1_8337_out0;
assign v$MUX3_9953_out0 = v$G2_15036_out0 ? v$FF7_8301_out0 : v$_14514_out1;
assign v$MUX3_9959_out0 = v$G2_15042_out0 ? v$FF7_8307_out0 : v$_14520_out1;
assign v$S_10347_out0 = v$S_12819_out0;
assign v$S_10348_out0 = v$S_12820_out0;
assign v$MUX6_10391_out0 = v$G2_15036_out0 ? v$FF1_16077_out0 : v$_1642_out1;
assign v$MUX6_10397_out0 = v$G2_15042_out0 ? v$FF1_16083_out0 : v$_1648_out1;
assign v$_10787_out0 = v$B_8316_out0[1:1];
assign v$_10788_out0 = v$B_8317_out0[1:1];
assign v$G67_11059_out0 = v$G71_15274_out0 && v$G68_15184_out0;
assign v$G67_11060_out0 = v$G71_15275_out0 && v$G68_15185_out0;
assign v$EQUAL_11623_out0 = v$G32_11884_out0;
assign v$EQUAL_11624_out0 = v$G32_11885_out0;
assign v$TX_11681_out0 = v$TX_1298_out0;
assign v$TX_11682_out0 = v$TX_1299_out0;
assign v$IR1$IS$LDST_13203_out0 = v$EQ1_12945_out0;
assign v$IR1$IS$LDST_13204_out0 = v$EQ1_12946_out0;
assign v$MUX2_13822_out0 = v$G2_15036_out0 ? v$FF8_14463_out0 : v$_11861_out1;
assign v$MUX2_13828_out0 = v$G2_15042_out0 ? v$FF8_14469_out0 : v$_11867_out1;
assign v$_14324_out0 = v$B_8316_out0[3:3];
assign v$_14325_out0 = v$B_8317_out0[3:3];
assign v$N_14507_out0 = v$_7720_out0;
assign v$N_14508_out0 = v$_7721_out0;
assign v$G10_14566_out0 = v$EQ2_12874_out0 && v$EQ4_5414_out0;
assign v$G10_14567_out0 = v$EQ2_12875_out0 && v$EQ4_5415_out0;
assign v$IR2$VALID_14823_out0 = v$IR2$VALID_7421_out0;
assign v$IR2$VALID_14824_out0 = v$IR2$VALID_7422_out0;
assign v$_15138_out0 = v$B_8316_out0[0:0];
assign v$_15139_out0 = v$B_8317_out0[0:0];
assign v$EQ3_15281_out0 = v$XOR1_8327_out0 == 2'h0;
assign v$EQ3_15282_out0 = v$XOR1_8328_out0 == 2'h0;
assign v$STP$DECODED_16534_out0 = v$EQ9_7979_out0;
assign v$STP$DECODED_16535_out0 = v$EQ9_7980_out0;
assign v$MUX4_16850_out0 = v$G2_15036_out0 ? v$FF6_2624_out0 : v$_11861_out0;
assign v$MUX4_16856_out0 = v$G2_15042_out0 ? v$FF6_2630_out0 : v$_11867_out0;
assign v$S_16937_out0 = v$RXset_1701_out0;
assign v$S_16948_out0 = v$RXset_1702_out0;
assign v$G16_16990_out0 = v$RXset_1701_out0 && v$RXlast_12821_out0;
assign v$G16_16991_out0 = v$RXset_1702_out0 && v$RXlast_12822_out0;
assign v$G9_17008_out0 = v$NQ2_2980_out0 && v$NR_16656_out0;
assign v$G9_17009_out0 = v$NQ2_2981_out0 && v$NR_16657_out0;
assign v$G3_17690_out0 = ! v$R_1586_out0;
assign v$OP_17803_out0 = v$_304_out0;
assign v$OP_17804_out0 = v$_305_out0;
assign v$MUX7_17906_out0 = v$G2_15036_out0 ? v$FF3_9974_out0 : v$_1642_out0;
assign v$MUX7_17912_out0 = v$G2_15042_out0 ? v$FF3_9980_out0 : v$_1648_out0;
assign v$S_17947_out0 = v$S_9424_out0;
assign v$S_17948_out0 = v$S_9425_out0;
assign v$G20_18281_out0 = v$NR_16656_out0 || v$Q3_18289_out0;
assign v$G20_18282_out0 = v$NR_16657_out0 || v$Q3_18290_out0;
assign v$G1_18647_out0 = v$ShiftEN_5827_out0 && v$CLK4_8834_out0;
assign v$G1_18648_out0 = v$ShiftEN_5828_out0 && v$CLK4_8835_out0;
assign v$G1_166_out0 = v$S_2443_out0 && v$ISMOV_8767_out0;
assign v$G1_167_out0 = v$S_2444_out0 && v$ISMOV_8768_out0;
assign v$G1_1249_out0 = v$S_901_out0 && v$ISMOV_4078_out0;
assign v$G1_1250_out0 = v$S_902_out0 && v$ISMOV_4079_out0;
assign v$G30_1717_out0 = v$EQ15_17047_out0 && v$G29_681_out0;
assign v$G30_1718_out0 = v$EQ15_17048_out0 && v$G29_682_out0;
assign v$G2_2425_out0 = v$EQUAL_11623_out0 && v$G3_10988_out0;
assign v$G2_2426_out0 = v$EQUAL_11624_out0 && v$G3_10989_out0;
assign v$G15_2677_out0 = v$IR1$IS$LDST_13203_out0 && v$IR1$S$WB_322_out0;
assign v$G15_2678_out0 = v$IR1$IS$LDST_13204_out0 && v$IR1$S$WB_323_out0;
assign v$IS$IR1$FMUL_2964_out0 = v$G10_14566_out0;
assign v$IS$IR1$FMUL_2965_out0 = v$G10_14567_out0;
assign v$G24_3401_out0 = v$IR1$IS$LDST_13203_out0 && v$IR1$S$WB_322_out0;
assign v$G24_3402_out0 = v$IR1$IS$LDST_13204_out0 && v$IR1$S$WB_323_out0;
assign v$SR_4368_out0 = v$SR_9927_out0;
assign v$SR_4369_out0 = v$SR_9927_out0;
assign v$SR_4370_out0 = v$SR_9927_out0;
assign v$SR_4371_out0 = v$SR_9927_out0;
assign v$SR_4372_out0 = v$SR_9928_out0;
assign v$SR_4373_out0 = v$SR_9928_out0;
assign v$SR_4374_out0 = v$SR_9928_out0;
assign v$SR_4375_out0 = v$SR_9928_out0;
assign v$OP_5038_out0 = v$OP_17803_out0;
assign v$OP_5039_out0 = v$OP_17804_out0;
assign v$G33_5131_out0 = v$NQ2_18563_out0 && v$G34_1570_out0;
assign v$G33_5132_out0 = v$NQ2_18564_out0 && v$G34_1571_out0;
assign v$IR2$VALID_6455_out0 = v$IR2$VALID_14823_out0;
assign v$IR2$VALID_6456_out0 = v$IR2$VALID_14824_out0;
assign v$G1_7325_out0 = v$G2_17663_out0 && v$_15138_out0;
assign v$G1_7326_out0 = v$G2_17664_out0 && v$_15139_out0;
assign v$IR1_7613_out0 = v$IR1_22_out0;
assign v$IR1_7614_out0 = v$IR1_23_out0;
assign v$G18_8420_out0 = v$G20_18281_out0 && v$G19_2412_out0;
assign v$G18_8421_out0 = v$G20_18282_out0 && v$G19_2413_out0;
assign v$G11_9603_out0 = v$EQ6_3957_out0 || v$EQ5_4856_out0;
assign v$G11_9604_out0 = v$EQ6_3958_out0 || v$EQ5_4857_out0;
assign v$Shift_9605_out0 = v$G1_18647_out0;
assign v$Shift_9606_out0 = v$G1_18648_out0;
assign v$EXEC2_9863_out0 = v$IR2$VALID_14823_out0;
assign v$EXEC2_9864_out0 = v$IR2$VALID_14824_out0;
assign v$IR2$VALID_10666_out0 = v$IR2$VALID_14823_out0;
assign v$IR2$VALID_10667_out0 = v$IR2$VALID_14824_out0;
assign v$G8_11068_out0 = v$Q1_10923_out0 && v$G9_17008_out0;
assign v$G8_11069_out0 = v$Q1_10924_out0 && v$G9_17009_out0;
assign v$FINISHED_11641_out0 = v$FINISHED_2255_out0;
assign v$G13_12160_out0 = v$G14_18435_out0 && v$NE_3429_out0;
assign v$G13_12161_out0 = v$G14_18436_out0 && v$NE_3430_out0;
assign v$ERR_12774_out0 = v$RXErrorSet_3480_out0;
assign v$ERR_12775_out0 = v$RXErrorSet_3481_out0;
assign v$G1_12982_out0 = v$STATE_16013_out0 && v$G3_17690_out0;
assign v$G15_13603_out0 = v$NE_3429_out0 && v$G16_3022_out0;
assign v$G15_13604_out0 = v$NE_3430_out0 && v$G16_3023_out0;
assign v$G32_14201_out0 = v$IR1$IS$LDST_13203_out0 && v$G34_4880_out0;
assign v$G32_14202_out0 = v$IR1$IS$LDST_13204_out0 && v$G34_4881_out0;
assign v$G25_14659_out0 = v$G21_7484_out0 && v$EQ7_3506_out0;
assign v$G25_14660_out0 = v$G21_7485_out0 && v$EQ7_3507_out0;
assign v$G4_14683_out0 = v$NE_3429_out0 && v$G5_10690_out0;
assign v$G4_14684_out0 = v$NE_3430_out0 && v$G5_10691_out0;
assign v$G17_14794_out0 = v$IR2$VALID_14823_out0 && v$G20_5451_out0;
assign v$G17_14795_out0 = v$IR2$VALID_14824_out0 && v$G20_5452_out0;
assign v$N_14843_out0 = v$N_14507_out0;
assign v$N_14844_out0 = v$N_14508_out0;
assign v$EQUAL_15828_out0 = v$EQUAL_11623_out0;
assign v$EQUAL_15829_out0 = v$EQUAL_11624_out0;
assign v$EXEC2_15883_out0 = v$IR2$VALID_14823_out0;
assign v$EXEC2_15884_out0 = v$IR2$VALID_14824_out0;
assign v$TXRST_16379_out0 = v$G67_11059_out0;
assign v$TXRST_16380_out0 = v$G67_11060_out0;
assign v$EN_16386_out0 = v$_10787_out0;
assign v$EN_16387_out0 = v$_893_out0;
assign v$EN_16388_out0 = v$_14324_out0;
assign v$EN_16390_out0 = v$_10788_out0;
assign v$EN_16391_out0 = v$_894_out0;
assign v$EN_16392_out0 = v$_14325_out0;
assign v$S_16939_out0 = v$G16_16990_out0;
assign v$S_16950_out0 = v$G16_16991_out0;
assign v$G14_17038_out0 = v$IR1$IS$LDST_13203_out0 && v$G9_16037_out0;
assign v$G14_17039_out0 = v$IR1$IS$LDST_13204_out0 && v$G9_16038_out0;
assign v$G36_17349_out0 = ! v$STP$DECODED_16534_out0;
assign v$G36_17350_out0 = ! v$STP$DECODED_16535_out0;
assign v$EDGE1_17407_out0 = v$INTERRUPT1_8284_out0;
assign v$EDGE1_17408_out0 = v$INTERRUPT1_8285_out0;
assign v$EXEC2_429_out0 = v$EXEC2_15883_out0;
assign v$EXEC2_430_out0 = v$EXEC2_15884_out0;
assign v$IR1$IS$FPU$ARITHMETIC_1370_out0 = v$G30_1717_out0;
assign v$IR1$IS$FPU$ARITHMETIC_1371_out0 = v$G30_1718_out0;
assign v$G1_1915_out0 = v$EXEC2_15883_out0 && v$IR15_10986_out0;
assign v$G1_1916_out0 = v$EXEC2_15884_out0 && v$IR15_10987_out0;
assign v$EXEC2_1945_out0 = v$EXEC2_9863_out0;
assign v$EXEC2_1946_out0 = v$EXEC2_9864_out0;
assign v$G12_2215_out0 = v$G13_12160_out0 || v$G15_13603_out0;
assign v$G12_2216_out0 = v$G13_12161_out0 || v$G15_13604_out0;
assign v$G3_2441_out0 = v$G15_2677_out0 && v$IS$IR2$DATA$PROCESSING_9944_out0;
assign v$G3_2442_out0 = v$G15_2678_out0 && v$IS$IR2$DATA$PROCESSING_9945_out0;
assign v$G29_3624_out0 = v$G30_2466_out0 || v$G33_5131_out0;
assign v$G29_3625_out0 = v$G30_2467_out0 || v$G33_5132_out0;
assign v$G3_3941_out0 = v$G8_11068_out0 || v$G10_18186_out0;
assign v$G3_3942_out0 = v$G8_11069_out0 || v$G10_18187_out0;
assign v$SEL1_5240_out0 = v$IR1_7613_out0[9:8];
assign v$SEL1_5241_out0 = v$IR1_7614_out0[9:8];
assign v$G12_6167_out0 = v$IS$IR1$FMUL_2964_out0 && v$G11_9603_out0;
assign v$G12_6168_out0 = v$IS$IR1$FMUL_2965_out0 && v$G11_9604_out0;
assign v$_6182_out0 = v$IR1_7613_out0[1:0];
assign v$_6183_out0 = v$IR1_7614_out0[1:0];
assign v$IR2$VALID$AND$NOT$FLOAD_7285_out0 = v$G17_14794_out0;
assign v$IR2$VALID$AND$NOT$FLOAD_7286_out0 = v$G17_14795_out0;
assign v$FINISHED_8010_out0 = v$FINISHED_11641_out0;
assign v$TXRST_8044_out0 = v$TXRST_16379_out0;
assign v$TXRST_8045_out0 = v$TXRST_16380_out0;
assign v$N_8269_out0 = v$N_14843_out0;
assign v$N_8270_out0 = v$N_14844_out0;
assign v$S_10442_out0 = v$G1_1249_out0;
assign v$S_10443_out0 = v$G1_1250_out0;
assign v$S_10699_out0 = v$G1_166_out0;
assign v$S_10700_out0 = v$G1_167_out0;
assign v$N_11963_out0 = v$N_14843_out0;
assign v$N_11964_out0 = v$N_14844_out0;
assign v$_12772_out0 = v$IR1_7613_out0[15:15];
assign v$_12773_out0 = v$IR1_7614_out0[15:15];
assign v$G26_13177_out0 = v$G24_3401_out0 && v$G25_2464_out0;
assign v$G26_13178_out0 = v$G24_3402_out0 && v$G25_2465_out0;
assign v$SEL13_13249_out0 = v$IR1_7613_out0[5:5];
assign v$IR2$VALID_13250_out0 = v$IR2$VALID_6455_out0;
assign v$IR2$VALID_13251_out0 = v$IR2$VALID_6456_out0;
assign v$_13542_out0 = v$IR1_7613_out0[8:8];
assign v$_13543_out0 = v$IR1_7614_out0[8:8];
assign v$G23_14080_out0 = ! v$G25_14659_out0;
assign v$G23_14081_out0 = ! v$G25_14660_out0;
assign v$G37_14088_out0 = v$IS$IR1$FMUL_2964_out0 && v$IS$IR2$DATA$PROCESSING_9944_out0;
assign v$G37_14089_out0 = v$IS$IR1$FMUL_2965_out0 && v$IS$IR2$DATA$PROCESSING_9945_out0;
assign v$SEL13_14655_out0 = v$IR1_7614_out0[5:5];
assign v$OP_14780_out0 = v$OP_5038_out0;
assign v$OP_14781_out0 = v$OP_5039_out0;
assign v$COUNTERINTERRUPT_14849_out0 = v$G2_2425_out0;
assign v$COUNTERINTERRUPT_14850_out0 = v$G2_2426_out0;
assign v$IR2$VALID_15878_out0 = v$IR2$VALID_10666_out0;
assign v$IR2$VALID_15879_out0 = v$IR2$VALID_10667_out0;
assign v$_15923_out0 = v$IR1_7613_out0[11:10];
assign v$_15924_out0 = v$IR1_7614_out0[11:10];
assign v$EN_16385_out0 = v$G1_7325_out0;
assign v$EN_16389_out0 = v$G1_7326_out0;
assign v$_16682_out0 = v$IR1_7613_out0[14:12];
assign v$_16683_out0 = v$IR1_7614_out0[14:12];
assign v$SR_16801_out0 = v$SR_4368_out0;
assign v$SR_16802_out0 = v$SR_4369_out0;
assign v$SR_16803_out0 = v$SR_4370_out0;
assign v$SR_16804_out0 = v$SR_4371_out0;
assign v$SR_16805_out0 = v$SR_4372_out0;
assign v$SR_16806_out0 = v$SR_4373_out0;
assign v$SR_16807_out0 = v$SR_4374_out0;
assign v$SR_16808_out0 = v$SR_4375_out0;
assign v$EN_16966_out0 = v$EN_16386_out0;
assign v$EN_16967_out0 = v$EN_16387_out0;
assign v$EN_16968_out0 = v$EN_16388_out0;
assign v$EN_16970_out0 = v$EN_16390_out0;
assign v$EN_16971_out0 = v$EN_16391_out0;
assign v$EN_16972_out0 = v$EN_16392_out0;
assign v$G16_16978_out0 = v$EQ3_15281_out0 && v$G32_14201_out0;
assign v$G16_16979_out0 = v$EQ3_15282_out0 && v$G32_14202_out0;
assign v$INTERRUPT1_17700_out0 = v$EDGE1_17407_out0;
assign v$INTERRUPT1_17701_out0 = v$EDGE1_17408_out0;
assign v$G15_17828_out0 = v$G17_11683_out0 || v$G18_8420_out0;
assign v$G15_17829_out0 = v$G17_11684_out0 || v$G18_8421_out0;
assign v$IR1_18034_out0 = v$IR1_7613_out0;
assign v$IR1_18035_out0 = v$IR1_7614_out0;
assign v$IR1_646_out0 = v$IR1_18034_out0;
assign v$IR1_647_out0 = v$IR1_18035_out0;
assign v$R_1488_out0 = v$FINISHED_8010_out0;
assign v$G31_1822_out0 = v$G28_14668_out0 && v$IR1$IS$FPU$ARITHMETIC_1370_out0;
assign v$G31_1823_out0 = v$G28_14669_out0 && v$IR1$IS$FPU$ARITHMETIC_1371_out0;
assign v$SEL2_2434_out0 = v$IR1_18034_out0[15:12];
assign v$SEL2_2435_out0 = v$IR1_18035_out0[15:12];
assign v$EQ1_2818_out0 = v$SR_16802_out0 == 2'h1;
assign v$EQ1_2819_out0 = v$SR_16806_out0 == 2'h1;
assign v$EQ2_3209_out0 = v$SR_16804_out0 == 2'h2;
assign v$EQ2_3210_out0 = v$SR_16808_out0 == 2'h2;
assign v$G18_3399_out0 = v$INTERRUPT1_17700_out0 && v$G17_5476_out0;
assign v$G18_3400_out0 = v$INTERRUPT1_17701_out0 && v$G17_5477_out0;
assign v$TXINTERRUPT_3634_out0 = v$TXRST_8044_out0;
assign v$TXINTERRUPT_3635_out0 = v$TXRST_8045_out0;
assign v$IR1$FPU$OP_3837_out0 = v$SEL1_5240_out0;
assign v$IR1$FPU$OP_3838_out0 = v$SEL1_5241_out0;
assign v$IR1$D_4219_out0 = v$_15923_out0;
assign v$IR1$D_4220_out0 = v$_15924_out0;
assign v$G2_5047_out0 = v$Q3_18289_out0 && v$G3_3941_out0;
assign v$G2_5048_out0 = v$Q3_18290_out0 && v$G3_3942_out0;
assign v$EQ1_5072_out0 = v$SR_16803_out0 == 2'h1;
assign v$EQ1_5073_out0 = v$SR_16807_out0 == 2'h1;
assign v$EQ1_5080_out0 = v$SR_16801_out0 == 2'h3;
assign v$EQ1_5081_out0 = v$SR_16805_out0 == 2'h3;
assign v$G26_5127_out0 = v$G25_10273_out0 || v$FINISHED_8010_out0;
assign v$G14_5384_out0 = v$G16_6407_out0 || v$G15_17828_out0;
assign v$G14_5385_out0 = v$G16_6408_out0 || v$G15_17829_out0;
assign v$EQ3_5436_out0 = v$SR_16803_out0 == 2'h3;
assign v$EQ3_5437_out0 = v$SR_16807_out0 == 2'h3;
assign v$IR1$32$BITS_5454_out0 = v$SEL13_14655_out0;
assign v$IR1$OP_5519_out0 = v$_16682_out0;
assign v$IR1$OP_5520_out0 = v$_16683_out0;
assign v$IR1$15_5758_out0 = v$_12772_out0;
assign v$IR1$15_5759_out0 = v$_12773_out0;
assign v$MUX3_6131_out0 = v$G47_1531_out0 ? v$C3_18552_out0 : v$G29_3624_out0;
assign v$MUX3_6132_out0 = v$G47_1532_out0 ? v$C3_18553_out0 : v$G29_3625_out0;
assign v$G4_7548_out0 = v$G3_2441_out0 || v$G16_16978_out0;
assign v$G4_7549_out0 = v$G3_2442_out0 || v$G16_16979_out0;
assign v$IR1$S_7842_out0 = v$_13542_out0;
assign v$IR1$S_7843_out0 = v$_13543_out0;
assign v$IR1$32$BITS_7867_out0 = v$SEL13_13249_out0;
assign v$EQ3_7898_out0 = v$SR_16801_out0 == 2'h1;
assign v$EQ3_7899_out0 = v$SR_16805_out0 == 2'h1;
assign v$EQ1_10409_out0 = v$SR_16804_out0 == 2'h3;
assign v$EQ1_10410_out0 = v$SR_16808_out0 == 2'h3;
assign v$OP_10992_out0 = v$OP_14780_out0;
assign v$OP_10993_out0 = v$OP_14781_out0;
assign v$_11757_out0 = { v$N_11963_out0,v$C1_5412_out0 };
assign v$_11758_out0 = { v$N_11964_out0,v$C1_5413_out0 };
assign v$G6_11934_out0 = v$IR2$VALID_13250_out0 && v$IR2$L_12464_out0;
assign v$G6_11935_out0 = v$IR2$VALID_13251_out0 && v$IR2$L_12465_out0;
assign v$EQ3_12136_out0 = v$SR_16804_out0 == 2'h1;
assign v$EQ3_12137_out0 = v$SR_16808_out0 == 2'h1;
assign v$IR1$M_13247_out0 = v$_6182_out0;
assign v$IR1$M_13248_out0 = v$_6183_out0;
assign v$G7_13559_out0 = v$G1_1915_out0 && v$G8_2414_out0;
assign v$G7_13560_out0 = v$G1_1916_out0 && v$G8_2415_out0;
assign v$EQ2_13623_out0 = v$SR_16802_out0 == 2'h2;
assign v$EQ2_13624_out0 = v$SR_16806_out0 == 2'h2;
assign v$EQ2_14300_out0 = v$SR_16801_out0 == 2'h2;
assign v$EQ2_14301_out0 = v$SR_16805_out0 == 2'h2;
assign v$FMUL$FINISHED_14472_out0 = v$FINISHED_8010_out0;
assign v$G14_14681_out0 = ! v$INTERRUPT1_17700_out0;
assign v$G14_14682_out0 = ! v$INTERRUPT1_17701_out0;
assign v$EXEC2_16363_out0 = v$EXEC2_1945_out0;
assign v$EXEC2_16364_out0 = v$EXEC2_1946_out0;
assign v$EQ2_16393_out0 = v$SR_16803_out0 == 2'h2;
assign v$EQ2_16394_out0 = v$SR_16807_out0 == 2'h2;
assign v$G32_16412_out0 = v$INTERRUPT3_3508_out0 || v$COUNTERINTERRUPT_14849_out0;
assign v$G32_16413_out0 = v$INTERRUPT3_3509_out0 || v$COUNTERINTERRUPT_14850_out0;
assign v$EQ3_16544_out0 = v$SR_16802_out0 == 2'h3;
assign v$EQ3_16545_out0 = v$SR_16806_out0 == 2'h3;
assign v$EN_16965_out0 = v$EN_16385_out0;
assign v$EN_16969_out0 = v$EN_16389_out0;
assign v$TXReset_17834_out0 = v$TXRST_8044_out0;
assign v$TXReset_17835_out0 = v$TXRST_8045_out0;
assign v$G24_17931_out0 = v$IR2$VALID_13250_out0 && v$G23_14080_out0;
assign v$G24_17932_out0 = v$IR2$VALID_13251_out0 && v$G23_14081_out0;
assign v$N_18295_out0 = v$N_8269_out0;
assign v$N_18296_out0 = v$N_8270_out0;
assign v$G21_18680_out0 = v$IR2$VALID$AND$NOT$FLOAD_7285_out0 && v$EQ11_11882_out0;
assign v$G21_18681_out0 = v$IR2$VALID$AND$NOT$FLOAD_7286_out0 && v$EQ11_11883_out0;
assign v$R_1587_out0 = v$R_1488_out0;
assign v$N_1621_out0 = v$N_18295_out0;
assign v$N_1622_out0 = v$N_18296_out0;
assign v$G8_1886_out0 = v$EQ1_5080_out0 && v$EN_16965_out0;
assign v$G8_1887_out0 = v$EQ3_16544_out0 && v$EN_16966_out0;
assign v$G8_1888_out0 = v$EQ3_5436_out0 && v$EN_16967_out0;
assign v$G8_1889_out0 = v$EQ1_10409_out0 && v$EN_16968_out0;
assign v$G8_1890_out0 = v$EQ1_5081_out0 && v$EN_16969_out0;
assign v$G8_1891_out0 = v$EQ3_16545_out0 && v$EN_16970_out0;
assign v$G8_1892_out0 = v$EQ3_5437_out0 && v$EN_16971_out0;
assign v$G8_1893_out0 = v$EQ1_10410_out0 && v$EN_16972_out0;
assign v$NEXTENDED_1909_out0 = v$_11757_out0;
assign v$NEXTENDED_1910_out0 = v$_11758_out0;
assign v$G3_2605_out0 = v$EQ3_7898_out0 && v$EN_16965_out0;
assign v$G3_2606_out0 = v$EQ1_2818_out0 && v$EN_16966_out0;
assign v$G3_2607_out0 = v$EQ1_5072_out0 && v$EN_16967_out0;
assign v$G3_2608_out0 = v$EQ3_12136_out0 && v$EN_16968_out0;
assign v$G3_2609_out0 = v$EQ3_7899_out0 && v$EN_16969_out0;
assign v$G3_2610_out0 = v$EQ1_2819_out0 && v$EN_16970_out0;
assign v$G3_2611_out0 = v$EQ1_5073_out0 && v$EN_16971_out0;
assign v$G3_2612_out0 = v$EQ3_12137_out0 && v$EN_16972_out0;
assign v$MUX2_2884_out0 = v$IR2$VALID$AND$NOT$FLOAD_7285_out0 ? v$IR2$D_14491_out0 : v$IR1$M_13247_out0;
assign v$MUX2_2885_out0 = v$IR2$VALID$AND$NOT$FLOAD_7286_out0 ? v$IR2$D_14492_out0 : v$IR1$M_13248_out0;
assign v$OP_3690_out0 = v$OP_10992_out0;
assign v$OP_3691_out0 = v$OP_10993_out0;
assign v$EXEC2_3998_out0 = v$EXEC2_16363_out0;
assign v$EXEC2_3999_out0 = v$EXEC2_16364_out0;
assign v$G4_4029_out0 = v$EQ2_14300_out0 && v$EN_16965_out0;
assign v$G4_4030_out0 = v$EQ2_13623_out0 && v$EN_16966_out0;
assign v$G4_4031_out0 = v$EQ2_16393_out0 && v$EN_16967_out0;
assign v$G4_4032_out0 = v$EQ2_3209_out0 && v$EN_16968_out0;
assign v$G4_4033_out0 = v$EQ2_14301_out0 && v$EN_16969_out0;
assign v$G4_4034_out0 = v$EQ2_13624_out0 && v$EN_16970_out0;
assign v$G4_4035_out0 = v$EQ2_16394_out0 && v$EN_16971_out0;
assign v$G4_4036_out0 = v$EQ2_3210_out0 && v$EN_16972_out0;
assign v$EXEC2_4387_out0 = v$EXEC2_16363_out0;
assign v$EXEC2_4388_out0 = v$EXEC2_16364_out0;
assign v$G16_4469_out0 = v$FF2_16652_out0 && v$G14_14681_out0;
assign v$G16_4470_out0 = v$FF2_16653_out0 && v$G14_14682_out0;
assign v$TXINT_4911_out0 = v$TXINTERRUPT_3634_out0;
assign v$TXINT_4912_out0 = v$TXINTERRUPT_3635_out0;
assign v$Q2P_6039_out0 = v$MUX3_6131_out0;
assign v$Q2P_6040_out0 = v$MUX3_6132_out0;
assign v$G8_6064_out0 = v$G4_7548_out0 || v$G14_17038_out0;
assign v$G8_6065_out0 = v$G4_7549_out0 || v$G14_17039_out0;
assign v$EQ3_7234_out0 = v$IR1$FPU$OP_3837_out0 == 2'h2;
assign v$EQ3_7235_out0 = v$IR1$FPU$OP_3838_out0 == 2'h2;
assign v$EXEC2_8015_out0 = v$EXEC2_16363_out0;
assign v$EXEC2_8016_out0 = v$EXEC2_16364_out0;
assign v$G36_8050_out0 = v$G31_1822_out0 || v$G37_14088_out0;
assign v$G36_8051_out0 = v$G31_1823_out0 || v$G37_14089_out0;
assign v$EQ16_10749_out0 = v$IR1$FPU$OP_3837_out0 == 2'h3;
assign v$32BIT_10933_out0 = v$IR1$32$BITS_5454_out0;
assign v$RD_11793_out0 = v$IR1$D_4219_out0;
assign v$S_12649_out0 = v$IR1$S_7842_out0;
assign v$S_12650_out0 = v$IR1$S_7843_out0;
assign v$G15_13391_out0 = v$G18_3399_out0 && v$R1_15011_out0;
assign v$G15_13392_out0 = v$G18_3400_out0 && v$R1_15012_out0;
assign v$FINISHED_13867_out0 = v$FMUL$FINISHED_14472_out0;
assign v$INT3_14034_out0 = v$G32_16412_out0;
assign v$INT3_14035_out0 = v$G32_16413_out0;
assign v$G13_15105_out0 = v$NQ0_7796_out0 && v$G14_5384_out0;
assign v$G13_15106_out0 = v$NQ0_7797_out0 && v$G14_5385_out0;
assign v$G4_15824_out0 = ! v$IR1$15_5758_out0;
assign v$G4_15825_out0 = ! v$IR1$15_5759_out0;
assign v$IR1_15998_out0 = v$IR1_646_out0;
assign v$IR1_15999_out0 = v$IR1_647_out0;
assign v$EQ4_16505_out0 = v$IR1$FPU$OP_3837_out0 == 2'h2;
assign v$EQ4_16506_out0 = v$IR1$FPU$OP_3838_out0 == 2'h2;
assign v$IR1$FULL$OP$CODE_17055_out0 = v$SEL2_2434_out0;
assign v$IR1$FULL$OP$CODE_17056_out0 = v$SEL2_2435_out0;
assign v$EXEC2_17638_out0 = v$EXEC2_16363_out0;
assign v$EXEC2_17639_out0 = v$EXEC2_16364_out0;
assign v$N_17937_out0 = v$N_18295_out0;
assign v$N_17938_out0 = v$N_18296_out0;
assign v$R_18337_out0 = v$TXReset_17834_out0;
assign v$R_18348_out0 = v$TXReset_17835_out0;
assign v$WENALU_18660_out0 = v$G7_13559_out0;
assign v$WENALU_18661_out0 = v$G7_13560_out0;
assign v$_41_out0 = v$IR1_15998_out0[8:8];
assign v$_42_out0 = v$IR1_15999_out0[8:8];
assign v$FMUL$FINISHED_200_out0 = v$FINISHED_13867_out0;
assign v$EQ8_252_out0 = v$IR1$FULL$OP$CODE_17055_out0 == 4'h0;
assign v$EQ8_253_out0 = v$IR1$FULL$OP$CODE_17056_out0 == 4'h0;
assign v$_909_out0 = v$IR1_15998_out0[11:10];
assign v$_910_out0 = v$IR1_15999_out0[11:10];
assign v$EXEC2_1167_out0 = v$EXEC2_4387_out0;
assign v$EXEC2_1168_out0 = v$EXEC2_4388_out0;
assign v$EXEC2_1469_out0 = v$EXEC2_8015_out0;
assign v$EXEC2_1470_out0 = v$EXEC2_8016_out0;
assign v$EQ5_1503_out0 = v$IR1$FULL$OP$CODE_17055_out0 == 4'h1;
assign v$EQ5_1504_out0 = v$IR1$FULL$OP$CODE_17056_out0 == 4'h1;
assign v$INTERRUPT0_1805_out0 = v$TXINT_4911_out0;
assign v$INTERRUPT0_1806_out0 = v$TXINT_4912_out0;
assign v$_1838_out0 = v$IR1_15998_out0[5:2];
assign v$_1839_out0 = v$IR1_15999_out0[5:2];
assign v$EQ5_1911_out0 = v$OP_3690_out0 == 4'h6;
assign v$EQ5_1912_out0 = v$OP_3691_out0 == 4'h6;
assign v$_1966_out0 = v$IR1_15998_out0[6:6];
assign v$_1967_out0 = v$IR1_15999_out0[6:6];
assign v$EDGE3_2241_out0 = v$INT3_14034_out0;
assign v$EDGE3_2242_out0 = v$INT3_14035_out0;
assign v$_2447_out0 = v$IR1_15998_out0[9:9];
assign v$_2448_out0 = v$IR1_15999_out0[9:9];
assign v$_2669_out0 = { v$Q2P_6039_out0,v$Q3P_11672_out0 };
assign v$_2670_out0 = { v$Q2P_6040_out0,v$Q3P_11673_out0 };
assign v$WENALU_4072_out0 = v$WENALU_18660_out0;
assign v$WENALU_4073_out0 = v$WENALU_18661_out0;
assign v$EQ1_4110_out0 = v$OP_3690_out0 == 4'h2;
assign v$EQ1_4111_out0 = v$OP_3691_out0 == 4'h2;
assign v$EQ3_5731_out0 = v$OP_3690_out0 == 4'h4;
assign v$EQ3_5732_out0 = v$OP_3691_out0 == 4'h4;
assign v$_7289_out0 = v$IR1_15998_out0[7:7];
assign v$_7290_out0 = v$IR1_15999_out0[7:7];
assign v$EXEC2_8048_out0 = v$EXEC2_17638_out0;
assign v$EXEC2_8049_out0 = v$EXEC2_17639_out0;
assign v$MUX16_8689_out0 = v$FINISHED_13867_out0 ? v$RD$FPU_12947_out0 : v$MUX2_2884_out0;
assign v$EQ13_9341_out0 = v$IR1$FULL$OP$CODE_17055_out0 == 4'h1;
assign v$EQ13_9342_out0 = v$IR1$FULL$OP$CODE_17056_out0 == 4'h1;
assign v$EQ4_9358_out0 = v$OP_3690_out0 == 4'h5;
assign v$EQ4_9359_out0 = v$OP_3691_out0 == 4'h5;
assign v$EXEC2_9439_out0 = v$EXEC2_3998_out0;
assign v$EXEC2_9440_out0 = v$EXEC2_3999_out0;
assign v$_10791_out0 = v$IR1_15998_out0[1:0];
assign v$_10792_out0 = v$IR1_15999_out0[1:0];
assign v$EQ2_10797_out0 = v$OP_3690_out0 == 4'h3;
assign v$EQ2_10798_out0 = v$OP_3691_out0 == 4'h3;
assign v$N_11753_out0 = v$N_17937_out0;
assign v$N_11754_out0 = v$N_17938_out0;
assign v$EQ14_12122_out0 = v$IR1$FULL$OP$CODE_17055_out0 == 4'h1;
assign v$EQ14_12123_out0 = v$IR1$FULL$OP$CODE_17056_out0 == 4'h1;
assign v$_12764_out0 = v$IR1_15998_out0[15:15];
assign v$_12765_out0 = v$IR1_15999_out0[15:15];
assign v$NEXTENDED_14372_out0 = v$NEXTENDED_1909_out0;
assign v$NEXTENDED_14373_out0 = v$NEXTENDED_1910_out0;
assign v$G13_14852_out0 = v$G8_6064_out0 || v$G12_6167_out0;
assign v$G13_14853_out0 = v$G8_6065_out0 || v$G12_6168_out0;
assign v$AD3_15145_out0 = v$MUX2_2885_out0;
assign v$G1_15293_out0 = v$G2_5047_out0 || v$G13_15105_out0;
assign v$G1_15294_out0 = v$G2_5048_out0 || v$G13_15106_out0;
assign v$G6_15565_out0 = ! v$R_18337_out0;
assign v$G6_15576_out0 = ! v$R_18348_out0;
assign v$EQ15_15790_out0 = v$IR1$FULL$OP$CODE_17055_out0 == 4'h1;
assign v$EQ2_15802_out0 = v$IR1_15998_out0 == 16'h7000;
assign v$EQ2_15803_out0 = v$IR1_15999_out0 == 16'h7000;
assign v$32BIT_15873_out0 = v$32BIT_10933_out0;
assign v$_16041_out0 = v$IR1_15998_out0[15:12];
assign v$_16042_out0 = v$IR1_15999_out0[15:12];
assign v$EQ6_16250_out0 = v$OP_3690_out0 == 4'h7;
assign v$EQ6_16251_out0 = v$OP_3691_out0 == 4'h7;
assign v$S_16383_out0 = v$S_12649_out0;
assign v$S_16384_out0 = v$S_12650_out0;
assign v$G13_16532_out0 = v$G16_4469_out0 && v$F1_3488_out0;
assign v$G13_16533_out0 = v$G16_4470_out0 && v$F1_3489_out0;
assign v$END_16598_out0 = v$N_1621_out0;
assign v$END_16599_out0 = v$N_1622_out0;
assign v$G3_17691_out0 = ! v$R_1587_out0;
assign v$JMI_73_out0 = v$EQ4_9358_out0;
assign v$JMI_74_out0 = v$EQ4_9359_out0;
assign v$G5_1123_out0 = v$FF2_13045_out0 && v$G6_15565_out0;
assign v$G5_1128_out0 = v$FF2_13056_out0 && v$G6_15576_out0;
assign v$JMP_1667_out0 = v$EQ3_5731_out0;
assign v$JMP_1668_out0 = v$EQ3_5732_out0;
assign v$JLS_1955_out0 = v$EQ2_10797_out0;
assign v$JLS_1956_out0 = v$EQ2_10798_out0;
assign v$G15_2283_out0 = v$32BIT_15873_out0 && v$IR2$IS$FPU_11844_out0;
assign v$INTERRUPT3_2816_out0 = v$EDGE3_2241_out0;
assign v$INTERRUPT3_2817_out0 = v$EDGE3_2242_out0;
assign v$IR1$OPCODE_2895_out0 = v$_16041_out0;
assign v$IR1$OPCODE_2896_out0 = v$_16042_out0;
assign v$INT2_3161_out0 = v$FMUL$FINISHED_200_out0;
assign v$G25_3549_out0 = ! v$EQ14_12122_out0;
assign v$G25_3550_out0 = ! v$EQ14_12123_out0;
assign v$IR1$P_3692_out0 = v$_7289_out0;
assign v$IR1$P_3693_out0 = v$_7290_out0;
assign v$IR1$L_5138_out0 = v$_2447_out0;
assign v$IR1$L_5139_out0 = v$_2448_out0;
assign v$EDGE0_5740_out0 = v$INTERRUPT0_1805_out0;
assign v$EDGE0_5741_out0 = v$INTERRUPT0_1806_out0;
assign v$STP_6205_out0 = v$EQ6_16250_out0;
assign v$STP_6206_out0 = v$EQ6_16251_out0;
assign v$STOP$1_7810_out0 = v$EQ2_15802_out0;
assign v$STOP$1_7811_out0 = v$EQ2_15803_out0;
assign v$IS$32$BIT_11006_out0 = v$32BIT_15873_out0;
assign v$Q0P_12171_out0 = v$G1_15293_out0;
assign v$Q0P_12172_out0 = v$G1_15294_out0;
assign v$IR1$M_12632_out0 = v$_10791_out0;
assign v$IR1$M_12633_out0 = v$_10792_out0;
assign v$G1_12983_out0 = v$STATE_16014_out0 && v$G3_17691_out0;
assign v$AD3_13144_out0 = v$AD3_15145_out0;
assign v$EQ10_13408_out0 = v$N_11753_out0 == 12'h2;
assign v$EQ10_13409_out0 = v$N_11754_out0 == 12'h2;
assign v$EQ11_13605_out0 = v$N_11753_out0 == 12'h4;
assign v$EQ11_13606_out0 = v$N_11754_out0 == 12'h4;
assign v$G28_13787_out0 = v$EQ16_10749_out0 && v$EQ15_15790_out0;
assign v$IS$32$BITS_14039_out0 = v$32BIT_15873_out0;
assign v$EQ8_14328_out0 = v$N_11753_out0 == 12'h0;
assign v$EQ8_14329_out0 = v$N_11754_out0 == 12'h0;
assign v$IR1$U_14776_out0 = v$_1966_out0;
assign v$IR1$U_14777_out0 = v$_1967_out0;
assign v$IR1$D_14847_out0 = v$_909_out0;
assign v$IR1$D_14848_out0 = v$_910_out0;
assign v$JLO_14983_out0 = v$EQ1_4110_out0;
assign v$JLO_14984_out0 = v$EQ1_4111_out0;
assign v$AD3_15144_out0 = v$MUX16_8689_out0;
assign v$G22_15631_out0 = v$EQ4_16505_out0 && v$EQ13_9341_out0;
assign v$G22_15632_out0 = v$EQ4_16506_out0 && v$EQ13_9342_out0;
assign v$IR1$N_15765_out0 = v$_1838_out0;
assign v$IR1$N_15766_out0 = v$_1839_out0;
assign v$IR1$LS_16424_out0 = v$_12764_out0;
assign v$IR1$LS_16425_out0 = v$_12765_out0;
assign v$IR1$W_16548_out0 = v$_41_out0;
assign v$IR1$W_16549_out0 = v$_42_out0;
assign v$G5_16556_out0 = v$EQ3_7234_out0 && v$EQ5_1503_out0;
assign v$G5_16557_out0 = v$EQ3_7235_out0 && v$EQ5_1504_out0;
assign v$G19_16696_out0 = v$G15_13391_out0 || v$G13_16532_out0;
assign v$G19_16697_out0 = v$G15_13392_out0 || v$G13_16533_out0;
assign v$G23_16770_out0 = v$G13_14852_out0 || v$G26_13177_out0;
assign v$G23_16771_out0 = v$G13_14853_out0 || v$G26_13178_out0;
assign v$EQ7_16898_out0 = v$N_11753_out0 == 12'h1;
assign v$EQ7_16899_out0 = v$N_11754_out0 == 12'h1;
assign v$G2_17064_out0 = v$S_16383_out0 && v$EXEC2_429_out0;
assign v$G2_17065_out0 = v$S_16384_out0 && v$EXEC2_430_out0;
assign v$EQ9_17768_out0 = v$N_11753_out0 == 12'h3;
assign v$EQ9_17769_out0 = v$N_11754_out0 == 12'h3;
assign v$JEQ_18036_out0 = v$EQ5_1911_out0;
assign v$JEQ_18037_out0 = v$EQ5_1912_out0;
assign v$EQ13_18548_out0 = v$N_11753_out0 == 12'h5;
assign v$EQ13_18549_out0 = v$N_11754_out0 == 12'h5;
assign v$IS$32$BITS_1282_out0 = v$IS$32$BITS_14039_out0;
assign v$JEQ_1675_out0 = v$JEQ_18036_out0;
assign v$JEQ_1676_out0 = v$JEQ_18037_out0;
assign v$G32_1826_out0 = v$INTERRUPT3_2816_out0 && v$G31_9632_out0;
assign v$G32_1827_out0 = v$INTERRUPT3_2817_out0 && v$G31_9633_out0;
assign v$G3_2671_out0 = v$G2_17064_out0 && v$G4_11988_out0;
assign v$G3_2672_out0 = v$G2_17065_out0 && v$G4_11989_out0;
assign v$G28_3167_out0 = ! v$INTERRUPT3_2816_out0;
assign v$G28_3168_out0 = ! v$INTERRUPT3_2817_out0;
assign v$INTERRUPT2_3853_out0 = v$INT2_3161_out0;
assign v$JMP_4337_out0 = v$JMP_1667_out0;
assign v$JMP_4338_out0 = v$JMP_1668_out0;
assign v$_5082_out0 = { v$Q0P_12171_out0,v$Q1P_11007_out0 };
assign v$_5083_out0 = { v$Q0P_12172_out0,v$Q1P_11008_out0 };
assign v$JLO_8109_out0 = v$JLO_14983_out0;
assign v$JLO_8110_out0 = v$JLO_14984_out0;
assign v$IR1$IS$FPU$LOAD$STORE_8930_out0 = v$G28_13787_out0;
assign v$IS$32$BIT_10863_out0 = v$IS$32$BIT_11006_out0;
assign v$_11646_out0 = { v$IR1$N_15765_out0,v$C4_15906_out0 };
assign v$_11647_out0 = { v$IR1$N_15766_out0,v$C4_15907_out0 };
assign v$INTERRUPT0_11700_out0 = v$EDGE0_5740_out0;
assign v$INTERRUPT0_11701_out0 = v$EDGE0_5741_out0;
assign v$STP_11714_out0 = v$STP_6205_out0;
assign v$STP_11715_out0 = v$STP_6206_out0;
assign v$G16_11965_out0 = ! v$IR1$W_16548_out0;
assign v$G16_11966_out0 = ! v$IR1$W_16549_out0;
assign v$AD3_13143_out0 = v$AD3_15144_out0;
assign v$JMI_13149_out0 = v$JMI_73_out0;
assign v$JMI_13150_out0 = v$JMI_74_out0;
assign v$G24_13860_out0 = v$G25_3549_out0 && v$G4_15824_out0;
assign v$G24_13861_out0 = v$G25_3550_out0 && v$G4_15825_out0;
assign v$EQ5_14374_out0 = v$IR1$OPCODE_2895_out0 == 4'h0;
assign v$EQ5_14375_out0 = v$IR1$OPCODE_2896_out0 == 4'h0;
assign v$G10_14893_out0 = ! v$STOP$1_7810_out0;
assign v$G10_14894_out0 = ! v$STOP$1_7811_out0;
assign v$EDGE1_15272_out0 = v$G19_16696_out0;
assign v$EDGE1_15273_out0 = v$G19_16697_out0;
assign v$IS$IR1$FMUL_15296_out0 = v$G22_15631_out0;
assign v$IS$IR1$FMUL_15297_out0 = v$G22_15632_out0;
assign v$JLS_16442_out0 = v$JLS_1955_out0;
assign v$JLS_16443_out0 = v$JLS_1956_out0;
assign v$G27_16528_out0 = v$G23_16770_out0 || v$G36_8050_out0;
assign v$G27_16529_out0 = v$G23_16771_out0 || v$G36_8051_out0;
assign v$EQ3_17921_out0 = v$IR1$OPCODE_2895_out0 == 4'h0;
assign v$EQ3_17922_out0 = v$IR1$OPCODE_2896_out0 == 4'h0;
assign v$G2_18429_out0 = ! v$IR1$L_5138_out0;
assign v$G2_18430_out0 = ! v$IR1$L_5139_out0;
assign v$G8_18779_out0 = ! v$IR1$U_14776_out0;
assign v$G8_18780_out0 = ! v$IR1$U_14777_out0;
assign v$_1231_out0 = { v$_5082_out0,v$_13065_out0 };
assign v$_1232_out0 = { v$_5083_out0,v$_13066_out0 };
assign v$DIN_1723_out0 = v$_11646_out0;
assign v$DIN_1724_out0 = v$_11647_out0;
assign v$G27_3882_out0 = ! v$IR1$IS$FPU$LOAD$STORE_8930_out0;
assign v$MUX11_4488_out0 = v$IS$IR1$FMUL_15297_out0 ? v$IR1$FPU$OP_3838_out0 : v$IR2$FPU$OP_1688_out0;
assign v$G17_5460_out0 = v$JLO_8109_out0 && v$G18_13513_out0;
assign v$G17_5461_out0 = v$JLO_8110_out0 && v$G18_13514_out0;
assign v$G29_5485_out0 = v$G32_1826_out0 && v$R3_15314_out0;
assign v$G29_5486_out0 = v$G32_1827_out0 && v$R3_15315_out0;
assign v$G9_5798_out0 = ! v$INTERRUPT0_11700_out0;
assign v$G9_5799_out0 = ! v$INTERRUPT0_11701_out0;
assign v$MUX17_6531_out0 = v$IS$IR1$FMUL_15296_out0 ? v$IR1$32$BITS_7867_out0 : v$IR2$FPU$32BIT_11800_out0;
assign v$EDGE2_6999_out0 = v$INTERRUPT2_3853_out0;
assign v$G5_7583_out0 = v$G3_2671_out0 && v$IR15_10986_out0;
assign v$G5_7584_out0 = v$G3_2672_out0 && v$IR15_10987_out0;
assign v$G20_12209_out0 = v$EQ5_14374_out0 && v$IR1$L_5138_out0;
assign v$G20_12210_out0 = v$EQ5_14375_out0 && v$IR1$L_5139_out0;
assign v$SUBEN_12858_out0 = v$G8_18779_out0;
assign v$SUBEN_12859_out0 = v$G8_18780_out0;
assign v$STALL_13145_out0 = v$G27_16528_out0;
assign v$STALL_13146_out0 = v$G27_16529_out0;
assign v$G3_14181_out0 = v$EQ3_17921_out0 && v$G2_18429_out0;
assign v$G3_14182_out0 = v$EQ3_17922_out0 && v$G2_18430_out0;
assign v$G7_14673_out0 = v$INTERRUPT0_11700_out0 && v$G1_14473_out0;
assign v$G7_14674_out0 = v$INTERRUPT0_11701_out0 && v$G1_14474_out0;
assign v$G5_15792_out0 = ! v$IS$32$BIT_10863_out0;
assign v$G30_15903_out0 = v$FF4_18438_out0 && v$G28_3167_out0;
assign v$G30_15904_out0 = v$FF4_18439_out0 && v$G28_3168_out0;
assign v$IS$32$BITS_17584_out0 = v$IS$32$BITS_1282_out0;
assign v$STP_17762_out0 = v$STP_11714_out0;
assign v$STP_17763_out0 = v$STP_11715_out0;
assign v$G15_18535_out0 = v$IR1$P_3692_out0 || v$G16_11965_out0;
assign v$G15_18536_out0 = v$IR1$P_3693_out0 || v$G16_11966_out0;
assign v$OP_1324_out0 = v$MUX11_4488_out0;
assign v$INTERRUPT2_1663_out0 = v$EDGE2_6999_out0;
assign v$G27_2512_out0 = v$G30_15903_out0 && v$F3_8247_out0;
assign v$G27_2513_out0 = v$G30_15904_out0 && v$F3_8248_out0;
assign v$IS$32$BITS_4149_out0 = v$IS$32$BITS_17584_out0;
assign v$G8_6047_out0 = v$G7_14673_out0 && v$R0_15192_out0;
assign v$G8_6048_out0 = v$G7_14674_out0 && v$R0_15193_out0;
assign v$G43_7051_out0 = v$STALL_13145_out0 && v$IR2$VALID_4217_out0;
assign v$G43_7052_out0 = v$STALL_13146_out0 && v$IR2$VALID_4218_out0;
assign v$STP_10818_out0 = v$STP_17762_out0;
assign v$STP_10819_out0 = v$STP_17763_out0;
assign v$32BIT_10932_out0 = v$MUX17_6531_out0;
assign v$MUX1_11751_out0 = v$SUBEN_12858_out0 ? v$C2_12207_out0 : v$C1_18208_out0;
assign v$MUX1_11752_out0 = v$SUBEN_12859_out0 ? v$C2_12208_out0 : v$C1_18209_out0;
assign v$G10_13314_out0 = v$FF1_6026_out0 && v$G9_5798_out0;
assign v$G10_13315_out0 = v$FF1_6027_out0 && v$G9_5799_out0;
assign v$G26_18115_out0 = v$IS$IR1$FMUL_15296_out0 && v$G27_3882_out0;
assign v$QP_18537_out0 = v$_1231_out0;
assign v$QP_18538_out0 = v$_1232_out0;
assign v$G10_1182_out0 = v$EQ11_13605_out0 && v$STP_10818_out0;
assign v$G10_1183_out0 = v$EQ11_13606_out0 && v$STP_10819_out0;
assign v$G33_1233_out0 = v$G29_5485_out0 || v$G27_2512_out0;
assign v$G33_1234_out0 = v$G29_5486_out0 || v$G27_2513_out0;
assign v$G11_1619_out0 = v$G10_13314_out0 && v$F0_15834_out0;
assign v$G11_1620_out0 = v$G10_13315_out0 && v$F0_15835_out0;
assign v$G8_2243_out0 = v$EQ9_17768_out0 && v$STP_10818_out0;
assign v$G8_2244_out0 = v$EQ9_17769_out0 && v$STP_10819_out0;
assign v$G7_3159_out0 = v$EQ10_13408_out0 && v$STP_10818_out0;
assign v$G7_3160_out0 = v$EQ10_13409_out0 && v$STP_10819_out0;
assign v$MUX11_4487_out0 = v$G26_18115_out0 ? v$IR1$FPU$OP_3837_out0 : v$IR2$FPU$OP_1687_out0;
assign v$G12_4833_out0 = v$G43_7051_out0 && v$INITIAL$FETCH$OCCURRED_1537_out0;
assign v$G12_4834_out0 = v$G43_7052_out0 && v$INITIAL$FETCH$OCCURRED_1538_out0;
assign v$XOR1_5078_out0 = v$MUX1_11751_out0 ^ v$DIN_1723_out0;
assign v$XOR1_5079_out0 = v$MUX1_11752_out0 ^ v$DIN_1724_out0;
assign v$G6_5464_out0 = v$EQ7_16898_out0 && v$STP_10818_out0;
assign v$G6_5465_out0 = v$EQ7_16899_out0 && v$STP_10819_out0;
assign v$G14_6428_out0 = v$EQ13_18548_out0 && v$STP_10818_out0;
assign v$G14_6429_out0 = v$EQ13_18549_out0 && v$STP_10819_out0;
assign v$G21_7036_out0 = ! v$INTERRUPT2_1663_out0;
assign v$EQ5_10028_out0 = v$QP_18537_out0 == 4'hb;
assign v$EQ5_10029_out0 = v$QP_18538_out0 == 4'hb;
assign v$FPU$OP_14069_out0 = v$OP_1324_out0;
assign v$G25_14578_out0 = v$INTERRUPT2_1663_out0 && v$G24_12087_out0;
assign v$G9_15125_out0 = v$EQ8_14328_out0 && v$STP_10818_out0;
assign v$G9_15126_out0 = v$EQ8_14329_out0 && v$STP_10819_out0;
assign v$32BIT_15872_out0 = v$32BIT_10932_out0;
assign v$OP_1323_out0 = v$MUX11_4487_out0;
assign v$G37_1360_out0 = v$G12_4833_out0 && v$G48_4876_out0;
assign v$G37_1361_out0 = v$G12_4834_out0 && v$G48_4877_out0;
assign v$EQ5_2969_out0 = v$FPU$OP_14069_out0 == 2'h3;
assign v$EQ2_4230_out0 = v$FPU$OP_14069_out0 == 2'h0;
assign v$INTDISABLE_4999_out0 = v$G7_3159_out0;
assign v$INTDISABLE_5000_out0 = v$G7_3160_out0;
assign v$G22_5462_out0 = v$G25_14578_out0 && v$R2_3845_out0;
assign v$NEXTINT_7001_out0 = v$G10_1182_out0;
assign v$NEXTINT_7002_out0 = v$G10_1183_out0;
assign v$INTCLEAR_7775_out0 = v$G8_2243_out0;
assign v$INTCLEAR_7776_out0 = v$G8_2244_out0;
assign v$G23_9601_out0 = v$FF3_15030_out0 && v$G21_7036_out0;
assign v$G29_10829_out0 = v$32BIT_15872_out0 && v$IR2$IS$FPU_11843_out0;
assign v$IS$32$BIT_11005_out0 = v$32BIT_15872_out0;
assign v$EDGE3_11040_out0 = v$G33_1233_out0;
assign v$EDGE3_11041_out0 = v$G33_1234_out0;
assign v$FPU$OP_12763_out0 = v$FPU$OP_14069_out0;
assign v$LDMAINPC_13634_out0 = v$G14_6428_out0;
assign v$LDMAINPC_13635_out0 = v$G14_6429_out0;
assign v$EQ3_13794_out0 = v$FPU$OP_14069_out0 == 2'h2;
assign v$IS$32$BITS_14038_out0 = v$32BIT_15872_out0;
assign v$G12_14705_out0 = v$G8_6047_out0 || v$G11_1619_out0;
assign v$G12_14706_out0 = v$G8_6048_out0 || v$G11_1620_out0;
assign v$EQ1_15290_out0 = v$FPU$OP_14069_out0 == 2'h1;
assign v$EQ6_16172_out0 = v$FPU$OP_14069_out0 == 2'h3;
assign v$EQ4_16702_out0 = v$FPU$OP_14069_out0 == 2'h3;
assign v$G66_16844_out0 = !(v$G69_1206_out0 && v$EQ5_10028_out0);
assign v$G66_16845_out0 = !(v$G69_1207_out0 && v$EQ5_10029_out0);
assign v$NEXTINTERRUPT_18546_out0 = v$G10_1182_out0;
assign v$NEXTINTERRUPT_18547_out0 = v$G10_1183_out0;
assign v$INTCLR_214_out0 = v$INTCLEAR_7775_out0;
assign v$INTCLR_215_out0 = v$INTCLEAR_7776_out0;
assign v$G35_1145_out0 = v$G37_1360_out0 && v$G36_17349_out0;
assign v$G35_1146_out0 = v$G37_1361_out0 && v$G36_17350_out0;
assign v$G8_1248_out0 = v$EQ4_16702_out0 && v$LOADA_5077_out0;
assign v$INTDISABLE_2684_out0 = v$INTDISABLE_4999_out0;
assign v$INTDISABLE_2685_out0 = v$INTDISABLE_5000_out0;
assign v$G16_3839_out0 = ! v$EQ6_16172_out0;
assign v$EDGE0_3990_out0 = v$G12_14705_out0;
assign v$EDGE0_3991_out0 = v$G12_14706_out0;
assign v$G34_4917_out0 = v$NEXTINTERRUPT_18546_out0 || v$FF2_1180_out0;
assign v$G34_4918_out0 = v$NEXTINTERRUPT_18547_out0 || v$FF2_1181_out0;
assign v$ADD_8220_out0 = v$EQ2_4230_out0;
assign v$IS$32$BIT_10862_out0 = v$IS$32$BIT_11005_out0;
assign v$FPU$LOAD$STORE_10980_out0 = v$EQ4_16702_out0;
assign v$G20_11710_out0 = v$G23_9601_out0 && v$F2_12096_out0;
assign v$G12_11979_out0 = v$G11_13407_out0 && v$EQ5_2969_out0;
assign v$G15_13420_out0 = v$G6_5464_out0 || v$NEXTINT_7001_out0;
assign v$G15_13421_out0 = v$G6_5465_out0 || v$NEXTINT_7002_out0;
assign v$SUB_13791_out0 = v$EQ1_15290_out0;
assign v$LDMAIN_13807_out0 = v$LDMAINPC_13634_out0;
assign v$LDMAIN_13808_out0 = v$LDMAINPC_13635_out0;
assign v$FPU$OP_14068_out0 = v$OP_1323_out0;
assign v$G65_14120_out0 = v$G66_16844_out0 && v$CLK4_2531_out0;
assign v$G65_14121_out0 = v$G66_16845_out0 && v$CLK4_2532_out0;
assign v$EQ1_16220_out0 = v$FPU$OP_12763_out0 == 2'h1;
assign v$G9_16964_out0 = v$EQ4_16702_out0 && v$G10_14589_out0;
assign v$MUL_17035_out0 = v$EQ3_13794_out0;
assign v$CLRINTERRUPTS_340_out0 = v$INTCLR_214_out0;
assign v$CLRINTERRUPTS_341_out0 = v$INTCLR_215_out0;
assign v$INTENABLE_2939_out0 = v$G15_13420_out0;
assign v$INTENABLE_2940_out0 = v$G15_13421_out0;
assign v$EQ5_2968_out0 = v$FPU$OP_14068_out0 == 2'h3;
assign v$G2_3725_out0 = v$ADD_8220_out0 || v$SUB_13791_out0;
assign v$EQ2_4229_out0 = v$FPU$OP_14068_out0 == 2'h0;
assign v$G17_5521_out0 = v$G15_2283_out0 && v$G16_3839_out0;
assign v$G13_7895_out0 = v$G9_16964_out0 && v$IR2$IS$FPU_11844_out0;
assign v$G6_7940_out0 = v$ADD_8220_out0 || v$SUB_13791_out0;
assign v$G26_10319_out0 = v$G22_5462_out0 || v$G20_11710_out0;
assign v$G35_10321_out0 = v$INTDISABLE_2684_out0 || v$AUTODISABLE_18213_out0;
assign v$G35_10322_out0 = v$INTDISABLE_2685_out0 || v$AUTODISABLE_18214_out0;
assign v$STOPBITERROR_11727_out0 = v$G65_14120_out0;
assign v$STOPBITERROR_11728_out0 = v$G65_14121_out0;
assign v$FPU$OP_12762_out0 = v$FPU$OP_14068_out0;
assign v$EQ7_13602_out0 = v$FPU$OP_14068_out0 == 2'h2;
assign v$EQ3_13793_out0 = v$FPU$OP_14068_out0 == 2'h2;
assign v$G21_14711_out0 = v$G20_12293_out0 && v$FPU$LOAD$STORE_10980_out0;
assign v$EQ1_15289_out0 = v$FPU$OP_14068_out0 == 2'h1;
assign v$G5_15791_out0 = ! v$IS$32$BIT_10862_out0;
assign v$G14_15816_out0 = v$G8_1248_out0 && v$IR2$IS$FPU_11844_out0;
assign v$EQ8_16018_out0 = v$FPU$OP_14068_out0 == 2'h3;
assign v$EQ4_16701_out0 = v$FPU$OP_14068_out0 == 2'h3;
assign v$STALL_17890_out0 = v$G35_1145_out0;
assign v$STALL_17891_out0 = v$G35_1146_out0;
assign v$NEXTINTERRUPT_18433_out0 = v$G34_4917_out0;
assign v$NEXTINTERRUPT_18434_out0 = v$G34_4918_out0;
assign v$STOPERROR_294_out0 = v$STOPBITERROR_11727_out0;
assign v$STOPERROR_295_out0 = v$STOPBITERROR_11728_out0;
assign v$G30_3764_out0 = ! v$EQ8_16018_out0;
assign v$CLR_4434_out0 = v$CLRINTERRUPTS_340_out0;
assign v$CLR_4435_out0 = v$CLRINTERRUPTS_341_out0;
assign v$G49_5244_out0 = ! v$STALL_17890_out0;
assign v$G49_5245_out0 = ! v$STALL_17891_out0;
assign v$G18_7510_out0 = v$G17_5521_out0 && v$IR2$VALID_15879_out0;
assign v$ADD_8219_out0 = v$EQ2_4229_out0;
assign v$G3_9357_out0 = v$MUL_17035_out0 || v$G6_7940_out0;
assign v$FPU$LOAD$STORE_10979_out0 = v$EQ4_16701_out0;
assign v$G12_11978_out0 = v$G11_13406_out0 && v$EQ5_2968_out0;
assign v$NEXTINTERRUPT_12752_out0 = v$NEXTINTERRUPT_18433_out0;
assign v$NEXTINTERRUPT_12753_out0 = v$NEXTINTERRUPT_18434_out0;
assign v$SUB_13790_out0 = v$EQ1_15289_out0;
assign v$DISABLEINTERRUPTS_14974_out0 = v$G35_10321_out0;
assign v$DISABLEINTERRUPTS_14975_out0 = v$G35_10322_out0;
assign v$STALL_15494_out0 = v$STALL_17890_out0;
assign v$STALL_15495_out0 = v$STALL_17891_out0;
assign v$EQ1_16219_out0 = v$FPU$OP_12762_out0 == 2'h1;
assign v$MUL_17034_out0 = v$EQ3_13793_out0;
assign v$INTENABLE_17402_out0 = v$INTENABLE_2939_out0;
assign v$INTENABLE_17403_out0 = v$INTENABLE_2940_out0;
assign v$EDGE2_18118_out0 = v$G26_10319_out0;
assign v$G31_2344_out0 = v$G29_10829_out0 && v$G30_3764_out0;
assign v$G2_3724_out0 = v$ADD_8219_out0 || v$SUB_13790_out0;
assign v$G4_4900_out0 = v$ERR_12774_out0 || v$STOPERROR_294_out0;
assign v$G4_4901_out0 = v$ERR_12775_out0 || v$STOPERROR_295_out0;
assign v$G6_7939_out0 = v$ADD_8219_out0 || v$SUB_13790_out0;
assign v$G28_8690_out0 = v$FPU$LOAD$STORE_10979_out0 && v$LOAD_6190_out0;
assign v$G27_10726_out0 = v$FPU$LOAD$STORE_10979_out0 && v$LOAD_6190_out0;
assign v$G27_11708_out0 = v$STP$DECODED_16534_out0 || v$G49_5244_out0;
assign v$G27_11709_out0 = v$STP$DECODED_16535_out0 || v$G49_5245_out0;
assign v$STALL_12230_out0 = v$STALL_15494_out0;
assign v$STALL_12231_out0 = v$STALL_15495_out0;
assign v$ENABLEINTERRUPTS_12547_out0 = v$INTENABLE_17402_out0;
assign v$ENABLEINTERRUPTS_12548_out0 = v$INTENABLE_17403_out0;
assign v$G21_14710_out0 = v$G20_12292_out0 && v$FPU$LOAD$STORE_10979_out0;
assign v$G19_15875_out0 = v$G21_14711_out0 || v$G3_9357_out0;
assign v$NEXTINTERRUPT_16777_out0 = v$NEXTINTERRUPT_12752_out0;
assign v$NEXTINTERRUPT_16778_out0 = v$NEXTINTERRUPT_12753_out0;
assign v$R_18332_out0 = v$DISABLEINTERRUPTS_14974_out0;
assign v$R_18335_out0 = v$CLR_4434_out0;
assign v$R_18343_out0 = v$DISABLEINTERRUPTS_14975_out0;
assign v$R_18346_out0 = v$CLR_4435_out0;
assign v$G8_1247_out0 = v$G27_10726_out0 && v$LOADA_5076_out0;
assign v$G7_1499_out0 = v$G19_15875_out0 && v$IR2$VALID_15879_out0;
assign v$G3_4104_out0 = v$I0P_4347_out0 && v$NEXTINTERRUPT_16777_out0;
assign v$G3_4105_out0 = v$I0P_4348_out0 && v$NEXTINTERRUPT_16778_out0;
assign v$G1_7223_out0 = v$I2P_7492_out0 && v$NEXTINTERRUPT_16777_out0;
assign v$G1_7224_out0 = v$I2P_7493_out0 && v$NEXTINTERRUPT_16778_out0;
assign v$G2_8334_out0 = v$I3P_10827_out0 && v$NEXTINTERRUPT_16777_out0;
assign v$G2_8335_out0 = v$I3P_10828_out0 && v$NEXTINTERRUPT_16778_out0;
assign v$G3_9940_out0 = v$INITIAL$FETCH$OCCURRED_1537_out0 && v$G27_11708_out0;
assign v$G3_9941_out0 = v$INITIAL$FETCH$OCCURRED_1538_out0 && v$G27_11709_out0;
assign v$PIPELINEHALT_14816_out0 = v$STALL_12230_out0;
assign v$PIPELINEHALT_14817_out0 = v$STALL_12231_out0;
assign v$G4_15457_out0 = v$I1P_2514_out0 && v$NEXTINTERRUPT_16777_out0;
assign v$G4_15458_out0 = v$I1P_2515_out0 && v$NEXTINTERRUPT_16778_out0;
assign v$G6_15560_out0 = ! v$R_18332_out0;
assign v$G6_15563_out0 = ! v$R_18335_out0;
assign v$G6_15571_out0 = ! v$R_18343_out0;
assign v$G6_15574_out0 = ! v$R_18346_out0;
assign v$G19_15874_out0 = v$G21_14710_out0 || v$G6_7939_out0;
assign v$G32_16333_out0 = v$G31_2344_out0 && v$IR2$VALID_15878_out0;
assign v$S_16931_out0 = v$ENABLEINTERRUPTS_12547_out0;
assign v$S_16942_out0 = v$ENABLEINTERRUPTS_12548_out0;
assign v$G9_16963_out0 = v$G28_8690_out0 && v$G10_14588_out0;
assign v$SetError_17573_out0 = v$G4_4900_out0;
assign v$SetError_17574_out0 = v$G4_4901_out0;
assign v$G7_1498_out0 = v$G19_15874_out0 && v$IR2$VALID_15878_out0;
assign v$G9_2527_out0 = v$CLR_4434_out0 || v$G4_15457_out0;
assign v$G9_2528_out0 = v$CLR_4435_out0 || v$G4_15458_out0;
assign v$G11_3012_out0 = v$CLR_4434_out0 || v$G2_8334_out0;
assign v$G11_3013_out0 = v$CLR_4435_out0 || v$G2_8335_out0;
assign v$G10_6689_out0 = v$CLR_4434_out0 || v$G1_7223_out0;
assign v$G10_6690_out0 = v$CLR_4435_out0 || v$G1_7224_out0;
assign v$G13_7894_out0 = v$G9_16963_out0 && v$IR2$IS$FPU_11843_out0;
assign v$SHOULD$STORE_12710_out0 = v$G32_16333_out0;
assign v$WENFPU_13740_out0 = v$G7_1499_out0;
assign v$G8_14257_out0 = v$FF2_13040_out0 || v$S_16931_out0;
assign v$G8_14263_out0 = v$FF2_13051_out0 || v$S_16942_out0;
assign v$G8_15479_out0 = v$CLR_4434_out0 || v$G3_4104_out0;
assign v$G8_15480_out0 = v$CLR_4435_out0 || v$G3_4105_out0;
assign v$G14_15815_out0 = v$G8_1247_out0 && v$IR2$IS$FPU_11843_out0;
assign v$G50_16361_out0 = v$G51_14015_out0 && v$G3_9940_out0;
assign v$G50_16362_out0 = v$G51_14016_out0 && v$G3_9941_out0;
assign v$S_16940_out0 = v$SetError_17573_out0;
assign v$S_16951_out0 = v$SetError_17574_out0;
assign v$G24_240_out0 = v$G7_1498_out0 && v$G26_5127_out0;
assign v$G33_324_out0 = v$FINISHED_8010_out0 || v$SHOULD$STORE_12710_out0;
assign v$WENFPU_3499_out0 = v$WENFPU_13740_out0;
assign v$G7_14123_out0 = v$G8_14257_out0 && v$G6_15560_out0;
assign v$G7_14129_out0 = v$G8_14263_out0 && v$G6_15571_out0;
assign v$IR1$VALID_17797_out0 = v$G50_16361_out0;
assign v$IR1$VALID_17798_out0 = v$G50_16362_out0;
assign v$R_18331_out0 = v$G8_15479_out0;
assign v$R_18333_out0 = v$G10_6689_out0;
assign v$R_18334_out0 = v$G11_3012_out0;
assign v$R_18336_out0 = v$G9_2527_out0;
assign v$R_18342_out0 = v$G8_15480_out0;
assign v$R_18344_out0 = v$G10_6690_out0;
assign v$R_18345_out0 = v$G11_3013_out0;
assign v$R_18347_out0 = v$G9_2528_out0;
assign v$IR1$VALID_9455_out0 = v$IR1$VALID_17797_out0;
assign v$IR1$VALID_9456_out0 = v$IR1$VALID_17798_out0;
assign v$WENFPU_13739_out0 = v$G24_240_out0;
assign v$Q_14141_out0 = v$G7_14123_out0;
assign v$Q_14152_out0 = v$G7_14129_out0;
assign v$G6_15559_out0 = ! v$R_18331_out0;
assign v$G6_15561_out0 = ! v$R_18333_out0;
assign v$G6_15562_out0 = ! v$R_18334_out0;
assign v$G6_15564_out0 = ! v$R_18336_out0;
assign v$G6_15570_out0 = ! v$R_18342_out0;
assign v$G6_15572_out0 = ! v$R_18344_out0;
assign v$G6_15573_out0 = ! v$R_18345_out0;
assign v$G6_15575_out0 = ! v$R_18347_out0;
assign v$WENFPU_3498_out0 = v$WENFPU_13739_out0;
assign v$IR1$VALID_5751_out0 = v$IR1$VALID_9455_out0;
assign v$IR1$VALID_5752_out0 = v$IR1$VALID_9456_out0;
assign v$ENABLEINTERRUPTS_17026_out0 = v$Q_14141_out0;
assign v$ENABLEINTERRUPTS_17027_out0 = v$Q_14152_out0;
assign v$G19_336_out0 = v$EDGE0_3990_out0 && v$ENABLEINTERRUPTS_17026_out0;
assign v$G19_337_out0 = v$EDGE0_3991_out0 && v$ENABLEINTERRUPTS_17027_out0;
assign v$G22_4882_out0 = v$EDGE3_11040_out0 && v$ENABLEINTERRUPTS_17026_out0;
assign v$G22_4883_out0 = v$EDGE3_11041_out0 && v$ENABLEINTERRUPTS_17027_out0;
assign v$IR1$VALID_14013_out0 = v$IR1$VALID_5751_out0;
assign v$IR1$VALID_14014_out0 = v$IR1$VALID_5752_out0;
assign v$G21_15822_out0 = v$EDGE2_18118_out0 && v$ENABLEINTERRUPTS_17026_out0;
assign v$G21_15823_out0 = v$EDGE2_18119_out0 && v$ENABLEINTERRUPTS_17027_out0;
assign v$G20_15936_out0 = v$EDGE1_15272_out0 && v$ENABLEINTERRUPTS_17026_out0;
assign v$G20_15937_out0 = v$EDGE1_15273_out0 && v$ENABLEINTERRUPTS_17027_out0;
assign v$G13_4351_out0 = v$G21_15822_out0 || v$G22_4882_out0;
assign v$G13_4352_out0 = v$G21_15823_out0 || v$G22_4883_out0;
assign v$G24_7896_out0 = v$LASTQ_12100_out0 && v$G21_15822_out0;
assign v$G24_7897_out0 = v$LASTQ_12111_out0 && v$G21_15823_out0;
assign v$G12_11896_out0 = v$G19_336_out0 || v$G20_15936_out0;
assign v$G12_11897_out0 = v$G19_337_out0 || v$G20_15937_out0;
assign v$G26_12654_out0 = v$LASTQ_12098_out0 && v$G19_336_out0;
assign v$G26_12655_out0 = v$LASTQ_12109_out0 && v$G19_337_out0;
assign v$G25_13011_out0 = v$LASTQ_12103_out0 && v$G20_15936_out0;
assign v$G25_13012_out0 = v$LASTQ_12114_out0 && v$G20_15937_out0;
assign v$S_16930_out0 = v$G19_336_out0;
assign v$S_16932_out0 = v$G21_15822_out0;
assign v$S_16933_out0 = v$G22_4882_out0;
assign v$S_16935_out0 = v$G20_15936_out0;
assign v$S_16941_out0 = v$G19_337_out0;
assign v$S_16943_out0 = v$G21_15823_out0;
assign v$S_16944_out0 = v$G22_4883_out0;
assign v$S_16946_out0 = v$G20_15937_out0;
assign v$IR1$VALID_18427_out0 = v$IR1$VALID_14013_out0;
assign v$IR1$VALID_18428_out0 = v$IR1$VALID_14014_out0;
assign v$G23_18654_out0 = v$LASTQ_12101_out0 && v$G22_4882_out0;
assign v$G23_18655_out0 = v$LASTQ_12112_out0 && v$G22_4883_out0;
assign v$G6_269_out0 = v$G5_16556_out0 && v$IR1$VALID_18427_out0;
assign v$G6_270_out0 = v$G5_16557_out0 && v$IR1$VALID_18428_out0;
assign v$IR1$VALID_3847_out0 = v$IR1$VALID_18427_out0;
assign v$IR1$VALID_3848_out0 = v$IR1$VALID_18428_out0;
assign v$G23_6992_out0 = v$EQ8_252_out0 && v$IR1$VALID_18427_out0;
assign v$G23_6993_out0 = v$EQ8_253_out0 && v$IR1$VALID_18428_out0;
assign v$G7_9938_out0 = v$IR1$VALID_18427_out0 && v$IS$IR1$FMUL_15296_out0;
assign v$G7_9939_out0 = v$IR1$VALID_18428_out0 && v$IS$IR1$FMUL_15297_out0;
assign v$G8_14256_out0 = v$FF2_13039_out0 || v$S_16930_out0;
assign v$G8_14258_out0 = v$FF2_13041_out0 || v$S_16932_out0;
assign v$G8_14259_out0 = v$FF2_13042_out0 || v$S_16933_out0;
assign v$G8_14261_out0 = v$FF2_13044_out0 || v$S_16935_out0;
assign v$G8_14262_out0 = v$FF2_13050_out0 || v$S_16941_out0;
assign v$G8_14264_out0 = v$FF2_13052_out0 || v$S_16943_out0;
assign v$G8_14265_out0 = v$FF2_13053_out0 || v$S_16944_out0;
assign v$G8_14267_out0 = v$FF2_13055_out0 || v$S_16946_out0;
assign v$G14_15291_out0 = v$G12_11896_out0 || v$G13_4351_out0;
assign v$G14_15292_out0 = v$G12_11897_out0 || v$G13_4352_out0;
assign v$G28_15384_out0 = v$G24_7896_out0 || v$G23_18654_out0;
assign v$G28_15385_out0 = v$G24_7897_out0 || v$G23_18655_out0;
assign v$G27_18489_out0 = v$G26_12654_out0 || v$G25_13011_out0;
assign v$G27_18490_out0 = v$G26_12655_out0 || v$G25_13012_out0;
assign v$IR1$VALID_61_out0 = v$IR1$VALID_3847_out0;
assign v$IR1$VALID_62_out0 = v$IR1$VALID_3848_out0;
assign v$INCOMINGINTERRUPT_1903_out0 = v$G14_15291_out0;
assign v$INCOMINGINTERRUPT_1904_out0 = v$G14_15292_out0;
assign v$MUX9_7648_out0 = v$G6_269_out0 ? v$IR1$D_4219_out0 : v$IR2$D_14491_out0;
assign v$MUX9_7649_out0 = v$G6_270_out0 ? v$IR1$D_4220_out0 : v$IR2$D_14492_out0;
assign v$G8_12482_out0 = v$G10_10271_out0 || v$G6_269_out0;
assign v$G8_12483_out0 = v$G10_10272_out0 || v$G6_270_out0;
assign v$EXEC1$FPU_13675_out0 = v$G7_9938_out0;
assign v$EXEC1$FPU_13676_out0 = v$G7_9939_out0;
assign v$G7_14122_out0 = v$G8_14256_out0 && v$G6_15559_out0;
assign v$G7_14124_out0 = v$G8_14258_out0 && v$G6_15561_out0;
assign v$G7_14125_out0 = v$G8_14259_out0 && v$G6_15562_out0;
assign v$G7_14127_out0 = v$G8_14261_out0 && v$G6_15564_out0;
assign v$G7_14128_out0 = v$G8_14262_out0 && v$G6_15570_out0;
assign v$G7_14130_out0 = v$G8_14264_out0 && v$G6_15572_out0;
assign v$G7_14131_out0 = v$G8_14265_out0 && v$G6_15573_out0;
assign v$G7_14133_out0 = v$G8_14267_out0 && v$G6_15575_out0;
assign v$G29_15774_out0 = v$G27_18489_out0 || v$G28_15384_out0;
assign v$G29_15775_out0 = v$G27_18490_out0 || v$G28_15385_out0;
assign v$INTERRUPTOVERFLOW_2233_out0 = v$G29_15774_out0;
assign v$INTERRUPTOVERFLOW_2234_out0 = v$G29_15775_out0;
assign v$G19_2826_out0 = v$G20_12209_out0 && v$IR1$VALID_61_out0;
assign v$G19_2827_out0 = v$G20_12210_out0 && v$IR1$VALID_62_out0;
assign v$AD1_6656_out0 = v$MUX9_7648_out0;
assign v$AD1_6657_out0 = v$MUX9_7649_out0;
assign v$G13_10230_out0 = v$G8_12482_out0 || v$G23_6992_out0;
assign v$G13_10231_out0 = v$G8_12483_out0 || v$G23_6993_out0;
assign v$EXEC1_10256_out0 = v$EXEC1$FPU_13675_out0;
assign v$EXEC1_10257_out0 = v$EXEC1$FPU_13676_out0;
assign v$G17_12139_out0 = v$INCOMINGINTERRUPT_1903_out0 && v$G18_2988_out0;
assign v$G17_12140_out0 = v$INCOMINGINTERRUPT_1904_out0 && v$G18_2989_out0;
assign v$Q_14140_out0 = v$G7_14122_out0;
assign v$Q_14142_out0 = v$G7_14124_out0;
assign v$Q_14143_out0 = v$G7_14125_out0;
assign v$Q_14145_out0 = v$G7_14127_out0;
assign v$Q_14151_out0 = v$G7_14128_out0;
assign v$Q_14153_out0 = v$G7_14130_out0;
assign v$Q_14154_out0 = v$G7_14131_out0;
assign v$Q_14156_out0 = v$G7_14133_out0;
assign v$G5_14649_out0 = v$IR1$VALID_61_out0 && v$IR1$W_16548_out0;
assign v$G5_14650_out0 = v$IR1$VALID_62_out0 && v$IR1$W_16549_out0;
assign v$G4_15544_out0 = v$G3_14181_out0 && v$IR1$VALID_61_out0;
assign v$G4_15545_out0 = v$G3_14182_out0 && v$IR1$VALID_62_out0;
assign v$MUX10_3626_out0 = v$G13_10230_out0 ? v$IR1$M_13247_out0 : v$IR2$M_12993_out0;
assign v$MUX10_3627_out0 = v$G13_10231_out0 ? v$IR1$M_13248_out0 : v$IR2$M_12994_out0;
assign v$I3_4823_out0 = v$Q_14143_out0;
assign v$I3_4824_out0 = v$Q_14154_out0;
assign v$I1_4890_out0 = v$Q_14145_out0;
assign v$I1_4891_out0 = v$Q_14156_out0;
assign v$NEWINTERRUPT_5432_out0 = v$G17_12139_out0;
assign v$NEWINTERRUPT_5433_out0 = v$G17_12140_out0;
assign v$G16_6391_out0 = v$NEXTINTERRUPT_16777_out0 || v$G17_12139_out0;
assign v$G16_6392_out0 = v$NEXTINTERRUPT_16778_out0 || v$G17_12140_out0;
assign v$G6_7480_out0 = v$Q_14142_out0 || v$Q_14143_out0;
assign v$G6_7481_out0 = v$Q_14153_out0 || v$Q_14154_out0;
assign v$G7_11796_out0 = v$G5_14649_out0 || v$G6_11934_out0;
assign v$G7_11797_out0 = v$G5_14650_out0 || v$G6_11935_out0;
assign v$READ$REQUEST_14458_out0 = v$G19_2826_out0;
assign v$READ$REQUEST_14459_out0 = v$G19_2827_out0;
assign v$I2_14493_out0 = v$Q_14142_out0;
assign v$I2_14494_out0 = v$Q_14153_out0;
assign v$G11_14584_out0 = v$G4_15544_out0 && v$G10_14893_out0;
assign v$G11_14585_out0 = v$G4_15545_out0 && v$G10_14894_out0;
assign v$G23_15947_out0 = v$EXEC1_10256_out0 && v$EQ7_13602_out0;
assign v$G5_16118_out0 = v$Q_14140_out0 || v$Q_14145_out0;
assign v$G5_16119_out0 = v$Q_14151_out0 || v$Q_14156_out0;
assign v$S_16934_out0 = v$INTERRUPTOVERFLOW_2233_out0;
assign v$S_16945_out0 = v$INTERRUPTOVERFLOW_2234_out0;
assign v$I0_18506_out0 = v$Q_14140_out0;
assign v$I0_18507_out0 = v$Q_14151_out0;
assign v$AD1_18672_out0 = v$AD1_6656_out0;
assign v$AD1_18673_out0 = v$AD1_6657_out0;
assign v$EXEC1_18719_out0 = v$EXEC1_10257_out0;
assign v$CAPTURE_242_out0 = v$G16_6391_out0;
assign v$CAPTURE_243_out0 = v$G16_6392_out0;
assign v$G7_1831_out0 = v$G5_16118_out0 || v$G6_7480_out0;
assign v$G7_1832_out0 = v$G5_16119_out0 || v$G6_7481_out0;
assign v$AD1_1840_out0 = v$AD1_18672_out0;
assign v$AD1_1841_out0 = v$AD1_18673_out0;
assign v$START_3700_out0 = v$G23_15947_out0;
assign v$NEWINTERRUPT_7025_out0 = v$NEWINTERRUPT_5432_out0;
assign v$NEWINTERRUPT_7026_out0 = v$NEWINTERRUPT_5433_out0;
assign v$G4_7739_out0 = ! v$I1_4890_out0;
assign v$G4_7740_out0 = ! v$I1_4891_out0;
assign v$RAMWEN_7764_out0 = v$G11_14584_out0;
assign v$RAMWEN_7765_out0 = v$G11_14585_out0;
assign v$G2_7777_out0 = ! v$I3_4823_out0;
assign v$G2_7778_out0 = ! v$I3_4824_out0;
assign v$G3_8822_out0 = ! v$I2_14493_out0;
assign v$G3_8823_out0 = ! v$I2_14494_out0;
assign v$AD2_9095_out0 = v$MUX10_3626_out0;
assign v$AD2_9096_out0 = v$MUX10_3627_out0;
assign v$WENLDST_12484_out0 = v$G7_11796_out0;
assign v$WENLDST_12485_out0 = v$G7_11797_out0;
assign v$I3P_13619_out0 = v$I3_4823_out0;
assign v$I3P_13620_out0 = v$I3_4824_out0;
assign v$G8_14260_out0 = v$FF2_13043_out0 || v$S_16934_out0;
assign v$G8_14266_out0 = v$FF2_13054_out0 || v$S_16945_out0;
assign v$READ$REQUEST_16552_out0 = v$READ$REQUEST_14458_out0;
assign v$READ$REQUEST_16553_out0 = v$READ$REQUEST_14459_out0;
assign v$EXEC1_18224_out0 = v$EXEC1_18719_out0;
assign v$EXEC1_3855_out0 = v$EXEC1_18224_out0;
assign v$NEWINTERRUPT_4431_out0 = v$NEWINTERRUPT_7025_out0;
assign v$NEWINTERRUPT_4432_out0 = v$NEWINTERRUPT_7026_out0;
assign v$MUX1_5013_out0 = v$G16_6391_out0 ? v$G7_1831_out0 : v$FF1_13095_out0;
assign v$MUX1_5014_out0 = v$G16_6392_out0 ? v$G7_1832_out0 : v$FF1_13096_out0;
assign v$READ$REQUEST_7806_out0 = v$READ$REQUEST_16552_out0;
assign v$READ$REQUEST_7807_out0 = v$READ$REQUEST_16553_out0;
assign v$G7_10967_out0 = v$I0_18506_out0 && v$G4_7739_out0;
assign v$G7_10968_out0 = v$I0_18507_out0 && v$G4_7740_out0;
assign v$_12080_out0 = v$AD1_1840_out0[0:0];
assign v$_12080_out1 = v$AD1_1840_out0[1:1];
assign v$_12081_out0 = v$AD1_1841_out0[0:0];
assign v$_12081_out1 = v$AD1_1841_out0[1:1];
assign v$G1_13546_out0 = v$I2_14493_out0 && v$G2_7777_out0;
assign v$G1_13547_out0 = v$I2_14494_out0 && v$G2_7778_out0;
assign v$G7_14126_out0 = v$G8_14260_out0 && v$G6_15563_out0;
assign v$G7_14132_out0 = v$G8_14266_out0 && v$G6_15574_out0;
assign v$S_15476_out0 = v$START_3700_out0;
assign v$AD2_15661_out0 = v$AD2_9095_out0;
assign v$AD2_15662_out0 = v$AD2_9096_out0;
assign v$RAMWEN_15663_out0 = v$RAMWEN_7764_out0;
assign v$RAMWEN_15664_out0 = v$RAMWEN_7765_out0;
assign v$G8_17897_out0 = v$G3_8822_out0 && v$G2_7777_out0;
assign v$G8_17898_out0 = v$G3_8823_out0 && v$G2_7778_out0;
assign v$WENLDST_18629_out0 = v$WENLDST_12484_out0;
assign v$WENLDST_18630_out0 = v$WENLDST_12485_out0;
assign v$START_18718_out0 = v$START_3700_out0;
assign v$WENRAM_4969_out0 = v$RAMWEN_15663_out0;
assign v$WENRAM_4970_out0 = v$RAMWEN_15664_out0;
assign v$START_5492_out0 = v$START_18718_out0;
assign v$MUX1_5819_out0 = v$_12080_out0 ? v$REG1_4894_out0 : v$REG0_16254_out0;
assign v$MUX1_5820_out0 = v$_12081_out0 ? v$REG1_4895_out0 : v$REG0_16255_out0;
assign v$AD2_6401_out0 = v$AD2_15661_out0;
assign v$AD2_6402_out0 = v$AD2_15662_out0;
assign v$I2P_6433_out0 = v$G1_13546_out0;
assign v$I2P_6434_out0 = v$G1_13547_out0;
assign v$WENLDST_6687_out0 = v$WENLDST_18629_out0;
assign v$WENLDST_6688_out0 = v$WENLDST_18630_out0;
assign v$S_8018_out0 = v$S_15476_out0;
assign v$G12_9942_out0 = !(v$NEWINTERRUPT_4431_out0 || v$FF1_1376_out0);
assign v$G12_9943_out0 = !(v$NEWINTERRUPT_4432_out0 || v$FF1_1377_out0);
assign v$MUX2_10668_out0 = v$_12080_out0 ? v$REG3_11001_out0 : v$REG2_17480_out0;
assign v$MUX2_10669_out0 = v$_12081_out0 ? v$REG3_11002_out0 : v$REG2_17481_out0;
assign v$ISINTERRUPTED_11968_out0 = v$MUX1_5013_out0;
assign v$ISINTERRUPTED_11969_out0 = v$MUX1_5014_out0;
assign v$G6_12126_out0 = v$G7_10967_out0 && v$G8_17897_out0;
assign v$G6_12127_out0 = v$G7_10968_out0 && v$G8_17898_out0;
assign v$Q_14144_out0 = v$G7_14126_out0;
assign v$Q_14155_out0 = v$G7_14132_out0;
assign v$G9_15531_out0 = v$I1_4890_out0 && v$G8_17897_out0;
assign v$G9_15532_out0 = v$I1_4891_out0 && v$G8_17898_out0;
assign v$READ$REQUEST1_16828_out0 = v$READ$REQUEST_7807_out0;
assign v$READ$REQUEST0_18478_out0 = v$READ$REQUEST_7806_out0;
assign v$EXEC1_18513_out0 = v$EXEC1_3855_out0;
assign v$ININTERRUPT_1133_out0 = v$ISINTERRUPTED_11968_out0;
assign v$ININTERRUPT_1134_out0 = v$ISINTERRUPTED_11969_out0;
assign v$MUX3_1584_out0 = v$_12080_out1 ? v$MUX2_10668_out0 : v$MUX1_5819_out0;
assign v$MUX3_1585_out0 = v$_12081_out1 ? v$MUX2_10669_out0 : v$MUX1_5820_out0;
assign v$G11_2287_out0 = v$G9_15125_out0 && v$G12_9942_out0;
assign v$G11_2288_out0 = v$G9_15126_out0 && v$G12_9943_out0;
assign v$I0P_2438_out0 = v$G6_12126_out0;
assign v$I0P_2439_out0 = v$G6_12127_out0;
assign v$G11_2978_out0 = v$I2P_6433_out0 || v$I3P_13619_out0;
assign v$G11_2979_out0 = v$I2P_6434_out0 || v$I3P_13620_out0;
assign v$G2_4089_out0 = v$G24_13860_out0 && v$WENLDST_6687_out0;
assign v$G2_4090_out0 = v$G24_13861_out0 && v$WENLDST_6688_out0;
assign v$MUX8_4349_out0 = v$IR2$15_7435_out0 ? v$WENALU_4072_out0 : v$WENLDST_6687_out0;
assign v$MUX8_4350_out0 = v$IR2$15_7436_out0 ? v$WENALU_4073_out0 : v$WENLDST_6688_out0;
assign v$XOR1_5009_out0 = v$AD3_13143_out0 ^ v$AD2_6401_out0;
assign v$XOR1_5010_out0 = v$AD3_13144_out0 ^ v$AD2_6402_out0;
assign v$READ$REQUEST1_6470_out0 = v$READ$REQUEST1_16828_out0;
assign v$_7245_out0 = v$AD2_6401_out0[0:0];
assign v$_7245_out1 = v$AD2_6401_out0[1:1];
assign v$_7246_out0 = v$AD2_6402_out0[0:0];
assign v$_7246_out1 = v$AD2_6402_out0[1:1];
assign v$G2_7575_out0 = v$G1_12983_out0 || v$S_8018_out0;
assign v$EXEC1_7960_out0 = v$EXEC1_18513_out0;
assign v$EXEC1_7961_out0 = v$EXEC1_18513_out0;
assign v$EXEC1_7962_out0 = v$EXEC1_18513_out0;
assign v$EXEC1_7963_out0 = v$EXEC1_18513_out0;
assign v$EXEC1_7964_out0 = v$EXEC1_18513_out0;
assign v$EXEC1_7965_out0 = v$EXEC1_18513_out0;
assign v$EXEC1_7966_out0 = v$EXEC1_18513_out0;
assign v$EXEC1_7967_out0 = v$EXEC1_18513_out0;
assign v$EXEC1_7968_out0 = v$EXEC1_18513_out0;
assign v$EXEC1_7969_out0 = v$EXEC1_18513_out0;
assign v$EXEC1_7970_out0 = v$EXEC1_18513_out0;
assign v$READ$REQUEST0_11394_out0 = v$READ$REQUEST0_18478_out0;
assign v$I1P_14818_out0 = v$G9_15531_out0;
assign v$I1P_14819_out0 = v$G9_15532_out0;
assign v$INTERRUPTOVERFLOW_15112_out0 = v$Q_14144_out0;
assign v$INTERRUPTOVERFLOW_15113_out0 = v$Q_14155_out0;
assign v$MUX15_15925_out0 = v$START_5492_out0 ? v$IS$32$BITS_14038_out0 : v$FF1_4339_out0;
assign v$START_16352_out0 = v$START_5492_out0;
assign v$WENRAM_17082_out0 = v$WENRAM_4969_out0;
assign v$WENRAM_17083_out0 = v$WENRAM_4970_out0;
assign v$G3_0_out0 = v$G2_4089_out0 && v$IR1$VALID_18427_out0;
assign v$G3_1_out0 = v$G2_4090_out0 && v$IR1$VALID_18428_out0;
assign v$MUX4_1651_out0 = v$_7245_out0 ? v$R1_13766_out0 : v$R0_3278_out0;
assign v$MUX4_1652_out0 = v$_7246_out0 ? v$R1_13767_out0 : v$R0_3279_out0;
assign v$WENRAM_2342_out0 = v$WENRAM_17082_out0;
assign v$WENRAM_2343_out0 = v$WENRAM_17083_out0;
assign v$IS$32$BITS_2992_out0 = v$MUX15_15925_out0;
assign v$DOUT1_3157_out0 = v$MUX3_1584_out0;
assign v$DOUT1_3158_out0 = v$MUX3_1585_out0;
assign v$EQ1_3211_out0 = v$XOR1_5009_out0 == 2'h0;
assign v$EQ1_3212_out0 = v$XOR1_5010_out0 == 2'h0;
assign v$G10_3803_out0 = v$I1P_14818_out0 || v$I3P_13619_out0;
assign v$G10_3804_out0 = v$I1P_14819_out0 || v$I3P_13620_out0;
assign v$START_4238_out0 = v$START_16352_out0;
assign v$G14_5129_out0 = ! v$ININTERRUPT_1133_out0;
assign v$G14_5130_out0 = ! v$ININTERRUPT_1134_out0;
assign v$G52_7887_out0 = v$READ$REQUEST0_11394_out0 || v$FF2_13458_out0;
assign v$G44_8251_out0 = v$READ$REQUEST1_6470_out0 || v$FF1_5448_out0;
assign v$ARR1_9067_out0 = v$READ$REQUEST1_6470_out0;
assign v$ENCODED1_9520_out0 = v$G11_2978_out0;
assign v$ENCODED1_9521_out0 = v$G11_2979_out0;
assign v$G31_10793_out0 = v$NEXTINTERRUPT_18433_out0 && v$ININTERRUPT_1133_out0;
assign v$G31_10794_out0 = v$NEXTINTERRUPT_18434_out0 && v$ININTERRUPT_1134_out0;
assign v$ARR0_10978_out0 = v$READ$REQUEST0_11394_out0;
assign v$MUX5_11847_out0 = v$EQ1_18594_out0 ? v$WENFPU_3498_out0 : v$MUX8_4349_out0;
assign v$MUX5_11848_out0 = v$EQ1_18595_out0 ? v$WENFPU_3499_out0 : v$MUX8_4350_out0;
assign v$WEN_12173_out0 = v$WENRAM_17082_out0;
assign v$WEN_12174_out0 = v$WENRAM_17083_out0;
assign v$NEXTSTATE_13536_out0 = v$G2_7575_out0;
assign v$MUX5_14082_out0 = v$_7245_out0 ? v$R3_10746_out0 : v$R2_7958_out0;
assign v$MUX5_14083_out0 = v$_7246_out0 ? v$R3_10747_out0 : v$R2_7959_out0;
assign v$WEN_14218_out0 = v$WENRAM_17082_out0;
assign v$WEN_14219_out0 = v$WENRAM_17083_out0;
assign v$INTOVERFLOW_16039_out0 = v$INTERRUPTOVERFLOW_15112_out0;
assign v$INTOVERFLOW_16040_out0 = v$INTERRUPTOVERFLOW_15113_out0;
assign v$STPHALT_18124_out0 = v$G11_2287_out0;
assign v$STPHALT_18125_out0 = v$G11_2288_out0;
assign v$WENRAM1_1719_out0 = v$WENRAM_2343_out0;
assign v$RR1_1947_out0 = v$G44_8251_out0;
assign v$RD_2226_out0 = v$DOUT1_3157_out0;
assign v$RD_2227_out0 = v$DOUT1_3158_out0;
assign v$WEN_3683_out0 = v$WEN_14218_out0;
assign v$WEN_3684_out0 = v$WEN_14219_out0;
assign v$WEN_3801_out0 = v$WEN_12173_out0;
assign v$WEN_3802_out0 = v$WEN_12174_out0;
assign v$STPHALT_4317_out0 = v$STPHALT_18124_out0;
assign v$STPHALT_4318_out0 = v$STPHALT_18125_out0;
assign v$MUX6_5051_out0 = v$_7245_out1 ? v$MUX5_14082_out0 : v$MUX4_1651_out0;
assign v$MUX6_5052_out0 = v$_7246_out1 ? v$MUX5_14083_out0 : v$MUX4_1652_out0;
assign v$G29_7851_out0 = v$NEWINTERRUPT_7025_out0 || v$G31_10793_out0;
assign v$G29_7852_out0 = v$NEWINTERRUPT_7026_out0 || v$G31_10794_out0;
assign v$RR0_8089_out0 = v$G52_7887_out0;
assign v$WENRAM0_9919_out0 = v$WENRAM_2342_out0;
assign v$G33_10750_out0 = v$LDMAIN_13807_out0 || v$G14_5129_out0;
assign v$G33_10751_out0 = v$LDMAIN_13808_out0 || v$G14_5130_out0;
assign v$MUX7_10965_out0 = v$IR2$VALID$AND$NOT$FLOAD_7285_out0 ? v$MUX5_11847_out0 : v$G3_0_out0;
assign v$MUX7_10966_out0 = v$IR2$VALID$AND$NOT$FLOAD_7286_out0 ? v$MUX5_11848_out0 : v$G3_1_out0;
assign v$START_14012_out0 = v$START_4238_out0;
assign v$ENCODED0_14022_out0 = v$G10_3803_out0;
assign v$ENCODED0_14023_out0 = v$G10_3804_out0;
assign v$AD3$EQUALS$AD2_14557_out0 = v$EQ1_3211_out0;
assign v$AD3$EQUALS$AD2_14558_out0 = v$EQ1_3212_out0;
assign v$OP1_15212_out0 = v$DOUT1_3157_out0;
assign v$OP1_15213_out0 = v$DOUT1_3158_out0;
assign v$IS$32$BITS_17583_out0 = v$IS$32$BITS_2992_out0;
assign v$WEN3_3285_out0 = v$MUX7_10966_out0;
assign v$DOUT2_3513_out0 = v$MUX6_5051_out0;
assign v$DOUT2_3514_out0 = v$MUX6_5052_out0;
assign v$IS$32$BITS_4148_out0 = v$IS$32$BITS_17583_out0;
assign v$OP1_5416_out0 = v$OP1_15212_out0;
assign v$OP1_5417_out0 = v$OP1_15213_out0;
assign v$A_8693_out0 = v$RD_2226_out0;
assign v$A_8694_out0 = v$RD_2227_out0;
assign v$MUX15_9403_out0 = v$FINISHED_13867_out0 ? v$WENFPU_3498_out0 : v$MUX7_10965_out0;
assign v$RDOUT_10345_out0 = v$RD_2226_out0;
assign v$RDOUT_10346_out0 = v$RD_2227_out0;
assign v$RAMWEN1_10766_out0 = v$WENRAM1_1719_out0;
assign v$WEN_12333_out0 = v$WEN_3801_out0;
assign v$WEN_12334_out0 = v$WEN_3802_out0;
assign v$_14612_out0 = { v$ENCODED0_14022_out0,v$ENCODED1_9520_out0 };
assign v$_14613_out0 = { v$ENCODED0_14023_out0,v$ENCODED1_9521_out0 };
assign v$S_15475_out0 = v$START_14012_out0;
assign v$RAMWEN0_16569_out0 = v$WENRAM0_9919_out0;
assign v$INTERRUPTNUMBER_39_out0 = v$_14612_out0;
assign v$INTERRUPTNUMBER_40_out0 = v$_14613_out0;
assign v$AWR0_1798_out0 = v$RAMWEN0_16569_out0;
assign v$WEN3_3284_out0 = v$MUX15_9403_out0;
assign v$DATA$IN_7075_out0 = v$RDOUT_10345_out0;
assign v$DATA$IN_7076_out0 = v$RDOUT_10346_out0;
assign v$S_8017_out0 = v$S_15475_out0;
assign v$A_11042_out0 = v$A_8693_out0;
assign v$A_11043_out0 = v$A_8694_out0;
assign v$G55_13697_out0 = v$RAMWEN0_16569_out0 || v$FF3_3378_out0;
assign v$D1_14098_out0 = (v$AD3_13144_out0 == 2'b00) ? v$WEN3_3285_out0 : 1'h0;
assign v$D1_14098_out1 = (v$AD3_13144_out0 == 2'b01) ? v$WEN3_3285_out0 : 1'h0;
assign v$D1_14098_out2 = (v$AD3_13144_out0 == 2'b10) ? v$WEN3_3285_out0 : 1'h0;
assign v$D1_14098_out3 = (v$AD3_13144_out0 == 2'b11) ? v$WEN3_3285_out0 : 1'h0;
assign v$AWR1_15889_out0 = v$RAMWEN1_10766_out0;
assign v$RM_16193_out0 = v$DOUT2_3513_out0;
assign v$RM_16194_out0 = v$DOUT2_3514_out0;
assign v$A_16420_out0 = v$OP1_5416_out0;
assign v$A_16421_out0 = v$OP1_5417_out0;
assign v$G56_17676_out0 = v$RAMWEN1_10766_out0 || v$FF4_13548_out0;
assign v$WEN_18392_out0 = v$WEN_12333_out0;
assign v$WEN_18393_out0 = v$WEN_12334_out0;
assign v$RM_18596_out0 = v$DOUT2_3513_out0;
assign v$RM_18597_out0 = v$DOUT2_3514_out0;
assign v$WR1_303_out0 = v$G56_17676_out0;
assign v$G6_668_out0 = ! v$WEN_18392_out0;
assign v$G6_669_out0 = ! v$WEN_18393_out0;
assign v$G84_1235_out0 = v$AWR1_15889_out0 || v$ARR1_9067_out0;
assign v$NINTERRUPT_1595_out0 = v$INTERRUPTNUMBER_39_out0;
assign v$NINTERRUPT_1596_out0 = v$INTERRUPTNUMBER_40_out0;
assign v$DATA$IN_1607_out0 = v$DATA$IN_7075_out0;
assign v$DATA$IN_1608_out0 = v$DATA$IN_7076_out0;
assign v$MUX1_1811_out0 = v$C_6062_out0 ? v$_12228_out0 : v$RM_16193_out0;
assign v$MUX1_1812_out0 = v$C_6063_out0 ? v$_12229_out0 : v$RM_16194_out0;
assign v$A_2547_out0 = v$A_16420_out0;
assign v$A_2548_out0 = v$A_16421_out0;
assign v$MUX13_2549_out0 = v$B$IS$RD_14084_out0 ? v$RD_2226_out0 : v$RM_18596_out0;
assign v$MUX13_2550_out0 = v$B$IS$RD_14085_out0 ? v$RD_2227_out0 : v$RM_18597_out0;
assign v$A_4196_out0 = v$A_11042_out0;
assign v$A_4197_out0 = v$A_11043_out0;
assign v$RAMDIN_7038_out0 = v$DATA$IN_7075_out0;
assign v$RAMDIN_7039_out0 = v$DATA$IN_7076_out0;
assign v$G88_7401_out0 = v$ARR0_10978_out0 || v$AWR0_1798_out0;
assign v$G2_7574_out0 = v$G1_12982_out0 || v$S_8017_out0;
assign v$RM_10242_out0 = v$RM_18596_out0;
assign v$RM_10243_out0 = v$RM_18597_out0;
assign v$G8_13403_out0 = ! v$WEN_18392_out0;
assign v$G8_13404_out0 = ! v$WEN_18393_out0;
assign v$DATA_14086_out0 = v$DATA$IN_7075_out0;
assign v$DATA_14087_out0 = v$DATA$IN_7076_out0;
assign v$D1_14097_out0 = (v$AD3_13143_out0 == 2'b00) ? v$WEN3_3284_out0 : 1'h0;
assign v$D1_14097_out1 = (v$AD3_13143_out0 == 2'b01) ? v$WEN3_3284_out0 : 1'h0;
assign v$D1_14097_out2 = (v$AD3_13143_out0 == 2'b10) ? v$WEN3_3284_out0 : 1'h0;
assign v$D1_14097_out3 = (v$AD3_13143_out0 == 2'b11) ? v$WEN3_3284_out0 : 1'h0;
assign v$WR0_14268_out0 = v$G55_13697_out0;
assign v$A_18293_out0 = v$A_11042_out0;
assign v$A_18294_out0 = v$A_11043_out0;
assign v$IN_193_out0 = v$MUX1_1811_out0;
assign v$IN_194_out0 = v$MUX1_1812_out0;
assign v$_683_out0 = v$A_2547_out0[7:4];
assign v$_684_out0 = v$A_2548_out0[7:4];
assign v$WR0_1316_out0 = v$WR0_14268_out0;
assign v$DIN_1803_out0 = v$RAMDIN_7038_out0;
assign v$DIN_1804_out0 = v$RAMDIN_7039_out0;
assign v$_1852_out0 = { v$A$SAVED_9967_out0,v$A_4196_out0 };
assign v$A_3242_out0 = v$A_18293_out0;
assign v$A_3243_out0 = v$A_18294_out0;
assign v$_3799_out0 = v$A_2547_out0[15:12];
assign v$_3800_out0 = v$A_2548_out0[15:12];
assign v$_4164_out0 = v$A_2547_out0[3:0];
assign v$_4165_out0 = v$A_2548_out0[3:0];
assign v$DATA_4354_out0 = v$DATA_14086_out0;
assign v$DATA_4355_out0 = v$DATA_14087_out0;
assign v$_8691_out0 = v$A_2547_out0[11:8];
assign v$_8692_out0 = v$A_2548_out0[11:8];
assign v$SEL2_9428_out0 = v$NINTERRUPT_1595_out0[0:0];
assign v$SEL2_9429_out0 = v$NINTERRUPT_1596_out0[0:0];
assign v$DATA$IN0_10404_out0 = v$DATA$IN_1607_out0;
assign v$G79_12737_out0 = v$RR0_8089_out0 || v$WR0_14268_out0;
assign v$NEXTSTATE_13535_out0 = v$G2_7574_out0;
assign v$B_14066_out0 = v$MUX13_2549_out0;
assign v$B_14067_out0 = v$MUX13_2550_out0;
assign v$WR1_14336_out0 = v$WR1_303_out0;
assign v$DATA$IN1_15283_out0 = v$DATA$IN_1608_out0;
assign v$A_16090_out0 = v$A_4197_out0;
assign v$G36_16700_out0 = v$RR1_1947_out0 || v$WR1_303_out0;
assign v$SEL3_17400_out0 = v$NINTERRUPT_1595_out0[1:1];
assign v$SEL3_17401_out0 = v$NINTERRUPT_1596_out0[1:1];
assign v$RM_18197_out0 = v$RM_10242_out0;
assign v$RM_18198_out0 = v$RM_10243_out0;
assign v$SEL5_313_out0 = v$A_3242_out0[15:15];
assign v$SEL5_314_out0 = v$A_3243_out0[15:15];
assign v$MUX7_1135_out0 = v$SEL2_9428_out0 ? v$INT3_271_out0 : v$INT2_256_out0;
assign v$MUX7_1136_out0 = v$SEL2_9429_out0 ? v$INT3_272_out0 : v$INT2_257_out0;
assign v$_1853_out0 = { v$A$SAVED_9968_out0,v$A_16090_out0 };
assign v$R0_2000_out0 = v$G79_12737_out0;
assign v$PIN_2935_out0 = v$DIN_1803_out0;
assign v$PIN_2936_out0 = v$DIN_1804_out0;
assign v$B_3366_out0 = v$B_14066_out0;
assign v$B_3367_out0 = v$B_14067_out0;
assign v$_3701_out0 = v$_683_out0[1:0];
assign v$_3701_out1 = v$_683_out0[3:2];
assign v$_3702_out0 = v$_684_out0[1:0];
assign v$_3702_out1 = v$_684_out0[3:2];
assign v$SEL1_3721_out0 = v$A_16090_out0[15:15];
assign v$IN_4360_out0 = v$IN_193_out0;
assign v$IN_4364_out0 = v$IN_194_out0;
assign v$A_9404_out0 = v$RM_18197_out0;
assign v$A_9405_out0 = v$RM_18198_out0;
assign v$DATAIN1_9634_out0 = v$DATA$IN1_15283_out0;
assign v$SEL9_9969_out0 = v$A_3242_out0[9:0];
assign v$SEL9_9970_out0 = v$A_3243_out0[9:0];
assign v$MUX13_10727_out0 = v$START_5492_out0 ? v$_1852_out0 : v$REG2_4047_out0;
assign v$DATAIN0_11058_out0 = v$DATA$IN0_10404_out0;
assign v$SEL4_11854_out0 = v$DATA_4354_out0[7:0];
assign v$SEL4_11855_out0 = v$DATA_4355_out0[7:0];
assign v$SEL1_11971_out0 = v$DATA_4354_out0[11:0];
assign v$SEL1_11972_out0 = v$DATA_4355_out0[11:0];
assign v$SEL7_12477_out0 = v$A_16090_out0[9:0];
assign v$_13256_out0 = v$_8691_out0[1:0];
assign v$_13256_out1 = v$_8691_out0[3:2];
assign v$_13257_out0 = v$_8692_out0[1:0];
assign v$_13257_out1 = v$_8692_out0[3:2];
assign v$A_13811_out0 = v$A_3242_out0;
assign v$A_13815_out0 = v$A_16090_out0;
assign v$A_13817_out0 = v$A_3243_out0;
assign v$MUX6_14420_out0 = v$SEL2_9428_out0 ? v$INT1_18533_out0 : v$INT0_15885_out0;
assign v$MUX6_14421_out0 = v$SEL2_9429_out0 ? v$INT1_18534_out0 : v$INT0_15886_out0;
assign v$_15018_out0 = v$_4164_out0[1:0];
assign v$_15018_out1 = v$_4164_out0[3:2];
assign v$_15019_out0 = v$_4165_out0[1:0];
assign v$_15019_out1 = v$_4165_out0[3:2];
assign v$THRESHOLD_15533_out0 = v$DATA_4354_out0;
assign v$THRESHOLD_15534_out0 = v$DATA_4355_out0;
assign v$SEL11_15556_out0 = v$A_3242_out0[15:15];
assign v$SEL11_15557_out0 = v$A_3243_out0[15:15];
assign v$_15826_out0 = { v$A$SAVED_14631_out0,v$A_3242_out0 };
assign v$_15827_out0 = { v$A$SAVED_14632_out0,v$A_3243_out0 };
assign v$_16231_out0 = v$_3799_out0[1:0];
assign v$_16231_out1 = v$_3799_out0[3:2];
assign v$_16232_out0 = v$_3800_out0[1:0];
assign v$_16232_out1 = v$_3800_out0[3:2];
assign v$SEL13_17581_out0 = v$A_3242_out0[15:15];
assign v$SEL13_17582_out0 = v$A_3243_out0[15:15];
assign v$R1_17899_out0 = v$G36_16700_out0;
assign v$SEL1_18247_out0 = v$DIN_1803_out0[3:0];
assign v$SEL1_18248_out0 = v$DIN_1804_out0[3:0];
assign v$MODE_48_out0 = v$SEL4_11854_out0;
assign v$MODE_49_out0 = v$SEL4_11855_out0;
assign v$_330_out0 = v$_13256_out0[0:0];
assign v$_330_out1 = v$_13256_out0[1:1];
assign v$_331_out0 = v$_13257_out0[0:0];
assign v$_331_out1 = v$_13257_out0[1:1];
assign v$SEL12_1192_out0 = v$MUX13_10727_out0[31:16];
assign v$_1686_out0 = { v$C6_1536_out0,v$SEL7_12477_out0 };
assign v$_2231_out0 = { v$C8_8206_out0,v$SEL9_9969_out0 };
assign v$_2232_out0 = { v$C8_8207_out0,v$SEL9_9970_out0 };
assign v$G59_2571_out0 = v$PHALT_15137_out0 && v$R1_17899_out0;
assign v$A$32BIT_2990_out0 = v$_15826_out0;
assign v$A$32BIT_2991_out0 = v$_15827_out0;
assign v$_3118_out0 = v$_16231_out1[0:0];
assign v$_3118_out1 = v$_16231_out1[1:1];
assign v$_3119_out0 = v$_16232_out1[0:0];
assign v$_3119_out1 = v$_16232_out1[1:1];
assign v$MUX4_3842_out0 = v$G68_14822_out0 ? v$REG10_16463_out0 : v$DATAIN0_11058_out0;
assign v$_4019_out0 = v$_3701_out0[0:0];
assign v$_4019_out1 = v$_3701_out0[1:1];
assign v$_4020_out0 = v$_3702_out0[0:0];
assign v$_4020_out1 = v$_3702_out0[1:1];
assign v$_4892_out0 = v$_13256_out1[0:0];
assign v$_4892_out1 = v$_13256_out1[1:1];
assign v$_4893_out0 = v$_13257_out1[0:0];
assign v$_4893_out1 = v$_13257_out1[1:1];
assign v$_5405_out0 = v$_15018_out1[0:0];
assign v$_5405_out1 = v$_15018_out1[1:1];
assign v$_5406_out0 = v$_15019_out1[0:0];
assign v$_5406_out1 = v$_15019_out1[1:1];
assign {v$A1_6409_out1,v$A1_6409_out0 } = v$XOR1_5078_out0 + v$A_9404_out0 + v$SUBEN_12858_out0;
assign {v$A1_6410_out1,v$A1_6410_out0 } = v$XOR1_5079_out0 + v$A_9405_out0 + v$SUBEN_12859_out0;
assign v$R0_6676_out0 = v$R0_2000_out0;
assign v$SEL1_7529_out0 = v$A_13811_out0[14:10];
assign v$SEL1_7533_out0 = v$A_13815_out0[14:10];
assign v$SEL1_7535_out0 = v$A_13817_out0[14:10];
assign v$_7902_out0 = v$PIN_2935_out0[7:0];
assign v$_7902_out1 = v$PIN_2935_out0[15:8];
assign v$_7903_out0 = v$PIN_2936_out0[7:0];
assign v$_7903_out1 = v$PIN_2936_out0[15:8];
assign v$IN_9566_out0 = v$IN_4360_out0;
assign v$IN_9570_out0 = v$IN_4364_out0;
assign v$_10244_out0 = v$_3701_out1[0:0];
assign v$_10244_out1 = v$_3701_out1[1:1];
assign v$_10245_out0 = v$_3702_out1[0:0];
assign v$_10245_out1 = v$_3702_out1[1:1];
assign v$MUX5_10896_out0 = v$G69_15812_out0 ? v$REG11_9622_out0 : v$DATAIN1_9634_out0;
assign v$_11056_out0 = v$_15018_out0[0:0];
assign v$_11056_out1 = v$_15018_out0[1:1];
assign v$_11057_out0 = v$_15019_out0[0:0];
assign v$_11057_out1 = v$_15019_out0[1:1];
assign v$R1_11886_out0 = v$R1_17899_out0;
assign v$G1_15142_out0 = ! v$SEL5_313_out0;
assign v$G1_15143_out0 = ! v$SEL5_314_out0;
assign v$_16550_out0 = v$_16231_out0[0:0];
assign v$_16550_out1 = v$_16231_out0[1:1];
assign v$_16551_out0 = v$_16232_out0[0:0];
assign v$_16551_out1 = v$_16232_out0[1:1];
assign v$A$32$BIT_16831_out0 = v$MUX13_10727_out0;
assign v$MUX5_16988_out0 = v$SEL3_17400_out0 ? v$MUX7_1135_out0 : v$MUX6_14420_out0;
assign v$MUX5_16989_out0 = v$SEL3_17401_out0 ? v$MUX7_1136_out0 : v$MUX6_14421_out0;
assign v$B_17051_out0 = v$B_3366_out0;
assign v$B_17052_out0 = v$B_3367_out0;
assign v$B_18099_out0 = v$B_3366_out0;
assign v$B_18100_out0 = v$B_3367_out0;
assign v$A$32$BIT_18440_out0 = v$_1853_out0;
assign v$A$EXP_284_out0 = v$SEL1_7529_out0;
assign v$A$EXP_288_out0 = v$SEL1_7533_out0;
assign v$A$EXP_290_out0 = v$SEL1_7535_out0;
assign v$_1197_out0 = v$IN_9566_out0[0:0];
assign v$_1198_out0 = v$IN_9570_out0[0:0];
assign v$A_2293_out0 = v$SEL12_1192_out0;
assign v$G6_3503_out0 = v$R0_6676_out0 && v$R1_11886_out0;
assign v$_4800_out0 = v$IN_9566_out0[14:0];
assign v$_4804_out0 = v$IN_9570_out0[14:0];
assign v$SEL2_6165_out0 = v$B_17051_out0[14:0];
assign v$SEL2_6166_out0 = v$B_17052_out0[14:0];
assign v$_7418_out0 = { v$_2231_out0,v$C2_1171_out0 };
assign v$_7419_out0 = { v$_2232_out0,v$C2_1172_out0 };
assign v$8LSB_7606_out0 = v$_7902_out0;
assign v$8LSB_7607_out0 = v$_7903_out0;
assign v$COUT_8292_out0 = v$A1_6409_out1;
assign v$COUT_8293_out0 = v$A1_6410_out1;
assign v$SUM_10304_out0 = v$A1_6409_out0;
assign v$SUM_10305_out0 = v$A1_6410_out0;
assign v$_10416_out0 = v$IN_9566_out0[15:15];
assign v$_10417_out0 = v$IN_9570_out0[15:15];
assign v$EQ1_11626_out0 = v$A$32$BIT_16831_out0 == 32'h0;
assign v$EQ1_11627_out0 = v$A$32$BIT_18440_out0 == 32'h0;
assign v$G62_11967_out0 = v$G59_2571_out0 && v$PCHALT_16563_out0;
assign v$B_12138_out0 = v$B_18100_out0;
assign v$_12523_out0 = { v$B$SAVED_3884_out0,v$B_18099_out0 };
assign v$END_12712_out0 = v$_7902_out1;
assign v$END_12713_out0 = v$_7903_out1;
assign v$SEL4_12976_out0 = v$A$32BIT_2990_out0[22:0];
assign v$SEL4_12977_out0 = v$A$32BIT_2991_out0[22:0];
assign v$_13269_out0 = v$IN_9566_out0[0:0];
assign v$_13272_out0 = v$IN_9570_out0[0:0];
assign v$A_13812_out0 = v$A$32BIT_2990_out0;
assign v$A_13814_out0 = v$A$32$BIT_16831_out0;
assign v$A_13816_out0 = v$A$32$BIT_18440_out0;
assign v$A_13818_out0 = v$A$32BIT_2991_out0;
assign v$EQ3_14302_out0 = v$A$32$BIT_16831_out0 == 32'h0;
assign v$EQ3_14303_out0 = v$A$32$BIT_18440_out0 == 32'h0;
assign v$SEL6_14456_out0 = v$B_17051_out0[15:15];
assign v$SEL6_14457_out0 = v$B_17052_out0[15:15];
assign v$_14599_out0 = v$IN_9566_out0[15:1];
assign v$_14603_out0 = v$IN_9570_out0[15:1];
assign v$_14633_out0 = v$IN_9566_out0[15:1];
assign v$_14637_out0 = v$IN_9570_out0[15:1];
assign v$_16747_out0 = v$IN_9566_out0[15:1];
assign v$_16751_out0 = v$IN_9570_out0[15:1];
assign v$SEL8_17494_out0 = v$A$32$BIT_16831_out0[22:0];
assign v$SEL8_17495_out0 = v$A$32$BIT_18440_out0[22:0];
assign v$MODE_17842_out0 = v$MODE_48_out0;
assign v$MODE_17843_out0 = v$MODE_49_out0;
assign v$MUX14_1189_out0 = v$START_5492_out0 ? v$_12523_out0 : v$REG1_7848_out0;
assign v$_1477_out0 = { v$C1_7971_out0,v$_4800_out0 };
assign v$_1481_out0 = { v$C1_7975_out0,v$_4804_out0 };
assign v$SEL1_3720_out0 = v$A_2293_out0[15:15];
assign v$G3_3950_out0 = ! v$SEL6_14456_out0;
assign v$G3_3951_out0 = ! v$SEL6_14457_out0;
assign v$B_4829_out0 = v$B_12138_out0;
assign v$RMN_6155_out0 = v$SUM_10304_out0;
assign v$RMN_6156_out0 = v$SUM_10305_out0;
assign v$MUX8_7078_out0 = v$IS$32$BITS_1282_out0 ? v$SEL8_17495_out0 : v$_1686_out0;
assign v$SEL1_7530_out0 = v$A_13812_out0[30:23];
assign v$SEL1_7532_out0 = v$A_13814_out0[30:23];
assign v$SEL1_7534_out0 = v$A_13816_out0[30:23];
assign v$SEL1_7536_out0 = v$A_13818_out0[30:23];
assign v$SEL5_7813_out0 = v$B_12138_out0[9:0];
assign v$_8213_out0 = v$8LSB_7606_out0[3:0];
assign v$_8213_out1 = v$8LSB_7606_out0[7:4];
assign v$_8214_out0 = v$8LSB_7607_out0[3:0];
assign v$_8214_out1 = v$8LSB_7607_out0[7:4];
assign v$_9445_out0 = { v$_16747_out0,v$LSB_7815_out0 };
assign v$_9449_out0 = { v$_16751_out0,v$LSB_7816_out0 };
assign v$MODE_10801_out0 = v$MODE_17842_out0;
assign v$MODE_10802_out0 = v$MODE_17843_out0;
assign v$A_11324_out0 = v$A$EXP_284_out0;
assign v$A_11332_out0 = v$A$EXP_288_out0;
assign v$A_11344_out0 = v$A$EXP_290_out0;
assign v$SEL7_12476_out0 = v$A_2293_out0[9:0];
assign v$_12524_out0 = { v$B$SAVED_3885_out0,v$B_12138_out0 };
assign v$HALTVALID_13286_out0 = v$G6_3503_out0;
assign v$_13304_out0 = { v$_14599_out0,v$_13269_out0 };
assign v$_13308_out0 = { v$_14603_out0,v$_13272_out0 };
assign v$SEL2_13434_out0 = v$B_12138_out0[15:15];
assign v$MUX6_13737_out0 = v$S$FF_10816_out0 ? v$LSB_7815_out0 : v$_10416_out0;
assign v$MUX6_13738_out0 = v$S$FF_10817_out0 ? v$LSB_7816_out0 : v$_10417_out0;
assign v$A_13813_out0 = v$A_2293_out0;
assign v$DM1_16244_out0 = v$HALTSEL_14742_out0 ? 1'h0 : v$G6_3503_out0;
assign v$DM1_16244_out1 = v$HALTSEL_14742_out0 ? v$G6_3503_out0 : 1'h0;
assign v$HALT_16371_out0 = v$G6_3503_out0;
assign v$MUX5_17066_out0 = v$S_10699_out0 ? v$_1197_out0 : v$C2_2666_out0;
assign v$MUX5_17067_out0 = v$S_10700_out0 ? v$_1198_out0 : v$C2_2667_out0;
assign v$_17770_out0 = { v$SEL4_12976_out0,v$C3_5386_out0 };
assign v$_17771_out0 = { v$SEL4_12977_out0,v$C3_5387_out0 };
assign v$A$EXP_285_out0 = v$SEL1_7530_out0;
assign v$A$EXP_287_out0 = v$SEL1_7532_out0;
assign v$A$EXP_289_out0 = v$SEL1_7534_out0;
assign v$A$EXP_291_out0 = v$SEL1_7536_out0;
assign v$_1685_out0 = { v$C6_1535_out0,v$SEL7_12476_out0 };
assign v$_1696_out0 = v$_8213_out0[1:0];
assign v$_1696_out1 = v$_8213_out0[3:2];
assign v$_1697_out0 = v$_8214_out0[1:0];
assign v$_1697_out1 = v$_8214_out0[3:2];
assign v$B$32$BIT_1896_out0 = v$_12524_out0;
assign v$MUX1_2603_out0 = v$G15_18535_out0 ? v$RMN_6155_out0 : v$RM_18197_out0;
assign v$MUX1_2604_out0 = v$G15_18536_out0 ? v$RMN_6156_out0 : v$RM_18198_out0;
assign v$SEL11_3703_out0 = v$MUX14_1189_out0[31:16];
assign v$MUX8_5397_out0 = v$IS$32$BIT_10862_out0 ? v$_17770_out0 : v$_7418_out0;
assign v$MUX8_5398_out0 = v$IS$32$BIT_10863_out0 ? v$_17771_out0 : v$_7419_out0;
assign v$SEL2_6972_out0 = v$B_4829_out0[14:10];
assign v$HALT1_7229_out0 = v$DM1_16244_out1;
assign v$SEL4_7340_out0 = v$A_11324_out0[1:1];
assign v$SEL4_7346_out0 = v$A_11332_out0[1:1];
assign v$SEL4_7355_out0 = v$A_11344_out0[1:1];
assign v$SEL1_7531_out0 = v$A_13813_out0[14:10];
assign v$HALTVALID_7744_out0 = v$HALTVALID_13286_out0;
assign v$SEL3_8430_out0 = v$A_11324_out0[2:2];
assign v$SEL3_8436_out0 = v$A_11332_out0[2:2];
assign v$SEL3_8445_out0 = v$A_11344_out0[2:2];
assign v$G7_9875_out0 = ! v$DM1_16244_out0;
assign v$HALT0_11685_out0 = v$DM1_16244_out0;
assign v$_11808_out0 = { v$_14633_out0,v$MUX6_13737_out0 };
assign v$_11812_out0 = { v$_14637_out0,v$MUX6_13738_out0 };
assign v$A$MANTISA_11826_out0 = v$MUX8_7078_out0;
assign v$SEL5_12782_out0 = v$A_11324_out0[0:0];
assign v$SEL5_12788_out0 = v$A_11332_out0[0:0];
assign v$SEL5_12797_out0 = v$A_11344_out0[0:0];
assign v$_13151_out0 = v$_8213_out1[1:0];
assign v$_13151_out1 = v$_8213_out1[3:2];
assign v$_13152_out0 = v$_8214_out1[1:0];
assign v$_13152_out1 = v$_8214_out1[3:2];
assign v$MUX4_15990_out0 = v$EN_16965_out0 ? v$_1477_out0 : v$IN_9566_out0;
assign v$MUX4_15994_out0 = v$EN_16969_out0 ? v$_1481_out0 : v$IN_9570_out0;
assign v$MUX10_16397_out0 = v$EQ1_16219_out0 ? v$G3_3950_out0 : v$SEL6_14456_out0;
assign v$MUX10_16398_out0 = v$EQ1_16220_out0 ? v$G3_3951_out0 : v$SEL6_14457_out0;
assign v$SEL2_16606_out0 = v$A_11324_out0[3:3];
assign v$SEL2_16612_out0 = v$A_11332_out0[3:3];
assign v$SEL2_16621_out0 = v$A_11344_out0[3:3];
assign v$B$32$BIT_17689_out0 = v$MUX14_1189_out0;
assign v$G1_17888_out0 = ((v$SEL1_3721_out0 && !v$SEL2_13434_out0) || (!v$SEL1_3721_out0) && v$SEL2_13434_out0);
assign v$SEL1_18044_out0 = v$A_11324_out0[4:4];
assign v$SEL1_18046_out0 = v$A_11332_out0[4:4];
assign v$SEL1_18047_out0 = v$A_11344_out0[4:4];
assign v$_18089_out0 = { v$C7_6038_out0,v$SEL5_7813_out0 };
assign v$A$EXP_286_out0 = v$SEL1_7531_out0;
assign v$HALT0_361_out0 = v$HALT0_11685_out0;
assign v$_1494_out0 = { v$SEL2_6165_out0,v$MUX10_16397_out0 };
assign v$_1495_out0 = { v$SEL2_6166_out0,v$MUX10_16398_out0 };
assign v$A0_1731_out0 = v$SEL5_12782_out0;
assign v$A0_1737_out0 = v$SEL5_12788_out0;
assign v$A0_1746_out0 = v$SEL5_12797_out0;
assign v$EQ4_3006_out0 = v$B$32$BIT_17689_out0 == 32'h0;
assign v$EQ4_3007_out0 = v$B$32$BIT_1896_out0 == 32'h0;
assign v$_3486_out0 = v$_1696_out0[0:0];
assign v$_3486_out1 = v$_1696_out0[1:1];
assign v$_3487_out0 = v$_1697_out0[0:0];
assign v$_3487_out1 = v$_1697_out0[1:1];
assign v$A$MANTISA_3756_out0 = v$MUX8_5397_out0;
assign v$A$MANTISA_3757_out0 = v$MUX8_5398_out0;
assign v$HALT1_4159_out0 = v$HALT1_7229_out0;
assign v$SEL6_4441_out0 = v$B$32$BIT_17689_out0[22:0];
assign v$SEL6_4442_out0 = v$B$32$BIT_1896_out0[22:0];
assign v$B_4828_out0 = v$B$32$BIT_17689_out0;
assign v$B_4830_out0 = v$B$32$BIT_1896_out0;
assign v$B_6548_out0 = v$SEL11_3703_out0;
assign v$MUX8_7077_out0 = v$IS$32$BITS_2992_out0 ? v$SEL8_17494_out0 : v$_1685_out0;
assign v$A2_8063_out0 = v$SEL3_8430_out0;
assign v$A2_8069_out0 = v$SEL3_8436_out0;
assign v$A2_8078_out0 = v$SEL3_8445_out0;
assign v$_8090_out0 = v$_13151_out0[0:0];
assign v$_8090_out1 = v$_13151_out0[1:1];
assign v$_8091_out0 = v$_13152_out0[0:0];
assign v$_8091_out1 = v$_13152_out0[1:1];
assign v$_9372_out0 = v$_13151_out1[0:0];
assign v$_9372_out1 = v$_13151_out1[1:1];
assign v$_9373_out0 = v$_13152_out1[0:0];
assign v$_9373_out1 = v$_13152_out1[1:1];
assign v$A3_10708_out0 = v$SEL2_16606_out0;
assign v$A3_10714_out0 = v$SEL2_16612_out0;
assign v$A3_10723_out0 = v$SEL2_16621_out0;
assign v$A_11325_out0 = v$A$EXP_285_out0;
assign v$A_11329_out0 = v$A$EXP_287_out0;
assign v$A_11333_out0 = v$A$EXP_289_out0;
assign v$A_11345_out0 = v$A$EXP_291_out0;
assign v$MUX2_12038_out0 = v$G3_2605_out0 ? v$_9445_out0 : v$MUX4_15990_out0;
assign v$MUX2_12042_out0 = v$G3_2609_out0 ? v$_9449_out0 : v$MUX4_15994_out0;
assign v$SIGN_12761_out0 = v$G1_17888_out0;
assign v$_14024_out0 = v$MUX1_2603_out0[11:0];
assign v$_14024_out1 = v$MUX1_2603_out0[15:4];
assign v$_14025_out0 = v$MUX1_2604_out0[11:0];
assign v$_14025_out1 = v$MUX1_2604_out0[15:4];
assign v$_14078_out0 = v$_1696_out1[0:0];
assign v$_14078_out1 = v$_1696_out1[1:1];
assign v$_14079_out0 = v$_1697_out1[0:0];
assign v$_14079_out1 = v$_1697_out1[1:1];
assign v$A1_14345_out0 = v$SEL4_7340_out0;
assign v$A1_14351_out0 = v$SEL4_7346_out0;
assign v$A1_14360_out0 = v$SEL4_7355_out0;
assign v$A4_15007_out0 = v$SEL1_18044_out0;
assign v$A4_15009_out0 = v$SEL1_18046_out0;
assign v$A4_15010_out0 = v$SEL1_18047_out0;
assign v$G8_15731_out0 = v$G7_9875_out0 && v$DM1_16244_out1;
assign v$EQ2_16156_out0 = v$B$32$BIT_17689_out0 == 32'h0;
assign v$EQ2_16157_out0 = v$B$32$BIT_1896_out0 == 32'h0;
assign v$B$EXP_16676_out0 = v$SEL2_6972_out0;
assign v$A$MANTISA_17916_out0 = v$A$MANTISA_11826_out0;
assign v$SIGN_1368_out0 = v$SIGN_12761_out0;
assign v$SIGN_1369_out0 = v$SIGN_12761_out0;
assign v$HALT1_3104_out0 = v$HALT1_4159_out0;
assign v$B_4827_out0 = v$B_6548_out0;
assign v$HALT0_5804_out0 = v$HALT0_361_out0;
assign v$G72_5901_out0 = ! v$HALT0_361_out0;
assign v$G5_6198_out0 = v$EQ3_14302_out0 || v$EQ4_3006_out0;
assign v$G5_6199_out0 = v$EQ3_14303_out0 || v$EQ4_3007_out0;
assign v$MUX1_6677_out0 = v$G4_4029_out0 ? v$_11808_out0 : v$MUX2_12038_out0;
assign v$MUX1_6681_out0 = v$G4_4033_out0 ? v$_11812_out0 : v$MUX2_12042_out0;
assign v$SEL2_6971_out0 = v$B_4828_out0[30:23];
assign v$SEL2_6973_out0 = v$B_4830_out0[30:23];
assign v$G78_7096_out0 = ! v$HALT1_4159_out0;
assign v$SEL5_7812_out0 = v$B_6548_out0[9:0];
assign v$SEL1_10292_out0 = v$A_11325_out0[3:0];
assign v$SEL1_10293_out0 = v$A_11329_out0[3:0];
assign v$SEL1_10294_out0 = v$A_11333_out0[3:0];
assign v$SEL1_10297_out0 = v$A_11345_out0[3:0];
assign v$A_11328_out0 = v$A$EXP_286_out0;
assign v$A$MANTISA_11825_out0 = v$MUX8_7077_out0;
assign v$MUX7_12743_out0 = v$IS$32$BITS_1282_out0 ? v$SEL6_4442_out0 : v$_18089_out0;
assign v$A$MANTISSA_13185_out0 = v$A$MANTISA_3756_out0;
assign v$A$MANTISSA_13186_out0 = v$A$MANTISA_3757_out0;
assign v$G54_13285_out0 = v$RAMWEN1_10766_out0 && v$HALT1_4159_out0;
assign v$G50_13303_out0 = ! v$HALT1_4159_out0;
assign v$SEL2_13433_out0 = v$B_6548_out0[15:15];
assign v$G63_13677_out0 = v$HALT0_361_out0 || v$HALT1_4159_out0;
assign v$HALT0_14137_out0 = v$HALT0_361_out0;
assign v$RAMADDRMUX_14376_out0 = v$_14024_out0;
assign v$RAMADDRMUX_14377_out0 = v$_14025_out0;
assign v$B_14440_out0 = v$B$EXP_16676_out0;
assign v$A$MANTISA_14550_out0 = v$A$MANTISA_17916_out0;
assign v$ADDRMSB_15028_out0 = v$_14024_out1;
assign v$ADDRMSB_15029_out0 = v$_14025_out1;
assign v$G45_15360_out0 = v$READ$REQUEST1_6470_out0 && v$HALT1_4159_out0;
assign v$G3_16009_out0 = v$EQ1_11626_out0 || v$EQ2_16156_out0;
assign v$G3_16010_out0 = v$EQ1_11627_out0 || v$EQ2_16157_out0;
assign v$SEL4_17332_out0 = v$A_11325_out0[7:4];
assign v$SEL4_17333_out0 = v$A_11329_out0[7:4];
assign v$SEL4_17334_out0 = v$A_11333_out0[7:4];
assign v$SEL4_17337_out0 = v$A_11345_out0[7:4];
assign v$G53_17493_out0 = v$RAMWEN0_16569_out0 && v$HALT0_361_out0;
assign v$B_17746_out0 = v$_1494_out0;
assign v$B_17747_out0 = v$_1495_out0;
assign v$HALT1_18308_out0 = v$HALT1_4159_out0;
assign v$G51_18762_out0 = v$READ$REQUEST0_11394_out0 && v$HALT0_361_out0;
assign v$SEL12_16_out0 = v$B_17746_out0[9:0];
assign v$SEL12_17_out0 = v$B_17747_out0[9:0];
assign v$SEL3_1251_out0 = v$A$MANTISSA_13185_out0[23:12];
assign v$SEL3_1252_out0 = v$A$MANTISSA_13186_out0[23:12];
assign v$HALT_1290_out0 = v$G63_13677_out0;
assign v$MUX3_1957_out0 = v$G8_1886_out0 ? v$_13304_out0 : v$MUX1_6677_out0;
assign v$MUX3_1961_out0 = v$G8_1890_out0 ? v$_13308_out0 : v$MUX1_6681_out0;
assign v$ARBHALT0_2908_out0 = v$HALT0_5804_out0;
assign v$B$MANTISA_3003_out0 = v$MUX7_12743_out0;
assign v$SEL1_3249_out0 = v$A$MANTISSA_13185_out0[11:0];
assign v$SEL1_3250_out0 = v$A$MANTISSA_13186_out0[11:0];
assign v$SEL7_4178_out0 = v$B_14440_out0[3:3];
assign v$RAMADDRMUX_4816_out0 = v$RAMADDRMUX_14376_out0;
assign v$RAMADDRMUX_4817_out0 = v$RAMADDRMUX_14377_out0;
assign v$B_4825_out0 = v$B_17746_out0;
assign v$B_4831_out0 = v$B_17747_out0;
assign v$ARBHALT1_5453_out0 = v$HALT1_3104_out0;
assign v$SEL6_5807_out0 = v$B_14440_out0[4:4];
assign v$G64_6432_out0 = v$G50_13303_out0 && v$R1_17899_out0;
assign v$SEL2_6970_out0 = v$B_4827_out0[14:10];
assign v$G1_7333_out0 = ! v$HALT1_18308_out0;
assign v$SEL4_7343_out0 = v$A_11328_out0[1:1];
assign v$G2_8130_out0 = ! v$HALT0_14137_out0;
assign v$SEL3_8433_out0 = v$A_11328_out0[2:2];
assign v$SEL9_10849_out0 = v$B_14440_out0[1:1];
assign v$A_11326_out0 = v$SEL4_17332_out0;
assign v$A_11327_out0 = v$SEL1_10292_out0;
assign v$A_11330_out0 = v$SEL4_17333_out0;
assign v$A_11331_out0 = v$SEL1_10293_out0;
assign v$A_11334_out0 = v$SEL4_17334_out0;
assign v$A_11335_out0 = v$SEL1_10294_out0;
assign v$A_11346_out0 = v$SEL4_17337_out0;
assign v$A_11347_out0 = v$SEL1_10297_out0;
assign v$SEL3_11895_out0 = v$A$MANTISA_14550_out0[22:0];
assign v$SEL10_12618_out0 = v$B_14440_out0[0:0];
assign v$SEL5_12785_out0 = v$A_11328_out0[0:0];
assign v$SEL8_12926_out0 = v$B_14440_out0[2:2];
assign v$SEL15_13612_out0 = v$B_17746_out0[15:15];
assign v$SEL15_13613_out0 = v$B_17747_out0[15:15];
assign v$G74_15740_out0 = v$REG4_10994_out0 && v$G72_5901_out0;
assign v$SEL1_15749_out0 = v$A$MANTISA_14550_out0[22:0];
assign v$SEL2_16609_out0 = v$A_11328_out0[3:3];
assign v$B$EXP_16675_out0 = v$SEL2_6971_out0;
assign v$B$EXP_16677_out0 = v$SEL2_6973_out0;
assign v$G1_17887_out0 = ((v$SEL1_3720_out0 && !v$SEL2_13433_out0) || (!v$SEL1_3720_out0) && v$SEL2_13433_out0);
assign v$A$MANTISA_17915_out0 = v$A$MANTISA_11825_out0;
assign v$SEL1_18045_out0 = v$A_11328_out0[4:4];
assign v$_18088_out0 = { v$C7_6037_out0,v$SEL5_7812_out0 };
assign v$G77_18210_out0 = v$REG7_6181_out0 && v$G78_7096_out0;
assign v$_18260_out0 = { v$B$SAVED_4358_out0,v$B_17746_out0 };
assign v$_18261_out0 = { v$B$SAVED_4359_out0,v$B_17747_out0 };
assign v$RAMADDRMUX_418_out0 = v$RAMADDRMUX_4816_out0;
assign v$RAMADDRMUX_419_out0 = v$RAMADDRMUX_4817_out0;
assign v$G83_428_out0 = v$G74_15740_out0 && v$G87_5144_out0;
assign v$A0_1734_out0 = v$SEL5_12785_out0;
assign v$A_2543_out0 = v$SEL3_1251_out0;
assign v$A_2544_out0 = v$SEL1_3249_out0;
assign v$A_2545_out0 = v$SEL3_1252_out0;
assign v$A_2546_out0 = v$SEL1_3250_out0;
assign v$G3_2977_out0 = v$G1_7333_out0 && v$WR1_14336_out0;
assign v$OUT_3176_out0 = v$MUX3_1957_out0;
assign v$OUT_3180_out0 = v$MUX3_1961_out0;
assign v$B0_3657_out0 = v$SEL10_12618_out0;
assign v$B$MANTISA_4071_out0 = v$B$MANTISA_3003_out0;
assign v$G85_6200_out0 = v$G77_18210_out0 && v$G86_13527_out0;
assign v$SEL2_6968_out0 = v$B_4825_out0[14:10];
assign v$SEL2_6974_out0 = v$B_4831_out0[14:10];
assign v$SEL4_7341_out0 = v$A_11326_out0[1:1];
assign v$SEL4_7342_out0 = v$A_11327_out0[1:1];
assign v$SEL4_7344_out0 = v$A_11330_out0[1:1];
assign v$SEL4_7345_out0 = v$A_11331_out0[1:1];
assign v$SEL4_7347_out0 = v$A_11334_out0[1:1];
assign v$SEL4_7348_out0 = v$A_11335_out0[1:1];
assign v$SEL4_7356_out0 = v$A_11346_out0[1:1];
assign v$SEL4_7357_out0 = v$A_11347_out0[1:1];
assign v$HALT_7572_out0 = v$ARBHALT0_2908_out0;
assign v$HALT_7573_out0 = v$ARBHALT1_5453_out0;
assign v$A2_8066_out0 = v$SEL3_8433_out0;
assign v$SEL3_8431_out0 = v$A_11326_out0[2:2];
assign v$SEL3_8432_out0 = v$A_11327_out0[2:2];
assign v$SEL3_8434_out0 = v$A_11330_out0[2:2];
assign v$SEL3_8435_out0 = v$A_11331_out0[2:2];
assign v$SEL3_8437_out0 = v$A_11334_out0[2:2];
assign v$SEL3_8438_out0 = v$A_11335_out0[2:2];
assign v$SEL3_8446_out0 = v$A_11346_out0[2:2];
assign v$SEL3_8447_out0 = v$A_11347_out0[2:2];
assign v$A3_10711_out0 = v$SEL2_16609_out0;
assign v$MUX7_12742_out0 = v$IS$32$BITS_2992_out0 ? v$SEL6_4441_out0 : v$_18088_out0;
assign v$SIGN_12760_out0 = v$G1_17887_out0;
assign v$SEL5_12783_out0 = v$A_11326_out0[0:0];
assign v$SEL5_12784_out0 = v$A_11327_out0[0:0];
assign v$SEL5_12786_out0 = v$A_11330_out0[0:0];
assign v$SEL5_12787_out0 = v$A_11331_out0[0:0];
assign v$SEL5_12789_out0 = v$A_11334_out0[0:0];
assign v$SEL5_12790_out0 = v$A_11335_out0[0:0];
assign v$SEL5_12798_out0 = v$A_11346_out0[0:0];
assign v$SEL5_12799_out0 = v$A_11347_out0[0:0];
assign v$G4_13187_out0 = v$G2_8130_out0 && v$WR0_1316_out0;
assign v$G6_13627_out0 = ((v$SEL11_15556_out0 && !v$SEL15_13612_out0) || (!v$SEL11_15556_out0) && v$SEL15_13612_out0);
assign v$G6_13628_out0 = ((v$SEL11_15557_out0 && !v$SEL15_13613_out0) || (!v$SEL11_15557_out0) && v$SEL15_13613_out0);
assign v$B1_14232_out0 = v$SEL9_10849_out0;
assign v$A1_14348_out0 = v$SEL4_7343_out0;
assign v$B_14437_out0 = v$B$EXP_16675_out0;
assign v$B_14441_out0 = v$B$EXP_16677_out0;
assign v$A$MANTISA_14549_out0 = v$A$MANTISA_17915_out0;
assign v$A4_15008_out0 = v$SEL1_18045_out0;
assign v$_16242_out0 = { v$C10_8949_out0,v$SEL12_16_out0 };
assign v$_16243_out0 = { v$C10_8950_out0,v$SEL12_17_out0 };
assign v$SEL2_16607_out0 = v$A_11326_out0[3:3];
assign v$SEL2_16608_out0 = v$A_11327_out0[3:3];
assign v$SEL2_16610_out0 = v$A_11330_out0[3:3];
assign v$SEL2_16611_out0 = v$A_11331_out0[3:3];
assign v$SEL2_16613_out0 = v$A_11334_out0[3:3];
assign v$SEL2_16614_out0 = v$A_11335_out0[3:3];
assign v$SEL2_16622_out0 = v$A_11346_out0[3:3];
assign v$SEL2_16623_out0 = v$A_11347_out0[3:3];
assign v$B2_16636_out0 = v$SEL8_12926_out0;
assign v$B$EXP_16674_out0 = v$SEL2_6970_out0;
assign v$B4_16928_out0 = v$SEL6_5807_out0;
assign v$B3_17862_out0 = v$SEL7_4178_out0;
assign v$G57_17955_out0 = v$G62_11967_out0 || v$G64_6432_out0;
assign v$B$32BIT_18471_out0 = v$_18260_out0;
assign v$B$32BIT_18472_out0 = v$_18261_out0;
assign v$SIGN_1366_out0 = v$SIGN_12760_out0;
assign v$SIGN_1367_out0 = v$SIGN_12760_out0;
assign v$G37_1519_out0 = !((v$B4_16928_out0 && !v$A4_15009_out0) || (!v$B4_16928_out0) && v$A4_15009_out0);
assign v$A0_1732_out0 = v$SEL5_12783_out0;
assign v$A0_1733_out0 = v$SEL5_12784_out0;
assign v$A0_1735_out0 = v$SEL5_12786_out0;
assign v$A0_1736_out0 = v$SEL5_12787_out0;
assign v$A0_1738_out0 = v$SEL5_12789_out0;
assign v$A0_1739_out0 = v$SEL5_12790_out0;
assign v$A0_1747_out0 = v$SEL5_12798_out0;
assign v$A0_1748_out0 = v$SEL5_12799_out0;
assign v$G5_2668_out0 = v$G4_13187_out0 || v$G3_2977_out0;
assign v$HALT_2899_out0 = v$HALT_7572_out0;
assign v$HALT_2900_out0 = v$HALT_7573_out0;
assign v$B$MANTISA_3002_out0 = v$MUX7_12742_out0;
assign v$G21_3534_out0 = ! v$B1_14232_out0;
assign v$G8_3738_out0 = !((v$A3_10714_out0 && !v$B3_17862_out0) || (!v$A3_10714_out0) && v$B3_17862_out0);
assign v$IN_4361_out0 = v$OUT_3176_out0;
assign v$IN_4365_out0 = v$OUT_3180_out0;
assign v$IS$SUB_4443_out0 = v$G6_13627_out0;
assign v$IS$SUB_4444_out0 = v$G6_13628_out0;
assign v$B_4826_out0 = v$B$32BIT_18471_out0;
assign v$B_4832_out0 = v$B$32BIT_18472_out0;
assign v$B$MANTISA_4909_out0 = v$B$MANTISA_4071_out0;
assign v$G36_5918_out0 = !((v$B3_17862_out0 && !v$A3_10714_out0) || (!v$B3_17862_out0) && v$A3_10714_out0);
assign v$G6_6561_out0 = ! v$B3_17862_out0;
assign v$SEL8_7275_out0 = v$B$32BIT_18471_out0[22:0];
assign v$SEL8_7276_out0 = v$B$32BIT_18472_out0[22:0];
assign v$G3_7488_out0 = !((v$A4_15009_out0 && !v$B4_16928_out0) || (!v$A4_15009_out0) && v$B4_16928_out0);
assign v$G90_8054_out0 = v$PHALT0$PREV_7612_out0 || v$G83_428_out0;
assign v$A2_8064_out0 = v$SEL3_8431_out0;
assign v$A2_8065_out0 = v$SEL3_8432_out0;
assign v$A2_8067_out0 = v$SEL3_8434_out0;
assign v$A2_8068_out0 = v$SEL3_8435_out0;
assign v$A2_8070_out0 = v$SEL3_8437_out0;
assign v$A2_8071_out0 = v$SEL3_8438_out0;
assign v$A2_8079_out0 = v$SEL3_8446_out0;
assign v$A2_8080_out0 = v$SEL3_8447_out0;
assign v$SEL1_8083_out0 = v$A_2543_out0[7:0];
assign v$SEL1_8084_out0 = v$A_2544_out0[7:0];
assign v$SEL1_8085_out0 = v$A_2545_out0[7:0];
assign v$SEL1_8086_out0 = v$A_2546_out0[7:0];
assign v$G17_8190_out0 = !((v$A0_1737_out0 && !v$B0_3657_out0) || (!v$A0_1737_out0) && v$B0_3657_out0);
assign v$SEL3_9050_out0 = v$B_14437_out0[7:4];
assign v$SEL3_9051_out0 = v$B_14441_out0[7:4];
assign v$A3_10709_out0 = v$SEL2_16607_out0;
assign v$A3_10710_out0 = v$SEL2_16608_out0;
assign v$A3_10712_out0 = v$SEL2_16610_out0;
assign v$A3_10713_out0 = v$SEL2_16611_out0;
assign v$A3_10715_out0 = v$SEL2_16613_out0;
assign v$A3_10716_out0 = v$SEL2_16614_out0;
assign v$A3_10724_out0 = v$SEL2_16622_out0;
assign v$A3_10725_out0 = v$SEL2_16623_out0;
assign v$SEL3_11894_out0 = v$A$MANTISA_14549_out0[22:0];
assign v$G23_12187_out0 = ! v$B0_3657_out0;
assign v$G33_13111_out0 = !((v$A0_1737_out0 && !v$B0_3657_out0) || (!v$A0_1737_out0) && v$B0_3657_out0);
assign v$G1_13190_out0 = ! v$B4_16928_out0;
assign v$G15_13655_out0 = !((v$A2_8069_out0 && !v$B2_16636_out0) || (!v$A2_8069_out0) && v$B2_16636_out0);
assign v$A1_14346_out0 = v$SEL4_7341_out0;
assign v$A1_14347_out0 = v$SEL4_7342_out0;
assign v$A1_14349_out0 = v$SEL4_7344_out0;
assign v$A1_14350_out0 = v$SEL4_7345_out0;
assign v$A1_14352_out0 = v$SEL4_7347_out0;
assign v$A1_14353_out0 = v$SEL4_7348_out0;
assign v$A1_14361_out0 = v$SEL4_7356_out0;
assign v$A1_14362_out0 = v$SEL4_7357_out0;
assign v$B_14436_out0 = v$B$EXP_16674_out0;
assign v$G35_14535_out0 = !((v$A2_8069_out0 && !v$B2_16636_out0) || (!v$A2_8069_out0) && v$B2_16636_out0);
assign v$RAM$ADDR_15228_out0 = v$RAMADDRMUX_418_out0;
assign v$RAM$ADDR_15229_out0 = v$RAMADDRMUX_419_out0;
assign v$_15349_out0 = { v$_16242_out0,v$C1_15921_out0 };
assign v$_15350_out0 = { v$_16243_out0,v$C1_15922_out0 };
assign v$SEL1_15748_out0 = v$A$MANTISA_14549_out0[22:0];
assign v$G12_16480_out0 = ! v$B2_16636_out0;
assign v$B$EXP_16672_out0 = v$SEL2_6968_out0;
assign v$B$EXP_16678_out0 = v$SEL2_6974_out0;
assign v$G16_16874_out0 = !((v$A1_14351_out0 && !v$B1_14232_out0) || (!v$A1_14351_out0) && v$B1_14232_out0);
assign v$G34_17304_out0 = !((v$A1_14351_out0 && !v$B1_14232_out0) || (!v$A1_14351_out0) && v$B1_14232_out0);
assign v$SEL2_17441_out0 = v$B_14437_out0[3:0];
assign v$SEL2_17442_out0 = v$B_14441_out0[3:0];
assign v$G89_17772_out0 = v$G85_6200_out0 || v$PHALT1$PREV_7363_out0;
assign v$SELIN_18215_out0 = v$G57_17955_out0;
assign v$SEL3_18618_out0 = v$A_2543_out0[11:8];
assign v$SEL3_18619_out0 = v$A_2544_out0[11:8];
assign v$SEL3_18620_out0 = v$A_2545_out0[11:8];
assign v$SEL3_18621_out0 = v$A_2546_out0[11:8];
assign v$A4XNORB4_1374_out0 = v$G3_7488_out0;
assign v$A0XNORB0_1444_out0 = v$G17_8190_out0;
assign v$SEL4_2280_out0 = v$B$MANTISA_4909_out0[22:0];
assign v$B$MANTISA_4070_out0 = v$B$MANTISA_3002_out0;
assign v$SEL7_4175_out0 = v$B_14436_out0[3:3];
assign v$A2XNORB2_4502_out0 = v$G15_13655_out0;
assign v$SEL6_5806_out0 = v$B_14436_out0[4:4];
assign v$RAM$ADDR_6413_out0 = v$RAM$ADDR_15228_out0;
assign v$RAM$ADDR_6414_out0 = v$RAM$ADDR_15229_out0;
assign v$G5_6946_out0 = v$A3_10714_out0 && v$G6_6561_out0;
assign v$SEL2_6969_out0 = v$B_4826_out0[30:23];
assign v$SEL2_6975_out0 = v$B_4832_out0[30:23];
assign v$RAMADDRESS_6988_out0 = v$RAM$ADDR_15228_out0;
assign v$RAMADDRESS_6989_out0 = v$RAM$ADDR_15229_out0;
assign v$G38_7303_out0 = v$G33_13111_out0 && v$G34_17304_out0;
assign v$V0_7423_out0 = v$G90_8054_out0;
assign v$_7615_out0 = { v$SEL8_7275_out0,v$C6_1568_out0 };
assign v$_7616_out0 = { v$SEL8_7276_out0,v$C6_1569_out0 };
assign v$IN_9567_out0 = v$IN_4361_out0;
assign v$IN_9571_out0 = v$IN_4365_out0;
assign v$G20_9894_out0 = v$A1_14351_out0 && v$G21_3534_out0;
assign v$G2_10402_out0 = v$A4_15009_out0 && v$G1_13190_out0;
assign v$SEL9_10846_out0 = v$B_14436_out0[1:1];
assign v$G25_10946_out0 = v$A0_1737_out0 && v$G23_12187_out0;
assign v$SEL2_11012_out0 = v$B$MANTISA_4909_out0[22:0];
assign v$A_11316_out0 = v$SEL3_18618_out0;
assign v$A_11317_out0 = v$SEL1_8083_out0;
assign v$A_11320_out0 = v$SEL3_18619_out0;
assign v$A_11321_out0 = v$SEL1_8084_out0;
assign v$A_11336_out0 = v$SEL3_18620_out0;
assign v$A_11337_out0 = v$SEL1_8085_out0;
assign v$A_11340_out0 = v$SEL3_18621_out0;
assign v$A_11341_out0 = v$SEL1_8086_out0;
assign v$SEL10_12615_out0 = v$B_14436_out0[0:0];
assign v$SEL8_12923_out0 = v$B_14436_out0[2:2];
assign v$B_14432_out0 = v$B$EXP_16672_out0;
assign v$B_14438_out0 = v$SEL3_9050_out0;
assign v$B_14439_out0 = v$SEL2_17441_out0;
assign v$B_14442_out0 = v$SEL3_9051_out0;
assign v$B_14443_out0 = v$SEL2_17442_out0;
assign v$B_14452_out0 = v$B$EXP_16678_out0;
assign v$A3XNORB3_14728_out0 = v$G8_3738_out0;
assign v$IS$SUB_15449_out0 = v$IS$SUB_4443_out0;
assign v$IS$SUB_15450_out0 = v$IS$SUB_4444_out0;
assign v$G11_15649_out0 = v$A2_8069_out0 && v$G12_16480_out0;
assign v$MUX2_15843_out0 = v$SELIN_18215_out0 ? v$MUX5_10896_out0 : v$MUX4_3842_out0;
assign v$ADDRESS_15901_out0 = v$RAM$ADDR_15228_out0;
assign v$ADDRESS_15902_out0 = v$RAM$ADDR_15229_out0;
assign v$A1XNORB1_16057_out0 = v$G16_16874_out0;
assign v$V1_16703_out0 = v$G89_17772_out0;
assign v$G39_17360_out0 = v$G36_5918_out0 && v$G37_1519_out0;
assign v$HALT_17681_out0 = v$HALT_2899_out0;
assign v$HALT_17682_out0 = v$HALT_2900_out0;
assign v$MEMHALT_17799_out0 = v$HALT_2899_out0;
assign v$MEMHALT_17800_out0 = v$HALT_2900_out0;
assign v$MUX5_1611_out0 = v$IS$32$BIT_10862_out0 ? v$_7615_out0 : v$_15349_out0;
assign v$MUX5_1612_out0 = v$IS$32$BIT_10863_out0 ? v$_7616_out0 : v$_15350_out0;
assign v$G7_2239_out0 = v$A4XNORB4_1374_out0 && v$G5_6946_out0;
assign v$B0_3654_out0 = v$SEL10_12615_out0;
assign v$SEL7_4172_out0 = v$B_14432_out0[3:3];
assign v$SEL7_4176_out0 = v$B_14438_out0[3:3];
assign v$SEL7_4177_out0 = v$B_14439_out0[3:3];
assign v$SEL7_4179_out0 = v$B_14442_out0[3:3];
assign v$SEL7_4180_out0 = v$B_14443_out0[3:3];
assign v$SEL7_4187_out0 = v$B_14452_out0[3:3];
assign v$G13_4411_out0 = v$A3XNORB3_14728_out0 && v$G11_15649_out0;
assign v$_4801_out0 = v$IN_9567_out0[13:0];
assign v$_4805_out0 = v$IN_9571_out0[13:0];
assign v$B$MANTISA_4908_out0 = v$B$MANTISA_4070_out0;
assign v$SEL6_5805_out0 = v$B_14432_out0[4:4];
assign v$SEL6_5808_out0 = v$B_14452_out0[4:4];
assign v$ADDRESS_5811_out0 = v$ADDRESS_15901_out0;
assign v$ADDRESS_5812_out0 = v$ADDRESS_15902_out0;
assign v$RAM$ADDR1_6454_out0 = v$RAM$ADDR_6414_out0;
assign v$SEL4_7334_out0 = v$A_11316_out0[1:1];
assign v$SEL4_7337_out0 = v$A_11320_out0[1:1];
assign v$SEL4_7349_out0 = v$A_11336_out0[1:1];
assign v$SEL4_7352_out0 = v$A_11340_out0[1:1];
assign v$A4$COMP$B4_7411_out0 = v$G2_10402_out0;
assign v$SEL3_8424_out0 = v$A_11316_out0[2:2];
assign v$SEL3_8427_out0 = v$A_11320_out0[2:2];
assign v$SEL3_8439_out0 = v$A_11336_out0[2:2];
assign v$SEL3_8442_out0 = v$A_11340_out0[2:2];
assign v$VALID1_8806_out0 = v$V1_16703_out0;
assign v$SEL1_10290_out0 = v$A_11317_out0[3:0];
assign v$SEL1_10291_out0 = v$A_11321_out0[3:0];
assign v$SEL1_10295_out0 = v$A_11337_out0[3:0];
assign v$SEL1_10296_out0 = v$A_11341_out0[3:0];
assign v$SEL9_10843_out0 = v$B_14432_out0[1:1];
assign v$SEL9_10847_out0 = v$B_14438_out0[1:1];
assign v$SEL9_10848_out0 = v$B_14439_out0[1:1];
assign v$SEL9_10850_out0 = v$B_14442_out0[1:1];
assign v$SEL9_10851_out0 = v$B_14443_out0[1:1];
assign v$SEL9_10858_out0 = v$B_14452_out0[1:1];
assign v$_11765_out0 = v$IN_9567_out0[15:15];
assign v$_11766_out0 = v$IN_9571_out0[15:15];
assign v$RAM$ADDR0_12525_out0 = v$RAM$ADDR_6413_out0;
assign v$SEL10_12612_out0 = v$B_14432_out0[0:0];
assign v$SEL10_12616_out0 = v$B_14438_out0[0:0];
assign v$SEL10_12617_out0 = v$B_14439_out0[0:0];
assign v$SEL10_12619_out0 = v$B_14442_out0[0:0];
assign v$SEL10_12620_out0 = v$B_14443_out0[0:0];
assign v$SEL10_12627_out0 = v$B_14452_out0[0:0];
assign v$RAMADDRESS_12721_out0 = v$RAMADDRESS_6988_out0;
assign v$RAMADDRESS_12722_out0 = v$RAMADDRESS_6989_out0;
assign v$SEL5_12776_out0 = v$A_11316_out0[0:0];
assign v$SEL5_12779_out0 = v$A_11320_out0[0:0];
assign v$SEL5_12791_out0 = v$A_11336_out0[0:0];
assign v$SEL5_12794_out0 = v$A_11340_out0[0:0];
assign v$HALT_12900_out0 = v$HALT_17681_out0;
assign v$HALT_12901_out0 = v$HALT_17682_out0;
assign v$SEL8_12920_out0 = v$B_14432_out0[2:2];
assign v$SEL8_12924_out0 = v$B_14438_out0[2:2];
assign v$SEL8_12925_out0 = v$B_14439_out0[2:2];
assign v$SEL8_12927_out0 = v$B_14442_out0[2:2];
assign v$SEL8_12928_out0 = v$B_14443_out0[2:2];
assign v$SEL8_12935_out0 = v$B_14452_out0[2:2];
assign v$G28_13027_out0 = v$A1XNORB1_16057_out0 && v$G25_10946_out0;
assign v$IS$SUB_13067_out0 = v$IS$SUB_15449_out0;
assign v$IS$SUB_13068_out0 = v$IS$SUB_15450_out0;
assign v$G22_13339_out0 = v$A2XNORB2_4502_out0 && v$G20_9894_out0;
assign v$G40_13372_out0 = v$G35_14535_out0 && v$G39_17360_out0;
assign v$VALID0_13405_out0 = v$V0_7423_out0;
assign v$_14164_out0 = v$IN_9567_out0[1:0];
assign v$_14165_out0 = v$IN_9571_out0[1:0];
assign v$B1_14229_out0 = v$SEL9_10846_out0;
assign v$_14600_out0 = v$IN_9567_out0[15:2];
assign v$_14604_out0 = v$IN_9571_out0[15:2];
assign v$_14634_out0 = v$IN_9567_out0[15:2];
assign v$_14638_out0 = v$IN_9571_out0[15:2];
assign v$SEL2_16600_out0 = v$A_11316_out0[3:3];
assign v$SEL2_16603_out0 = v$A_11320_out0[3:3];
assign v$SEL2_16615_out0 = v$A_11336_out0[3:3];
assign v$SEL2_16618_out0 = v$A_11340_out0[3:3];
assign v$B2_16633_out0 = v$SEL8_12923_out0;
assign v$B$EXP_16673_out0 = v$SEL2_6969_out0;
assign v$B$EXP_16679_out0 = v$SEL2_6975_out0;
assign v$_16748_out0 = v$IN_9567_out0[15:2];
assign v$_16752_out0 = v$IN_9571_out0[15:2];
assign v$B4_16927_out0 = v$SEL6_5806_out0;
assign v$_17057_out0 = v$IN_9567_out0[1:0];
assign v$_17058_out0 = v$IN_9571_out0[1:0];
assign v$SEL4_17330_out0 = v$A_11317_out0[7:4];
assign v$SEL4_17331_out0 = v$A_11321_out0[7:4];
assign v$SEL4_17335_out0 = v$A_11337_out0[7:4];
assign v$SEL4_17336_out0 = v$A_11341_out0[7:4];
assign v$B3_17859_out0 = v$SEL7_4175_out0;
assign v$G28_18550_out0 = v$MEMHALT_17799_out0 || v$PIPELINEHALT_14816_out0;
assign v$G28_18551_out0 = v$MEMHALT_17800_out0 || v$PIPELINEHALT_14817_out0;
assign v$_1478_out0 = { v$C1_7972_out0,v$_4801_out0 };
assign v$_1482_out0 = { v$C1_7976_out0,v$_4805_out0 };
assign v$G37_1518_out0 = !((v$B4_16927_out0 && !v$A4_15008_out0) || (!v$B4_16927_out0) && v$A4_15008_out0);
assign v$A0_1725_out0 = v$SEL5_12776_out0;
assign v$A0_1728_out0 = v$SEL5_12779_out0;
assign v$A0_1740_out0 = v$SEL5_12791_out0;
assign v$A0_1743_out0 = v$SEL5_12794_out0;
assign v$RAMAddress_2262_out0 = v$RAMADDRESS_12721_out0;
assign v$RAMAddress_2263_out0 = v$RAMADDRESS_12722_out0;
assign v$SEL4_2279_out0 = v$B$MANTISA_4908_out0[22:0];
assign v$EQ1_2953_out0 = v$ADDRESS_5811_out0 == 12'hff8;
assign v$EQ1_2954_out0 = v$ADDRESS_5812_out0 == 12'hff8;
assign v$G21_3531_out0 = ! v$B1_14229_out0;
assign v$EQ5_3551_out0 = v$ADDRESS_5811_out0 == 12'hff7;
assign v$EQ5_3552_out0 = v$ADDRESS_5812_out0 == 12'hff7;
assign v$B0_3651_out0 = v$SEL10_12612_out0;
assign v$B0_3655_out0 = v$SEL10_12616_out0;
assign v$B0_3656_out0 = v$SEL10_12617_out0;
assign v$B0_3658_out0 = v$SEL10_12619_out0;
assign v$B0_3659_out0 = v$SEL10_12620_out0;
assign v$B0_3666_out0 = v$SEL10_12627_out0;
assign v$G8_3735_out0 = !((v$A3_10711_out0 && !v$B3_17859_out0) || (!v$A3_10711_out0) && v$B3_17859_out0);
assign v$MUX3_3771_out0 = v$IS$SUB_13067_out0 ? v$C8_13621_out0 : v$C1_16233_out0;
assign v$MUX3_3772_out0 = v$IS$SUB_13068_out0 ? v$C8_13622_out0 : v$C1_16234_out0;
assign v$G27_4788_out0 = v$A2XNORB2_4502_out0 && v$G28_13027_out0;
assign v$A3$COMP$B3_4957_out0 = v$G7_2239_out0;
assign v$G18_4985_out0 = v$A3XNORB3_14728_out0 && v$G22_13339_out0;
assign v$G36_5915_out0 = !((v$B3_17859_out0 && !v$A3_10711_out0) || (!v$B3_17859_out0) && v$A3_10711_out0);
assign v$EXTHALT_6459_out0 = v$G28_18550_out0;
assign v$EXTHALT_6460_out0 = v$G28_18551_out0;
assign v$G6_6558_out0 = ! v$B3_17859_out0;
assign v$G3_7487_out0 = !((v$A4_15008_out0 && !v$B4_16927_out0) || (!v$A4_15008_out0) && v$B4_16927_out0);
assign v$MUX5_7954_out0 = v$S_10442_out0 ? v$_14164_out0 : v$C1_3018_out0;
assign v$MUX5_7955_out0 = v$S_10443_out0 ? v$_14165_out0 : v$C1_3019_out0;
assign v$A2_8057_out0 = v$SEL3_8424_out0;
assign v$A2_8060_out0 = v$SEL3_8427_out0;
assign v$A2_8072_out0 = v$SEL3_8439_out0;
assign v$A2_8075_out0 = v$SEL3_8442_out0;
assign v$G17_8187_out0 = !((v$A0_1734_out0 && !v$B0_3654_out0) || (!v$A0_1734_out0) && v$B0_3654_out0);
assign v$V0_9351_out0 = v$VALID0_13405_out0;
assign v$_9446_out0 = { v$_16748_out0,v$S$REG_3443_out0 };
assign v$_9450_out0 = { v$_16752_out0,v$S$REG_3444_out0 };
assign v$A3_10702_out0 = v$SEL2_16600_out0;
assign v$A3_10705_out0 = v$SEL2_16603_out0;
assign v$A3_10717_out0 = v$SEL2_16615_out0;
assign v$A3_10720_out0 = v$SEL2_16618_out0;
assign v$G41_10884_out0 = v$G38_7303_out0 && v$G40_13372_out0;
assign v$SEL2_11011_out0 = v$B$MANTISA_4908_out0[22:0];
assign v$A_11318_out0 = v$SEL4_17330_out0;
assign v$A_11319_out0 = v$SEL1_10290_out0;
assign v$A_11322_out0 = v$SEL4_17331_out0;
assign v$A_11323_out0 = v$SEL1_10291_out0;
assign v$A_11338_out0 = v$SEL4_17335_out0;
assign v$A_11339_out0 = v$SEL1_10295_out0;
assign v$A_11342_out0 = v$SEL4_17336_out0;
assign v$A_11343_out0 = v$SEL1_10296_out0;
assign v$EQ3_11712_out0 = v$ADDRESS_5811_out0 == 12'hffa;
assign v$EQ3_11713_out0 = v$ADDRESS_5812_out0 == 12'hffa;
assign v$G23_12184_out0 = ! v$B0_3654_out0;
assign v$G14_12645_out0 = v$A4XNORB4_1374_out0 && v$G13_4411_out0;
assign v$RAMADDR1_12657_out0 = v$RAM$ADDR1_6454_out0;
assign v$G33_13108_out0 = !((v$A0_1734_out0 && !v$B0_3654_out0) || (!v$A0_1734_out0) && v$B0_3654_out0);
assign v$G1_13189_out0 = ! v$B4_16927_out0;
assign v$_13221_out0 = { v$_11765_out0,v$_11765_out0 };
assign v$_13222_out0 = { v$_11766_out0,v$_11766_out0 };
assign v$_13305_out0 = { v$_14600_out0,v$_17057_out0 };
assign v$_13309_out0 = { v$_14604_out0,v$_17058_out0 };
assign v$G15_13652_out0 = !((v$A2_8066_out0 && !v$B2_16633_out0) || (!v$A2_8066_out0) && v$B2_16633_out0);
assign v$B1_14226_out0 = v$SEL9_10843_out0;
assign v$B1_14230_out0 = v$SEL9_10847_out0;
assign v$B1_14231_out0 = v$SEL9_10848_out0;
assign v$B1_14233_out0 = v$SEL9_10850_out0;
assign v$B1_14234_out0 = v$SEL9_10851_out0;
assign v$B1_14241_out0 = v$SEL9_10858_out0;
assign v$A1_14339_out0 = v$SEL4_7334_out0;
assign v$A1_14342_out0 = v$SEL4_7337_out0;
assign v$A1_14354_out0 = v$SEL4_7349_out0;
assign v$A1_14357_out0 = v$SEL4_7352_out0;
assign v$B_14433_out0 = v$B$EXP_16673_out0;
assign v$B_14453_out0 = v$B$EXP_16679_out0;
assign v$G35_14532_out0 = !((v$A2_8066_out0 && !v$B2_16633_out0) || (!v$A2_8066_out0) && v$B2_16633_out0);
assign v$CIN_15051_out0 = v$IS$SUB_13067_out0;
assign v$CIN_15054_out0 = v$IS$SUB_13068_out0;
assign v$EQ12_15107_out0 = v$ADDRESS_5811_out0 == 12'hff6;
assign v$EQ12_15108_out0 = v$ADDRESS_5812_out0 == 12'hff6;
assign v$S_15477_out0 = v$HALT_12900_out0;
assign v$S_15478_out0 = v$HALT_12901_out0;
assign v$B$MANTISA_15588_out0 = v$MUX5_1611_out0;
assign v$B$MANTISA_15589_out0 = v$MUX5_1612_out0;
assign v$G12_16477_out0 = ! v$B2_16633_out0;
assign v$EQ4_16578_out0 = v$ADDRESS_5811_out0 == 12'hffb;
assign v$EQ4_16579_out0 = v$ADDRESS_5812_out0 == 12'hffb;
assign v$B2_16630_out0 = v$SEL8_12920_out0;
assign v$B2_16634_out0 = v$SEL8_12924_out0;
assign v$B2_16635_out0 = v$SEL8_12925_out0;
assign v$B2_16637_out0 = v$SEL8_12927_out0;
assign v$B2_16638_out0 = v$SEL8_12928_out0;
assign v$B2_16645_out0 = v$SEL8_12935_out0;
assign v$G16_16871_out0 = !((v$A1_14348_out0 && !v$B1_14229_out0) || (!v$A1_14348_out0) && v$B1_14229_out0);
assign v$EQ2_16902_out0 = v$ADDRESS_5811_out0 == 12'hff9;
assign v$EQ2_16903_out0 = v$ADDRESS_5812_out0 == 12'hff9;
assign v$B4_16926_out0 = v$SEL6_5805_out0;
assign v$B4_16929_out0 = v$SEL6_5808_out0;
assign v$RAMADDR0_16982_out0 = v$RAM$ADDR0_12525_out0;
assign v$G34_17301_out0 = !((v$A1_14348_out0 && !v$B1_14229_out0) || (!v$A1_14348_out0) && v$B1_14229_out0);
assign v$V1_17836_out0 = v$VALID1_8806_out0;
assign v$B3_17856_out0 = v$SEL7_4172_out0;
assign v$B3_17860_out0 = v$SEL7_4176_out0;
assign v$B3_17861_out0 = v$SEL7_4177_out0;
assign v$B3_17863_out0 = v$SEL7_4179_out0;
assign v$B3_17864_out0 = v$SEL7_4180_out0;
assign v$B3_17871_out0 = v$SEL7_4187_out0;
assign v$G65_18211_out0 = v$HALT_12900_out0 || v$G64_6395_out0;
assign v$G65_18212_out0 = v$HALT_12901_out0 || v$G64_6396_out0;
assign v$G13_198_out0 = v$EQ12_15107_out0 && v$WEN_3683_out0;
assign v$G13_199_out0 = v$EQ12_15108_out0 && v$WEN_3684_out0;
assign v$MUX6_1311_out0 = v$FF1_16315_out0 ? v$S$REG_3443_out0 : v$_13221_out0;
assign v$MUX6_1312_out0 = v$FF1_16316_out0 ? v$S$REG_3444_out0 : v$_13222_out0;
assign v$A4XNORB4_1373_out0 = v$G3_7487_out0;
assign v$A0XNORB0_1441_out0 = v$G17_8187_out0;
assign v$G37_1517_out0 = !((v$B4_16926_out0 && !v$A4_15007_out0) || (!v$B4_16926_out0) && v$A4_15007_out0);
assign v$G37_1520_out0 = !((v$B4_16929_out0 && !v$A4_15010_out0) || (!v$B4_16929_out0) && v$A4_15010_out0);
assign v$A2$COMP$B2_1984_out0 = v$G14_12645_out0;
assign v$B$MANTISSA_2673_out0 = v$B$MANTISA_15588_out0;
assign v$B$MANTISSA_2674_out0 = v$B$MANTISA_15589_out0;
assign v$ADD_2955_out0 = v$RAMAddress_2262_out0;
assign v$ADD_2956_out0 = v$RAMAddress_2263_out0;
assign v$G21_3528_out0 = ! v$B1_14226_out0;
assign v$G21_3532_out0 = ! v$B1_14230_out0;
assign v$G21_3533_out0 = ! v$B1_14231_out0;
assign v$G21_3535_out0 = ! v$B1_14233_out0;
assign v$G21_3536_out0 = ! v$B1_14234_out0;
assign v$G21_3543_out0 = ! v$B1_14241_out0;
assign v$G8_3732_out0 = !((v$A3_10708_out0 && !v$B3_17856_out0) || (!v$A3_10708_out0) && v$B3_17856_out0);
assign v$G8_3736_out0 = !((v$A3_10712_out0 && !v$B3_17860_out0) || (!v$A3_10712_out0) && v$B3_17860_out0);
assign v$G8_3737_out0 = !((v$A3_10713_out0 && !v$B3_17861_out0) || (!v$A3_10713_out0) && v$B3_17861_out0);
assign v$G8_3739_out0 = !((v$A3_10715_out0 && !v$B3_17863_out0) || (!v$A3_10715_out0) && v$B3_17863_out0);
assign v$G8_3740_out0 = !((v$A3_10716_out0 && !v$B3_17864_out0) || (!v$A3_10716_out0) && v$B3_17864_out0);
assign v$G8_3747_out0 = !((v$A3_10723_out0 && !v$B3_17871_out0) || (!v$A3_10723_out0) && v$B3_17871_out0);
assign v$A2XNORB2_4499_out0 = v$G15_13652_out0;
assign v$G30_4923_out0 = !(v$EXTHALT_6459_out0 || v$STPHALT_4317_out0);
assign v$G30_4924_out0 = !(v$EXTHALT_6460_out0 || v$STPHALT_4318_out0);
assign v$G36_5912_out0 = !((v$B3_17856_out0 && !v$A3_10708_out0) || (!v$B3_17856_out0) && v$A3_10708_out0);
assign v$G36_5916_out0 = !((v$B3_17860_out0 && !v$A3_10712_out0) || (!v$B3_17860_out0) && v$A3_10712_out0);
assign v$G36_5917_out0 = !((v$B3_17861_out0 && !v$A3_10713_out0) || (!v$B3_17861_out0) && v$A3_10713_out0);
assign v$G36_5919_out0 = !((v$B3_17863_out0 && !v$A3_10715_out0) || (!v$B3_17863_out0) && v$A3_10715_out0);
assign v$G36_5920_out0 = !((v$B3_17864_out0 && !v$A3_10716_out0) || (!v$B3_17864_out0) && v$A3_10716_out0);
assign v$G36_5927_out0 = !((v$B3_17871_out0 && !v$A3_10723_out0) || (!v$B3_17871_out0) && v$A3_10723_out0);
assign v$G6_6555_out0 = ! v$B3_17856_out0;
assign v$G6_6559_out0 = ! v$B3_17860_out0;
assign v$G6_6560_out0 = ! v$B3_17861_out0;
assign v$G6_6562_out0 = ! v$B3_17863_out0;
assign v$G6_6563_out0 = ! v$B3_17864_out0;
assign v$G6_6570_out0 = ! v$B3_17871_out0;
assign v$MUX6_6903_out0 = v$G70_14028_out0 ? v$REG12_3330_out0 : v$RAMADDR1_12657_out0;
assign v$G5_6943_out0 = v$A3_10711_out0 && v$G6_6558_out0;
assign v$G38_7300_out0 = v$G33_13108_out0 && v$G34_17301_out0;
assign v$SEL4_7335_out0 = v$A_11318_out0[1:1];
assign v$SEL4_7336_out0 = v$A_11319_out0[1:1];
assign v$SEL4_7338_out0 = v$A_11322_out0[1:1];
assign v$SEL4_7339_out0 = v$A_11323_out0[1:1];
assign v$SEL4_7350_out0 = v$A_11338_out0[1:1];
assign v$SEL4_7351_out0 = v$A_11339_out0[1:1];
assign v$SEL4_7353_out0 = v$A_11342_out0[1:1];
assign v$SEL4_7354_out0 = v$A_11343_out0[1:1];
assign v$G3_7486_out0 = !((v$A4_15007_out0 && !v$B4_16926_out0) || (!v$A4_15007_out0) && v$B4_16926_out0);
assign v$G3_7489_out0 = !((v$A4_15010_out0 && !v$B4_16929_out0) || (!v$A4_15010_out0) && v$B4_16929_out0);
assign v$G3_7518_out0 = v$EQ2_16902_out0 && v$WEN_3683_out0;
assign v$G3_7519_out0 = v$EQ2_16903_out0 && v$WEN_3684_out0;
assign v$S_8019_out0 = v$S_15477_out0;
assign v$S_8020_out0 = v$S_15478_out0;
assign v$G17_8184_out0 = !((v$A0_1731_out0 && !v$B0_3651_out0) || (!v$A0_1731_out0) && v$B0_3651_out0);
assign v$G17_8188_out0 = !((v$A0_1735_out0 && !v$B0_3655_out0) || (!v$A0_1735_out0) && v$B0_3655_out0);
assign v$G17_8189_out0 = !((v$A0_1736_out0 && !v$B0_3656_out0) || (!v$A0_1736_out0) && v$B0_3656_out0);
assign v$G17_8191_out0 = !((v$A0_1738_out0 && !v$B0_3658_out0) || (!v$A0_1738_out0) && v$B0_3658_out0);
assign v$G17_8192_out0 = !((v$A0_1739_out0 && !v$B0_3659_out0) || (!v$A0_1739_out0) && v$B0_3659_out0);
assign v$G17_8199_out0 = !((v$A0_1746_out0 && !v$B0_3666_out0) || (!v$A0_1746_out0) && v$B0_3666_out0);
assign v$SEL3_8425_out0 = v$A_11318_out0[2:2];
assign v$SEL3_8426_out0 = v$A_11319_out0[2:2];
assign v$SEL3_8428_out0 = v$A_11322_out0[2:2];
assign v$SEL3_8429_out0 = v$A_11323_out0[2:2];
assign v$SEL3_8440_out0 = v$A_11338_out0[2:2];
assign v$SEL3_8441_out0 = v$A_11339_out0[2:2];
assign v$SEL3_8443_out0 = v$A_11342_out0[2:2];
assign v$SEL3_8444_out0 = v$A_11343_out0[2:2];
assign v$G66_8673_out0 = ! v$G65_18211_out0;
assign v$G66_8674_out0 = ! v$G65_18212_out0;
assign v$SEL3_9049_out0 = v$B_14433_out0[7:4];
assign v$SEL3_9054_out0 = v$B_14453_out0[7:4];
assign v$MUX3_9123_out0 = v$G66_8931_out0 ? v$REG9_16088_out0 : v$RAMADDR0_16982_out0;
assign v$G20_9891_out0 = v$A1_14348_out0 && v$G21_3531_out0;
assign v$G19_10248_out0 = v$A4XNORB4_1374_out0 && v$G18_4985_out0;
assign v$G2_10401_out0 = v$A4_15008_out0 && v$G1_13189_out0;
assign v$G25_10943_out0 = v$A0_1734_out0 && v$G23_12184_out0;
assign v$G23_12181_out0 = ! v$B0_3651_out0;
assign v$G23_12185_out0 = ! v$B0_3655_out0;
assign v$G23_12186_out0 = ! v$B0_3656_out0;
assign v$G23_12188_out0 = ! v$B0_3658_out0;
assign v$G23_12189_out0 = ! v$B0_3659_out0;
assign v$G23_12196_out0 = ! v$B0_3666_out0;
assign v$G5_12747_out0 = v$EQ5_3551_out0 && v$WEN_3683_out0;
assign v$G5_12748_out0 = v$EQ5_3552_out0 && v$WEN_3684_out0;
assign v$SEL5_12777_out0 = v$A_11318_out0[0:0];
assign v$SEL5_12778_out0 = v$A_11319_out0[0:0];
assign v$SEL5_12780_out0 = v$A_11322_out0[0:0];
assign v$SEL5_12781_out0 = v$A_11323_out0[0:0];
assign v$SEL5_12792_out0 = v$A_11338_out0[0:0];
assign v$SEL5_12793_out0 = v$A_11339_out0[0:0];
assign v$SEL5_12795_out0 = v$A_11342_out0[0:0];
assign v$SEL5_12796_out0 = v$A_11343_out0[0:0];
assign v$G33_13105_out0 = !((v$A0_1731_out0 && !v$B0_3651_out0) || (!v$A0_1731_out0) && v$B0_3651_out0);
assign v$G33_13109_out0 = !((v$A0_1735_out0 && !v$B0_3655_out0) || (!v$A0_1735_out0) && v$B0_3655_out0);
assign v$G33_13110_out0 = !((v$A0_1736_out0 && !v$B0_3656_out0) || (!v$A0_1736_out0) && v$B0_3656_out0);
assign v$G33_13112_out0 = !((v$A0_1738_out0 && !v$B0_3658_out0) || (!v$A0_1738_out0) && v$B0_3658_out0);
assign v$G33_13113_out0 = !((v$A0_1739_out0 && !v$B0_3659_out0) || (!v$A0_1739_out0) && v$B0_3659_out0);
assign v$G33_13120_out0 = !((v$A0_1746_out0 && !v$B0_3666_out0) || (!v$A0_1746_out0) && v$B0_3666_out0);
assign v$G1_13188_out0 = ! v$B4_16926_out0;
assign v$G1_13191_out0 = ! v$B4_16929_out0;
assign v$G15_13649_out0 = !((v$A2_8063_out0 && !v$B2_16630_out0) || (!v$A2_8063_out0) && v$B2_16630_out0);
assign v$G15_13653_out0 = !((v$A2_8067_out0 && !v$B2_16634_out0) || (!v$A2_8067_out0) && v$B2_16634_out0);
assign v$G15_13654_out0 = !((v$A2_8068_out0 && !v$B2_16635_out0) || (!v$A2_8068_out0) && v$B2_16635_out0);
assign v$G15_13656_out0 = !((v$A2_8070_out0 && !v$B2_16637_out0) || (!v$A2_8070_out0) && v$B2_16637_out0);
assign v$G15_13657_out0 = !((v$A2_8071_out0 && !v$B2_16638_out0) || (!v$A2_8071_out0) && v$B2_16638_out0);
assign v$G15_13664_out0 = !((v$A2_8078_out0 && !v$B2_16645_out0) || (!v$A2_8078_out0) && v$B2_16645_out0);
assign v$G2_13693_out0 = v$EQ3_11712_out0 && v$WEN_3683_out0;
assign v$G2_13694_out0 = v$EQ3_11713_out0 && v$WEN_3684_out0;
assign v$VALID_14495_out0 = v$V0_9351_out0;
assign v$VALID_14496_out0 = v$V1_17836_out0;
assign v$G35_14529_out0 = !((v$A2_8063_out0 && !v$B2_16630_out0) || (!v$A2_8063_out0) && v$B2_16630_out0);
assign v$G35_14533_out0 = !((v$A2_8067_out0 && !v$B2_16634_out0) || (!v$A2_8067_out0) && v$B2_16634_out0);
assign v$G35_14534_out0 = !((v$A2_8068_out0 && !v$B2_16635_out0) || (!v$A2_8068_out0) && v$B2_16635_out0);
assign v$G35_14536_out0 = !((v$A2_8070_out0 && !v$B2_16637_out0) || (!v$A2_8070_out0) && v$B2_16637_out0);
assign v$G35_14537_out0 = !((v$A2_8071_out0 && !v$B2_16638_out0) || (!v$A2_8071_out0) && v$B2_16638_out0);
assign v$G35_14544_out0 = !((v$A2_8078_out0 && !v$B2_16645_out0) || (!v$A2_8078_out0) && v$B2_16645_out0);
assign v$A3XNORB3_14725_out0 = v$G8_3735_out0;
assign v$G4_15127_out0 = v$EQ1_2953_out0 && v$WEN_3683_out0;
assign v$G4_15128_out0 = v$EQ1_2954_out0 && v$WEN_3684_out0;
assign v$G11_15646_out0 = v$A2_8066_out0 && v$G12_16477_out0;
assign v$G24_15696_out0 = v$A3XNORB3_14728_out0 && v$G27_4788_out0;
assign v$MUX4_15991_out0 = v$EN_16966_out0 ? v$_1478_out0 : v$IN_9567_out0;
assign v$MUX4_15995_out0 = v$EN_16970_out0 ? v$_1482_out0 : v$IN_9571_out0;
assign v$A1XNORB1_16054_out0 = v$G16_16871_out0;
assign v$G12_16474_out0 = ! v$B2_16630_out0;
assign v$G12_16478_out0 = ! v$B2_16634_out0;
assign v$G12_16479_out0 = ! v$B2_16635_out0;
assign v$G12_16481_out0 = ! v$B2_16637_out0;
assign v$G12_16482_out0 = ! v$B2_16638_out0;
assign v$G12_16489_out0 = ! v$B2_16645_out0;
assign v$G1_16496_out0 = v$EQ4_16578_out0 && v$WEN_3683_out0;
assign v$G1_16497_out0 = v$EQ4_16579_out0 && v$WEN_3684_out0;
assign v$SEL2_16601_out0 = v$A_11318_out0[3:3];
assign v$SEL2_16602_out0 = v$A_11319_out0[3:3];
assign v$SEL2_16604_out0 = v$A_11322_out0[3:3];
assign v$SEL2_16605_out0 = v$A_11323_out0[3:3];
assign v$SEL2_16616_out0 = v$A_11338_out0[3:3];
assign v$SEL2_16617_out0 = v$A_11339_out0[3:3];
assign v$SEL2_16619_out0 = v$A_11342_out0[3:3];
assign v$SEL2_16620_out0 = v$A_11343_out0[3:3];
assign v$G16_16868_out0 = !((v$A1_14345_out0 && !v$B1_14226_out0) || (!v$A1_14345_out0) && v$B1_14226_out0);
assign v$G16_16872_out0 = !((v$A1_14349_out0 && !v$B1_14230_out0) || (!v$A1_14349_out0) && v$B1_14230_out0);
assign v$G16_16873_out0 = !((v$A1_14350_out0 && !v$B1_14231_out0) || (!v$A1_14350_out0) && v$B1_14231_out0);
assign v$G16_16875_out0 = !((v$A1_14352_out0 && !v$B1_14233_out0) || (!v$A1_14352_out0) && v$B1_14233_out0);
assign v$G16_16876_out0 = !((v$A1_14353_out0 && !v$B1_14234_out0) || (!v$A1_14353_out0) && v$B1_14234_out0);
assign v$G16_16883_out0 = !((v$A1_14360_out0 && !v$B1_14241_out0) || (!v$A1_14360_out0) && v$B1_14241_out0);
assign v$G34_17298_out0 = !((v$A1_14345_out0 && !v$B1_14226_out0) || (!v$A1_14345_out0) && v$B1_14226_out0);
assign v$G34_17302_out0 = !((v$A1_14349_out0 && !v$B1_14230_out0) || (!v$A1_14349_out0) && v$B1_14230_out0);
assign v$G34_17303_out0 = !((v$A1_14350_out0 && !v$B1_14231_out0) || (!v$A1_14350_out0) && v$B1_14231_out0);
assign v$G34_17305_out0 = !((v$A1_14352_out0 && !v$B1_14233_out0) || (!v$A1_14352_out0) && v$B1_14233_out0);
assign v$G34_17306_out0 = !((v$A1_14353_out0 && !v$B1_14234_out0) || (!v$A1_14353_out0) && v$B1_14234_out0);
assign v$G34_17313_out0 = !((v$A1_14360_out0 && !v$B1_14241_out0) || (!v$A1_14360_out0) && v$B1_14241_out0);
assign v$CIN_17343_out0 = v$CIN_15051_out0;
assign v$CIN_17346_out0 = v$CIN_15054_out0;
assign v$G39_17359_out0 = v$G36_5915_out0 && v$G37_1518_out0;
assign v$SEL2_17440_out0 = v$B_14433_out0[3:0];
assign v$SEL2_17445_out0 = v$B_14453_out0[3:0];
assign v$SAME_18739_out0 = v$G41_10884_out0;
assign v$I3REGISTERWRITE_1264_out0 = v$G1_16496_out0;
assign v$I3REGISTERWRITE_1265_out0 = v$G1_16497_out0;
assign v$SEL4_1364_out0 = v$B$MANTISSA_2673_out0[23:12];
assign v$SEL4_1365_out0 = v$B$MANTISSA_2674_out0[23:12];
assign v$A4XNORB4_1372_out0 = v$G3_7486_out0;
assign v$A4XNORB4_1375_out0 = v$G3_7489_out0;
assign v$A0XNORB0_1438_out0 = v$G17_8184_out0;
assign v$A0XNORB0_1442_out0 = v$G17_8188_out0;
assign v$A0XNORB0_1443_out0 = v$G17_8189_out0;
assign v$A0XNORB0_1445_out0 = v$G17_8191_out0;
assign v$A0XNORB0_1446_out0 = v$G17_8192_out0;
assign v$A0XNORB0_1453_out0 = v$G17_8199_out0;
assign v$COUNTEREN_1625_out0 = v$G13_198_out0;
assign v$COUNTEREN_1626_out0 = v$G13_199_out0;
assign v$A0_1726_out0 = v$SEL5_12777_out0;
assign v$A0_1727_out0 = v$SEL5_12778_out0;
assign v$A0_1729_out0 = v$SEL5_12780_out0;
assign v$A0_1730_out0 = v$SEL5_12781_out0;
assign v$A0_1741_out0 = v$SEL5_12792_out0;
assign v$A0_1742_out0 = v$SEL5_12793_out0;
assign v$A0_1744_out0 = v$SEL5_12795_out0;
assign v$A0_1745_out0 = v$SEL5_12796_out0;
assign v$MUX1_1851_out0 = v$SELIN_18215_out0 ? v$MUX6_6903_out0 : v$MUX3_9123_out0;
assign v$G7_2238_out0 = v$A4XNORB4_1373_out0 && v$G5_6943_out0;
assign v$I1REGISTERWRITE_2931_out0 = v$G3_7518_out0;
assign v$I1REGISTERWRITE_2932_out0 = v$G3_7519_out0;
assign v$I0REGISTERWRITE_3355_out0 = v$G4_15127_out0;
assign v$I0REGISTERWRITE_3356_out0 = v$G4_15128_out0;
assign v$ModeRegAdd_4007_out0 = v$ADD_2955_out0 == 12'hffc;
assign v$ModeRegAdd_4008_out0 = v$ADD_2956_out0 == 12'hffc;
assign v$G13_4408_out0 = v$A3XNORB3_14725_out0 && v$G11_15646_out0;
assign v$A2XNORB2_4496_out0 = v$G15_13649_out0;
assign v$A2XNORB2_4500_out0 = v$G15_13653_out0;
assign v$A2XNORB2_4501_out0 = v$G15_13654_out0;
assign v$A2XNORB2_4503_out0 = v$G15_13656_out0;
assign v$A2XNORB2_4504_out0 = v$G15_13657_out0;
assign v$A2XNORB2_4511_out0 = v$G15_13664_out0;
assign v$MODEEN_5755_out0 = v$G5_12747_out0;
assign v$MODEEN_5756_out0 = v$G5_12748_out0;
assign v$G5_6940_out0 = v$A3_10708_out0 && v$G6_6555_out0;
assign v$G5_6944_out0 = v$A3_10712_out0 && v$G6_6559_out0;
assign v$G5_6945_out0 = v$A3_10713_out0 && v$G6_6560_out0;
assign v$G5_6947_out0 = v$A3_10715_out0 && v$G6_6562_out0;
assign v$G5_6948_out0 = v$A3_10716_out0 && v$G6_6563_out0;
assign v$G5_6955_out0 = v$A3_10723_out0 && v$G6_6570_out0;
assign v$G38_7297_out0 = v$G33_13105_out0 && v$G34_17298_out0;
assign v$G38_7301_out0 = v$G33_13109_out0 && v$G34_17302_out0;
assign v$G38_7302_out0 = v$G33_13110_out0 && v$G34_17303_out0;
assign v$G38_7304_out0 = v$G33_13112_out0 && v$G34_17305_out0;
assign v$G38_7305_out0 = v$G33_13113_out0 && v$G34_17306_out0;
assign v$G38_7312_out0 = v$G33_13120_out0 && v$G34_17313_out0;
assign v$A4$COMP$B4_7410_out0 = v$G2_10401_out0;
assign v$StatRegAdd_7741_out0 = v$ADD_2955_out0 == 12'hffd;
assign v$StatRegAdd_7742_out0 = v$ADD_2956_out0 == 12'hffd;
assign v$A2_8058_out0 = v$SEL3_8425_out0;
assign v$A2_8059_out0 = v$SEL3_8426_out0;
assign v$A2_8061_out0 = v$SEL3_8428_out0;
assign v$A2_8062_out0 = v$SEL3_8429_out0;
assign v$A2_8073_out0 = v$SEL3_8440_out0;
assign v$A2_8074_out0 = v$SEL3_8441_out0;
assign v$A2_8076_out0 = v$SEL3_8443_out0;
assign v$A2_8077_out0 = v$SEL3_8444_out0;
assign v$EN_9080_out0 = v$G30_4923_out0;
assign v$EN_9081_out0 = v$G30_4924_out0;
assign v$G20_9888_out0 = v$A1_14345_out0 && v$G21_3528_out0;
assign v$G20_9892_out0 = v$A1_14349_out0 && v$G21_3532_out0;
assign v$G20_9893_out0 = v$A1_14350_out0 && v$G21_3533_out0;
assign v$G20_9895_out0 = v$A1_14352_out0 && v$G21_3535_out0;
assign v$G20_9896_out0 = v$A1_14353_out0 && v$G21_3536_out0;
assign v$G20_9903_out0 = v$A1_14360_out0 && v$G21_3543_out0;
assign v$G2_10400_out0 = v$A4_15007_out0 && v$G1_13188_out0;
assign v$G2_10403_out0 = v$A4_15010_out0 && v$G1_13191_out0;
assign v$A3_10703_out0 = v$SEL2_16601_out0;
assign v$A3_10704_out0 = v$SEL2_16602_out0;
assign v$A3_10706_out0 = v$SEL2_16604_out0;
assign v$A3_10707_out0 = v$SEL2_16605_out0;
assign v$A3_10718_out0 = v$SEL2_16616_out0;
assign v$A3_10719_out0 = v$SEL2_16617_out0;
assign v$A3_10721_out0 = v$SEL2_16619_out0;
assign v$A3_10722_out0 = v$SEL2_16620_out0;
assign v$G25_10940_out0 = v$A0_1731_out0 && v$G23_12181_out0;
assign v$G25_10944_out0 = v$A0_1735_out0 && v$G23_12185_out0;
assign v$G25_10945_out0 = v$A0_1736_out0 && v$G23_12186_out0;
assign v$G25_10947_out0 = v$A0_1738_out0 && v$G23_12188_out0;
assign v$G25_10948_out0 = v$A0_1739_out0 && v$G23_12189_out0;
assign v$G25_10955_out0 = v$A0_1746_out0 && v$G23_12196_out0;
assign v$G26_11370_out0 = v$A4XNORB4_1374_out0 && v$G24_15696_out0;
assign v$_11809_out0 = { v$_14634_out0,v$MUX6_1311_out0 };
assign v$_11813_out0 = { v$_14638_out0,v$MUX6_1312_out0 };
assign v$I2REGISTERWRITE_11930_out0 = v$G2_13693_out0;
assign v$I2REGISTERWRITE_11931_out0 = v$G2_13694_out0;
assign v$MUX2_12039_out0 = v$G3_2606_out0 ? v$_9446_out0 : v$MUX4_15991_out0;
assign v$MUX2_12043_out0 = v$G3_2610_out0 ? v$_9450_out0 : v$MUX4_15995_out0;
assign v$A1$COMP$B1_12498_out0 = v$G19_10248_out0;
assign v$RXRegAdd_12974_out0 = v$ADD_2955_out0 == 12'hffe;
assign v$RXRegAdd_12975_out0 = v$ADD_2956_out0 == 12'hffe;
assign v$G28_13024_out0 = v$A1XNORB1_16054_out0 && v$G25_10943_out0;
assign v$G22_13336_out0 = v$A2XNORB2_4499_out0 && v$G20_9891_out0;
assign v$G40_13369_out0 = v$G35_14532_out0 && v$G39_17359_out0;
assign v$G40_13370_out0 = v$G35_14533_out0 && v$G36_5916_out0;
assign v$G40_13371_out0 = v$G35_14534_out0 && v$G36_5917_out0;
assign v$G40_13373_out0 = v$G35_14536_out0 && v$G36_5919_out0;
assign v$G40_13374_out0 = v$G35_14537_out0 && v$G36_5920_out0;
assign v$SEL2_13746_out0 = v$B$MANTISSA_2673_out0[11:0];
assign v$SEL2_13747_out0 = v$B$MANTISSA_2674_out0[11:0];
assign v$A1_14340_out0 = v$SEL4_7335_out0;
assign v$A1_14341_out0 = v$SEL4_7336_out0;
assign v$A1_14343_out0 = v$SEL4_7338_out0;
assign v$A1_14344_out0 = v$SEL4_7339_out0;
assign v$A1_14355_out0 = v$SEL4_7350_out0;
assign v$A1_14356_out0 = v$SEL4_7351_out0;
assign v$A1_14358_out0 = v$SEL4_7353_out0;
assign v$A1_14359_out0 = v$SEL4_7354_out0;
assign v$B_14434_out0 = v$SEL3_9049_out0;
assign v$B_14435_out0 = v$SEL2_17440_out0;
assign v$B_14454_out0 = v$SEL3_9054_out0;
assign v$B_14455_out0 = v$SEL2_17445_out0;
assign v$StatRegAdd1_14555_out0 = v$ADD_2955_out0 == 12'hffd;
assign v$StatRegAdd1_14556_out0 = v$ADD_2956_out0 == 12'hffd;
assign v$A3XNORB3_14722_out0 = v$G8_3732_out0;
assign v$A3XNORB3_14726_out0 = v$G8_3736_out0;
assign v$A3XNORB3_14727_out0 = v$G8_3737_out0;
assign v$A3XNORB3_14729_out0 = v$G8_3739_out0;
assign v$A3XNORB3_14730_out0 = v$G8_3740_out0;
assign v$A3XNORB3_14737_out0 = v$G8_3747_out0;
assign v$TXRegAdd_15600_out0 = v$ADD_2955_out0 == 12'hfff;
assign v$TXRegAdd_15601_out0 = v$ADD_2956_out0 == 12'hfff;
assign v$G11_15643_out0 = v$A2_8063_out0 && v$G12_16474_out0;
assign v$G11_15647_out0 = v$A2_8067_out0 && v$G12_16478_out0;
assign v$G11_15648_out0 = v$A2_8068_out0 && v$G12_16479_out0;
assign v$G11_15650_out0 = v$A2_8070_out0 && v$G12_16481_out0;
assign v$G11_15651_out0 = v$A2_8071_out0 && v$G12_16482_out0;
assign v$G11_15658_out0 = v$A2_8078_out0 && v$G12_16489_out0;
assign v$A1XNORB1_16051_out0 = v$G16_16868_out0;
assign v$A1XNORB1_16055_out0 = v$G16_16872_out0;
assign v$A1XNORB1_16056_out0 = v$G16_16873_out0;
assign v$A1XNORB1_16058_out0 = v$G16_16875_out0;
assign v$A1XNORB1_16059_out0 = v$G16_16876_out0;
assign v$A1XNORB1_16066_out0 = v$G16_16883_out0;
assign v$CIN_16107_out0 = v$CIN_17343_out0;
assign v$CIN_16110_out0 = v$CIN_17346_out0;
assign v$G39_17358_out0 = v$G36_5912_out0 && v$G37_1517_out0;
assign v$G39_17361_out0 = v$G36_5927_out0 && v$G37_1520_out0;
assign v$SAME_18367_out0 = v$SAME_18739_out0;
assign v$VALID_18670_out0 = v$VALID_14495_out0;
assign v$VALID_18671_out0 = v$VALID_14496_out0;
assign v$G7_2237_out0 = v$A4XNORB4_1372_out0 && v$G5_6940_out0;
assign v$G7_2240_out0 = v$A4XNORB4_1375_out0 && v$G5_6955_out0;
assign v$SEL7_4173_out0 = v$B_14434_out0[3:3];
assign v$SEL7_4174_out0 = v$B_14435_out0[3:3];
assign v$SEL7_4188_out0 = v$B_14454_out0[3:3];
assign v$SEL7_4189_out0 = v$B_14455_out0[3:3];
assign v$G13_4405_out0 = v$A3XNORB3_14722_out0 && v$G11_15643_out0;
assign v$G13_4409_out0 = v$A3XNORB3_14726_out0 && v$G11_15647_out0;
assign v$G13_4410_out0 = v$A3XNORB3_14727_out0 && v$G11_15648_out0;
assign v$G13_4412_out0 = v$A3XNORB3_14729_out0 && v$G11_15650_out0;
assign v$G13_4413_out0 = v$A3XNORB3_14730_out0 && v$G11_15651_out0;
assign v$G13_4420_out0 = v$A3XNORB3_14737_out0 && v$G11_15658_out0;
assign v$G27_4785_out0 = v$A2XNORB2_4499_out0 && v$G28_13024_out0;
assign v$A3$COMP$B3_4954_out0 = v$G7_2238_out0;
assign v$A3$COMP$B3_4955_out0 = v$G5_6944_out0;
assign v$A3$COMP$B3_4956_out0 = v$G5_6945_out0;
assign v$A3$COMP$B3_4958_out0 = v$G5_6947_out0;
assign v$A3$COMP$B3_4959_out0 = v$G5_6948_out0;
assign v$G18_4982_out0 = v$A3XNORB3_14725_out0 && v$G22_13336_out0;
assign v$MUX1_6678_out0 = v$G4_4030_out0 ? v$_11809_out0 : v$MUX2_12039_out0;
assign v$MUX1_6682_out0 = v$G4_4034_out0 ? v$_11813_out0 : v$MUX2_12043_out0;
assign v$A4$COMP$B4_7409_out0 = v$G2_10400_out0;
assign v$A4$COMP$B4_7412_out0 = v$G2_10403_out0;
assign v$G3_7598_out0 = v$TXRegAdd_15600_out0 && v$WEN_18392_out0;
assign v$G3_7599_out0 = v$TXRegAdd_15601_out0 && v$WEN_18393_out0;
assign v$G7_7726_out0 = v$StatRegAdd1_14555_out0 && v$G8_13403_out0;
assign v$G7_7727_out0 = v$StatRegAdd1_14556_out0 && v$G8_13404_out0;
assign v$A0$COMP$B0_7998_out0 = v$G26_11370_out0;
assign v$I0EN_8042_out0 = v$I0REGISTERWRITE_3355_out0;
assign v$I0EN_8043_out0 = v$I0REGISTERWRITE_3356_out0;
assign v$G5_8448_out0 = v$RXRegAdd_12974_out0 && v$G6_668_out0;
assign v$G5_8449_out0 = v$RXRegAdd_12975_out0 && v$G6_669_out0;
assign v$CINA_8509_out0 = v$CIN_16107_out0;
assign v$CINA_8632_out0 = v$CIN_16110_out0;
assign v$SEL9_10844_out0 = v$B_14434_out0[1:1];
assign v$SEL9_10845_out0 = v$B_14435_out0[1:1];
assign v$SEL9_10859_out0 = v$B_14454_out0[1:1];
assign v$SEL9_10860_out0 = v$B_14455_out0[1:1];
assign v$G41_10881_out0 = v$G38_7300_out0 && v$G40_13369_out0;
assign v$G41_10882_out0 = v$G38_7301_out0 && v$G40_13370_out0;
assign v$G41_10883_out0 = v$G38_7302_out0 && v$G40_13371_out0;
assign v$G41_10885_out0 = v$G38_7304_out0 && v$G40_13373_out0;
assign v$G41_10886_out0 = v$G38_7305_out0 && v$G40_13374_out0;
assign v$B_12130_out0 = v$SEL4_1364_out0;
assign v$B_12131_out0 = v$SEL2_13746_out0;
assign v$B_12132_out0 = v$SEL4_1365_out0;
assign v$B_12133_out0 = v$SEL2_13747_out0;
assign v$SEL10_12613_out0 = v$B_14434_out0[0:0];
assign v$SEL10_12614_out0 = v$B_14435_out0[0:0];
assign v$SEL10_12628_out0 = v$B_14454_out0[0:0];
assign v$SEL10_12629_out0 = v$B_14455_out0[0:0];
assign v$G14_12644_out0 = v$A4XNORB4_1373_out0 && v$G13_4408_out0;
assign v$SEL8_12921_out0 = v$B_14434_out0[2:2];
assign v$SEL8_12922_out0 = v$B_14435_out0[2:2];
assign v$SEL8_12936_out0 = v$B_14454_out0[2:2];
assign v$SEL8_12937_out0 = v$B_14455_out0[2:2];
assign v$G28_13021_out0 = v$A1XNORB1_16051_out0 && v$G25_10940_out0;
assign v$G28_13025_out0 = v$A1XNORB1_16055_out0 && v$G25_10944_out0;
assign v$G28_13026_out0 = v$A1XNORB1_16056_out0 && v$G25_10945_out0;
assign v$G28_13028_out0 = v$A1XNORB1_16058_out0 && v$G25_10947_out0;
assign v$G28_13029_out0 = v$A1XNORB1_16059_out0 && v$G25_10948_out0;
assign v$G28_13036_out0 = v$A1XNORB1_16066_out0 && v$G25_10955_out0;
assign v$G22_13333_out0 = v$A2XNORB2_4496_out0 && v$G20_9888_out0;
assign v$G22_13337_out0 = v$A2XNORB2_4500_out0 && v$G20_9892_out0;
assign v$G22_13338_out0 = v$A2XNORB2_4501_out0 && v$G20_9893_out0;
assign v$G22_13340_out0 = v$A2XNORB2_4503_out0 && v$G20_9895_out0;
assign v$G22_13341_out0 = v$A2XNORB2_4504_out0 && v$G20_9896_out0;
assign v$G22_13348_out0 = v$A2XNORB2_4511_out0 && v$G20_9903_out0;
assign v$G40_13366_out0 = v$G35_14529_out0 && v$G39_17358_out0;
assign v$G40_13381_out0 = v$G35_14544_out0 && v$G39_17361_out0;
assign v$COUNTEREN_13450_out0 = v$COUNTEREN_1625_out0;
assign v$COUNTEREN_13451_out0 = v$COUNTEREN_1626_out0;
assign v$RAMADDR_13607_out0 = v$MUX1_1851_out0;
assign v$ENMODE_14574_out0 = v$MODEEN_5755_out0;
assign v$ENMODE_14575_out0 = v$MODEEN_5756_out0;
assign v$G9_15590_out0 = v$ModeRegAdd_4007_out0 && v$WEN_18392_out0;
assign v$G9_15591_out0 = v$ModeRegAdd_4008_out0 && v$WEN_18393_out0;
assign v$I2EN_15746_out0 = v$I2REGISTERWRITE_11930_out0;
assign v$I2EN_15747_out0 = v$I2REGISTERWRITE_11931_out0;
assign v$G1_16401_out0 = v$StatRegAdd_7741_out0 && v$WEN_18392_out0;
assign v$G1_16402_out0 = v$StatRegAdd_7742_out0 && v$WEN_18393_out0;
assign v$I3EN_17775_out0 = v$I3REGISTERWRITE_1264_out0;
assign v$I3EN_17776_out0 = v$I3REGISTERWRITE_1265_out0;
assign v$VALID_17917_out0 = v$VALID_18670_out0;
assign v$VALID_17918_out0 = v$VALID_18671_out0;
assign v$I1EN_18402_out0 = v$I1REGISTERWRITE_2931_out0;
assign v$I1EN_18403_out0 = v$I1REGISTERWRITE_2932_out0;
assign v$G32_404_out0 = v$A1$COMP$B1_12498_out0 || v$A0$COMP$B0_7998_out0;
assign v$MUX3_1958_out0 = v$G8_1887_out0 ? v$_13305_out0 : v$MUX1_6678_out0;
assign v$MUX3_1962_out0 = v$G8_1891_out0 ? v$_13309_out0 : v$MUX1_6682_out0;
assign v$A2$COMP$B2_1981_out0 = v$G14_12644_out0;
assign v$A2$COMP$B2_1982_out0 = v$G13_4409_out0;
assign v$A2$COMP$B2_1983_out0 = v$G13_4410_out0;
assign v$A2$COMP$B2_1985_out0 = v$G13_4412_out0;
assign v$A2$COMP$B2_1986_out0 = v$G13_4413_out0;
assign v$B0_3652_out0 = v$SEL10_12613_out0;
assign v$B0_3653_out0 = v$SEL10_12614_out0;
assign v$B0_3667_out0 = v$SEL10_12628_out0;
assign v$B0_3668_out0 = v$SEL10_12629_out0;
assign v$VALID_3712_out0 = v$VALID_17917_out0;
assign v$VALID_3713_out0 = v$VALID_17918_out0;
assign v$ModeWrite_4452_out0 = v$G9_15590_out0;
assign v$ModeWrite_4453_out0 = v$G9_15591_out0;
assign v$G27_4782_out0 = v$A2XNORB2_4496_out0 && v$G28_13021_out0;
assign v$G27_4786_out0 = v$A2XNORB2_4500_out0 && v$G28_13025_out0;
assign v$G27_4787_out0 = v$A2XNORB2_4501_out0 && v$G28_13026_out0;
assign v$G27_4789_out0 = v$A2XNORB2_4503_out0 && v$G28_13028_out0;
assign v$G27_4790_out0 = v$A2XNORB2_4504_out0 && v$G28_13029_out0;
assign v$G27_4797_out0 = v$A2XNORB2_4511_out0 && v$G28_13036_out0;
assign v$A3$COMP$B3_4951_out0 = v$G7_2237_out0;
assign v$A3$COMP$B3_4966_out0 = v$G7_2240_out0;
assign v$G18_4979_out0 = v$A3XNORB3_14722_out0 && v$G22_13333_out0;
assign v$G18_4983_out0 = v$A3XNORB3_14726_out0 && v$G22_13337_out0;
assign v$G18_4984_out0 = v$A3XNORB3_14727_out0 && v$G22_13338_out0;
assign v$G18_4986_out0 = v$A3XNORB3_14729_out0 && v$G22_13340_out0;
assign v$G18_4987_out0 = v$A3XNORB3_14730_out0 && v$G22_13341_out0;
assign v$G18_4994_out0 = v$A3XNORB3_14737_out0 && v$G22_13348_out0;
assign v$THRESHOLD$WRITE_7236_out0 = v$COUNTEREN_13450_out0;
assign v$THRESHOLD$WRITE_7237_out0 = v$COUNTEREN_13451_out0;
assign v$ENMODE_7737_out0 = v$ENMODE_14574_out0;
assign v$ENMODE_7738_out0 = v$ENMODE_14575_out0;
assign v$RAMADDR_8766_out0 = v$RAMADDR_13607_out0;
assign v$SEL4_9574_out0 = v$B_12130_out0[11:8];
assign v$SEL4_9575_out0 = v$B_12131_out0[11:8];
assign v$SEL4_9576_out0 = v$B_12132_out0[11:8];
assign v$SEL4_9577_out0 = v$B_12133_out0[11:8];
assign v$STRead_9925_out0 = v$G7_7726_out0;
assign v$STRead_9926_out0 = v$G7_7727_out0;
assign v$STClr_10217_out0 = v$G1_16401_out0;
assign v$STClr_10218_out0 = v$G1_16402_out0;
assign v$G19_10247_out0 = v$A4XNORB4_1373_out0 && v$G18_4982_out0;
assign v$G41_10878_out0 = v$G38_7297_out0 && v$G40_13366_out0;
assign v$G41_10893_out0 = v$G38_7312_out0 && v$G40_13381_out0;
assign v$G14_12643_out0 = v$A4XNORB4_1372_out0 && v$G13_4405_out0;
assign v$G14_12646_out0 = v$A4XNORB4_1375_out0 && v$G13_4420_out0;
assign v$B1_14227_out0 = v$SEL9_10844_out0;
assign v$B1_14228_out0 = v$SEL9_10845_out0;
assign v$B1_14242_out0 = v$SEL9_10859_out0;
assign v$B1_14243_out0 = v$SEL9_10860_out0;
assign v$G24_15693_out0 = v$A3XNORB3_14725_out0 && v$G27_4785_out0;
assign v$RXRead_16365_out0 = v$G5_8448_out0;
assign v$RXRead_16366_out0 = v$G5_8449_out0;
assign v$B2_16631_out0 = v$SEL8_12921_out0;
assign v$B2_16632_out0 = v$SEL8_12922_out0;
assign v$B2_16646_out0 = v$SEL8_12936_out0;
assign v$B2_16647_out0 = v$SEL8_12937_out0;
assign v$TXWrite_17496_out0 = v$G3_7598_out0;
assign v$TXWrite_17497_out0 = v$G3_7599_out0;
assign v$SEL2_17517_out0 = v$B_12130_out0[7:0];
assign v$SEL2_17518_out0 = v$B_12131_out0[7:0];
assign v$SEL2_17519_out0 = v$B_12132_out0[7:0];
assign v$SEL2_17520_out0 = v$B_12133_out0[7:0];
assign v$B3_17857_out0 = v$SEL7_4173_out0;
assign v$B3_17858_out0 = v$SEL7_4174_out0;
assign v$B3_17872_out0 = v$SEL7_4188_out0;
assign v$B3_17873_out0 = v$SEL7_4189_out0;
assign v$SAME_18735_out0 = v$G41_10881_out0;
assign v$SAME_18737_out0 = v$G41_10882_out0;
assign v$SAME_18738_out0 = v$G41_10883_out0;
assign v$SAME_18741_out0 = v$G41_10885_out0;
assign v$SAME_18742_out0 = v$G41_10886_out0;
assign v$R_1489_out0 = v$VALID_3712_out0;
assign v$R_1490_out0 = v$VALID_3713_out0;
assign v$STATUSREAD_1637_out0 = v$STRead_9925_out0;
assign v$STATUSREAD_1638_out0 = v$STRead_9926_out0;
assign v$A2$COMP$B2_1978_out0 = v$G14_12643_out0;
assign v$A2$COMP$B2_1993_out0 = v$G14_12646_out0;
assign v$OUT_3177_out0 = v$MUX3_1958_out0;
assign v$OUT_3181_out0 = v$MUX3_1962_out0;
assign v$G21_3529_out0 = ! v$B1_14227_out0;
assign v$G21_3530_out0 = ! v$B1_14228_out0;
assign v$G21_3544_out0 = ! v$B1_14242_out0;
assign v$G21_3545_out0 = ! v$B1_14243_out0;
assign v$G8_3733_out0 = !((v$A3_10709_out0 && !v$B3_17857_out0) || (!v$A3_10709_out0) && v$B3_17857_out0);
assign v$G8_3734_out0 = !((v$A3_10710_out0 && !v$B3_17858_out0) || (!v$A3_10710_out0) && v$B3_17858_out0);
assign v$G8_3748_out0 = !((v$A3_10724_out0 && !v$B3_17872_out0) || (!v$A3_10724_out0) && v$B3_17872_out0);
assign v$G8_3749_out0 = !((v$A3_10725_out0 && !v$B3_17873_out0) || (!v$A3_10725_out0) && v$B3_17873_out0);
assign v$G36_5913_out0 = !((v$B3_17857_out0 && !v$A3_10709_out0) || (!v$B3_17857_out0) && v$A3_10709_out0);
assign v$G36_5914_out0 = !((v$B3_17858_out0 && !v$A3_10710_out0) || (!v$B3_17858_out0) && v$A3_10710_out0);
assign v$G36_5928_out0 = !((v$B3_17872_out0 && !v$A3_10724_out0) || (!v$B3_17872_out0) && v$A3_10724_out0);
assign v$G36_5929_out0 = !((v$B3_17873_out0 && !v$A3_10725_out0) || (!v$B3_17873_out0) && v$A3_10725_out0);
assign v$STATUSCLR_5953_out0 = v$STClr_10217_out0;
assign v$STATUSCLR_5954_out0 = v$STClr_10218_out0;
assign v$G6_6556_out0 = ! v$B3_17857_out0;
assign v$G6_6557_out0 = ! v$B3_17858_out0;
assign v$G6_6571_out0 = ! v$B3_17872_out0;
assign v$G6_6572_out0 = ! v$B3_17873_out0;
assign v$G17_8185_out0 = !((v$A0_1732_out0 && !v$B0_3652_out0) || (!v$A0_1732_out0) && v$B0_3652_out0);
assign v$G17_8186_out0 = !((v$A0_1733_out0 && !v$B0_3653_out0) || (!v$A0_1733_out0) && v$B0_3653_out0);
assign v$G17_8200_out0 = !((v$A0_1747_out0 && !v$B0_3667_out0) || (!v$A0_1747_out0) && v$B0_3667_out0);
assign v$G17_8201_out0 = !((v$A0_1748_out0 && !v$B0_3668_out0) || (!v$A0_1748_out0) && v$B0_3668_out0);
assign v$LOWER$SAME_10184_out0 = v$SAME_18738_out0;
assign v$LOWER$SAME_10185_out0 = v$SAME_18742_out0;
assign v$G19_10246_out0 = v$A4XNORB4_1372_out0 && v$G18_4979_out0;
assign v$G19_10249_out0 = v$A4XNORB4_1375_out0 && v$G18_4994_out0;
assign v$TXWRITE_11109_out0 = v$TXWrite_17496_out0;
assign v$TXWRITE_11110_out0 = v$TXWrite_17497_out0;
assign v$G26_11369_out0 = v$A4XNORB4_1373_out0 && v$G24_15693_out0;
assign v$G23_12182_out0 = ! v$B0_3652_out0;
assign v$G23_12183_out0 = ! v$B0_3653_out0;
assign v$G23_12197_out0 = ! v$B0_3667_out0;
assign v$G23_12198_out0 = ! v$B0_3668_out0;
assign v$A1$COMP$B1_12495_out0 = v$G19_10247_out0;
assign v$A1$COMP$B1_12496_out0 = v$G18_4983_out0;
assign v$A1$COMP$B1_12497_out0 = v$G18_4984_out0;
assign v$A1$COMP$B1_12499_out0 = v$G18_4986_out0;
assign v$A1$COMP$B1_12500_out0 = v$G18_4987_out0;
assign v$G33_13106_out0 = !((v$A0_1732_out0 && !v$B0_3652_out0) || (!v$A0_1732_out0) && v$B0_3652_out0);
assign v$G33_13107_out0 = !((v$A0_1733_out0 && !v$B0_3653_out0) || (!v$A0_1733_out0) && v$B0_3653_out0);
assign v$G33_13121_out0 = !((v$A0_1747_out0 && !v$B0_3667_out0) || (!v$A0_1747_out0) && v$B0_3667_out0);
assign v$G33_13122_out0 = !((v$A0_1748_out0 && !v$B0_3668_out0) || (!v$A0_1748_out0) && v$B0_3668_out0);
assign v$G5_13549_out0 = v$EQUAL_15828_out0 || v$THRESHOLD$WRITE_7236_out0;
assign v$G5_13550_out0 = v$EQUAL_15829_out0 || v$THRESHOLD$WRITE_7237_out0;
assign v$G15_13650_out0 = !((v$A2_8064_out0 && !v$B2_16631_out0) || (!v$A2_8064_out0) && v$B2_16631_out0);
assign v$G15_13651_out0 = !((v$A2_8065_out0 && !v$B2_16632_out0) || (!v$A2_8065_out0) && v$B2_16632_out0);
assign v$G15_13665_out0 = !((v$A2_8079_out0 && !v$B2_16646_out0) || (!v$A2_8079_out0) && v$B2_16646_out0);
assign v$G15_13666_out0 = !((v$A2_8080_out0 && !v$B2_16647_out0) || (!v$A2_8080_out0) && v$B2_16647_out0);
assign v$B_14424_out0 = v$SEL4_9574_out0;
assign v$B_14425_out0 = v$SEL2_17517_out0;
assign v$B_14428_out0 = v$SEL4_9575_out0;
assign v$B_14429_out0 = v$SEL2_17518_out0;
assign v$B_14444_out0 = v$SEL4_9576_out0;
assign v$B_14445_out0 = v$SEL2_17519_out0;
assign v$B_14448_out0 = v$SEL4_9577_out0;
assign v$B_14449_out0 = v$SEL2_17520_out0;
assign v$G35_14530_out0 = !((v$A2_8064_out0 && !v$B2_16631_out0) || (!v$A2_8064_out0) && v$B2_16631_out0);
assign v$G35_14531_out0 = !((v$A2_8065_out0 && !v$B2_16632_out0) || (!v$A2_8065_out0) && v$B2_16632_out0);
assign v$G35_14545_out0 = !((v$A2_8079_out0 && !v$B2_16646_out0) || (!v$A2_8079_out0) && v$B2_16646_out0);
assign v$G35_14546_out0 = !((v$A2_8080_out0 && !v$B2_16647_out0) || (!v$A2_8080_out0) && v$B2_16647_out0);
assign v$MODEWRITE_14714_out0 = v$ModeWrite_4452_out0;
assign v$MODEWRITE_14715_out0 = v$ModeWrite_4453_out0;
assign v$HIGHER$SAME_15023_out0 = v$SAME_18737_out0;
assign v$HIGHER$SAME_15024_out0 = v$SAME_18741_out0;
assign v$G31_15518_out0 = v$A2$COMP$B2_1984_out0 || v$G32_404_out0;
assign v$G24_15690_out0 = v$A3XNORB3_14722_out0 && v$G27_4782_out0;
assign v$G24_15694_out0 = v$A3XNORB3_14726_out0 && v$G27_4786_out0;
assign v$G24_15695_out0 = v$A3XNORB3_14727_out0 && v$G27_4787_out0;
assign v$G24_15697_out0 = v$A3XNORB3_14729_out0 && v$G27_4789_out0;
assign v$G24_15698_out0 = v$A3XNORB3_14730_out0 && v$G27_4790_out0;
assign v$G24_15705_out0 = v$A3XNORB3_14737_out0 && v$G27_4797_out0;
assign v$RXREAD_15854_out0 = v$RXRead_16365_out0;
assign v$RXREAD_15855_out0 = v$RXRead_16366_out0;
assign v$EN_15897_out0 = v$ENMODE_7737_out0;
assign v$EN_15898_out0 = v$ENMODE_7738_out0;
assign v$G12_16475_out0 = ! v$B2_16631_out0;
assign v$G12_16476_out0 = ! v$B2_16632_out0;
assign v$G12_16490_out0 = ! v$B2_16646_out0;
assign v$G12_16491_out0 = ! v$B2_16647_out0;
assign v$G16_16869_out0 = !((v$A1_14346_out0 && !v$B1_14227_out0) || (!v$A1_14346_out0) && v$B1_14227_out0);
assign v$G16_16870_out0 = !((v$A1_14347_out0 && !v$B1_14228_out0) || (!v$A1_14347_out0) && v$B1_14228_out0);
assign v$G16_16884_out0 = !((v$A1_14361_out0 && !v$B1_14242_out0) || (!v$A1_14361_out0) && v$B1_14242_out0);
assign v$G16_16885_out0 = !((v$A1_14362_out0 && !v$B1_14243_out0) || (!v$A1_14362_out0) && v$B1_14243_out0);
assign v$G34_17299_out0 = !((v$A1_14346_out0 && !v$B1_14227_out0) || (!v$A1_14346_out0) && v$B1_14227_out0);
assign v$G34_17300_out0 = !((v$A1_14347_out0 && !v$B1_14228_out0) || (!v$A1_14347_out0) && v$B1_14228_out0);
assign v$G34_17314_out0 = !((v$A1_14361_out0 && !v$B1_14242_out0) || (!v$A1_14361_out0) && v$B1_14242_out0);
assign v$G34_17315_out0 = !((v$A1_14362_out0 && !v$B1_14243_out0) || (!v$A1_14362_out0) && v$B1_14243_out0);
assign v$SAME_18365_out0 = v$SAME_18735_out0;
assign v$RAMADDR_18656_out0 = v$RAMADDR_8766_out0;
assign v$SAME_18731_out0 = v$G41_10878_out0;
assign v$SAME_18751_out0 = v$G41_10893_out0;
assign v$A0XNORB0_1439_out0 = v$G17_8185_out0;
assign v$A0XNORB0_1440_out0 = v$G17_8186_out0;
assign v$A0XNORB0_1454_out0 = v$G17_8200_out0;
assign v$A0XNORB0_1455_out0 = v$G17_8201_out0;
assign v$R_1588_out0 = v$R_1489_out0;
assign v$R_1589_out0 = v$R_1490_out0;
assign v$G30_1781_out0 = v$A3$COMP$B3_4957_out0 || v$G31_15518_out0;
assign v$WREN_2534_out0 = v$TXWRITE_11109_out0;
assign v$WREN_2535_out0 = v$TXWRITE_11110_out0;
assign v$SEL7_4166_out0 = v$B_14424_out0[3:3];
assign v$SEL7_4169_out0 = v$B_14428_out0[3:3];
assign v$SEL7_4181_out0 = v$B_14444_out0[3:3];
assign v$SEL7_4184_out0 = v$B_14448_out0[3:3];
assign v$G1_4213_out0 = v$STATUSREAD_1637_out0 || v$RXREAD_15854_out0;
assign v$G1_4214_out0 = v$STATUSREAD_1638_out0 || v$RXREAD_15855_out0;
assign v$IN_4362_out0 = v$OUT_3177_out0;
assign v$IN_4366_out0 = v$OUT_3181_out0;
assign v$A2XNORB2_4497_out0 = v$G15_13650_out0;
assign v$A2XNORB2_4498_out0 = v$G15_13651_out0;
assign v$A2XNORB2_4512_out0 = v$G15_13665_out0;
assign v$A2XNORB2_4513_out0 = v$G15_13666_out0;
assign v$RXreset_5959_out0 = v$RXREAD_15854_out0;
assign v$RXreset_5960_out0 = v$RXREAD_15855_out0;
assign v$G5_6941_out0 = v$A3_10709_out0 && v$G6_6556_out0;
assign v$G5_6942_out0 = v$A3_10710_out0 && v$G6_6557_out0;
assign v$G5_6956_out0 = v$A3_10724_out0 && v$G6_6571_out0;
assign v$G5_6957_out0 = v$A3_10725_out0 && v$G6_6572_out0;
assign v$_7277_out0 = v$RAMADDR_18656_out0[3:0];
assign v$_7277_out1 = v$RAMADDR_18656_out0[11:8];
assign v$G38_7298_out0 = v$G33_13106_out0 && v$G34_17299_out0;
assign v$G38_7299_out0 = v$G33_13107_out0 && v$G34_17300_out0;
assign v$G38_7313_out0 = v$G33_13121_out0 && v$G34_17314_out0;
assign v$G38_7314_out0 = v$G33_13122_out0 && v$G34_17315_out0;
assign v$A0$COMP$B0_7995_out0 = v$G26_11369_out0;
assign v$A0$COMP$B0_7996_out0 = v$G24_15694_out0;
assign v$A0$COMP$B0_7997_out0 = v$G24_15695_out0;
assign v$A0$COMP$B0_7999_out0 = v$G24_15697_out0;
assign v$A0$COMP$B0_8000_out0 = v$G24_15698_out0;
assign v$SEL3_9047_out0 = v$B_14425_out0[7:4];
assign v$SEL3_9048_out0 = v$B_14429_out0[7:4];
assign v$SEL3_9052_out0 = v$B_14445_out0[7:4];
assign v$SEL3_9053_out0 = v$B_14449_out0[7:4];
assign v$G1_9389_out0 = v$LOWER$SAME_10184_out0 && v$HIGHER$SAME_15023_out0;
assign v$G1_9390_out0 = v$LOWER$SAME_10185_out0 && v$HIGHER$SAME_15024_out0;
assign v$G20_9889_out0 = v$A1_14346_out0 && v$G21_3529_out0;
assign v$G20_9890_out0 = v$A1_14347_out0 && v$G21_3530_out0;
assign v$G20_9904_out0 = v$A1_14361_out0 && v$G21_3544_out0;
assign v$G20_9905_out0 = v$A1_14362_out0 && v$G21_3545_out0;
assign v$SEL9_10837_out0 = v$B_14424_out0[1:1];
assign v$SEL9_10840_out0 = v$B_14428_out0[1:1];
assign v$SEL9_10852_out0 = v$B_14444_out0[1:1];
assign v$SEL9_10855_out0 = v$B_14448_out0[1:1];
assign v$G25_10941_out0 = v$A0_1732_out0 && v$G23_12182_out0;
assign v$G25_10942_out0 = v$A0_1733_out0 && v$G23_12183_out0;
assign v$G25_10956_out0 = v$A0_1747_out0 && v$G23_12197_out0;
assign v$G25_10957_out0 = v$A0_1748_out0 && v$G23_12198_out0;
assign v$G26_11368_out0 = v$A4XNORB4_1372_out0 && v$G24_15690_out0;
assign v$G26_11371_out0 = v$A4XNORB4_1375_out0 && v$G24_15705_out0;
assign v$A1$COMP$B1_12492_out0 = v$G19_10246_out0;
assign v$A1$COMP$B1_12507_out0 = v$G19_10249_out0;
assign v$SEL10_12606_out0 = v$B_14424_out0[0:0];
assign v$SEL10_12609_out0 = v$B_14428_out0[0:0];
assign v$SEL10_12621_out0 = v$B_14444_out0[0:0];
assign v$SEL10_12624_out0 = v$B_14448_out0[0:0];
assign v$Clear_12750_out0 = v$STATUSCLR_5953_out0;
assign v$Clear_12751_out0 = v$STATUSCLR_5954_out0;
assign v$SEL8_12914_out0 = v$B_14424_out0[2:2];
assign v$SEL8_12917_out0 = v$B_14428_out0[2:2];
assign v$SEL8_12929_out0 = v$B_14444_out0[2:2];
assign v$SEL8_12932_out0 = v$B_14448_out0[2:2];
assign v$G40_13367_out0 = v$G35_14530_out0 && v$G36_5913_out0;
assign v$G40_13368_out0 = v$G35_14531_out0 && v$G36_5914_out0;
assign v$G40_13382_out0 = v$G35_14545_out0 && v$G36_5928_out0;
assign v$G40_13383_out0 = v$G35_14546_out0 && v$G36_5929_out0;
assign v$TXSet_14337_out0 = v$TXWRITE_11109_out0;
assign v$TXSet_14338_out0 = v$TXWRITE_11110_out0;
assign v$A3XNORB3_14723_out0 = v$G8_3733_out0;
assign v$A3XNORB3_14724_out0 = v$G8_3734_out0;
assign v$A3XNORB3_14738_out0 = v$G8_3748_out0;
assign v$A3XNORB3_14739_out0 = v$G8_3749_out0;
assign v$G11_15644_out0 = v$A2_8064_out0 && v$G12_16475_out0;
assign v$G11_15645_out0 = v$A2_8065_out0 && v$G12_16476_out0;
assign v$G11_15659_out0 = v$A2_8079_out0 && v$G12_16490_out0;
assign v$G11_15660_out0 = v$A2_8080_out0 && v$G12_16491_out0;
assign v$A1XNORB1_16052_out0 = v$G16_16869_out0;
assign v$A1XNORB1_16053_out0 = v$G16_16870_out0;
assign v$A1XNORB1_16067_out0 = v$G16_16884_out0;
assign v$A1XNORB1_16068_out0 = v$G16_16885_out0;
assign v$SEL2_17438_out0 = v$B_14425_out0[3:0];
assign v$SEL2_17439_out0 = v$B_14429_out0[3:0];
assign v$SEL2_17443_out0 = v$B_14445_out0[3:0];
assign v$SEL2_17444_out0 = v$B_14449_out0[3:0];
assign v$MUX1_18328_out0 = v$G5_13549_out0 ? v$C3_12205_out0 : v$A1_13701_out0;
assign v$MUX1_18329_out0 = v$G5_13550_out0 ? v$C3_12206_out0 : v$A1_13702_out0;
assign v$SAME_18363_out0 = v$SAME_18731_out0;
assign v$SAME_18369_out0 = v$SAME_18751_out0;
assign v$G32_401_out0 = v$A1$COMP$B1_12495_out0 || v$A0$COMP$B0_7995_out0;
assign v$G32_402_out0 = v$A1$COMP$B1_12496_out0 || v$A0$COMP$B0_7996_out0;
assign v$G32_403_out0 = v$A1$COMP$B1_12497_out0 || v$A0$COMP$B0_7997_out0;
assign v$G32_405_out0 = v$A1$COMP$B1_12499_out0 || v$A0$COMP$B0_7999_out0;
assign v$G32_406_out0 = v$A1$COMP$B1_12500_out0 || v$A0$COMP$B0_8000_out0;
assign v$SEL8_1968_out0 = v$_7277_out1[7:7];
assign v$SEL3_3126_out0 = v$_7277_out1[2:2];
assign v$B0_3645_out0 = v$SEL10_12606_out0;
assign v$B0_3648_out0 = v$SEL10_12609_out0;
assign v$B0_3660_out0 = v$SEL10_12621_out0;
assign v$B0_3663_out0 = v$SEL10_12624_out0;
assign v$G13_4406_out0 = v$A3XNORB3_14723_out0 && v$G11_15644_out0;
assign v$G13_4407_out0 = v$A3XNORB3_14724_out0 && v$G11_15645_out0;
assign v$G13_4421_out0 = v$A3XNORB3_14738_out0 && v$G11_15659_out0;
assign v$G13_4422_out0 = v$A3XNORB3_14739_out0 && v$G11_15660_out0;
assign v$A3$COMP$B3_4952_out0 = v$G5_6941_out0;
assign v$A3$COMP$B3_4953_out0 = v$G5_6942_out0;
assign v$A3$COMP$B3_4967_out0 = v$G5_6956_out0;
assign v$A3$COMP$B3_4968_out0 = v$G5_6957_out0;
assign v$SEL1_7005_out0 = v$_7277_out1[0:0];
assign v$A0$COMP$B0_7992_out0 = v$G26_11368_out0;
assign v$A0$COMP$B0_8007_out0 = v$G26_11371_out0;
assign v$IN_9568_out0 = v$IN_4362_out0;
assign v$IN_9572_out0 = v$IN_4366_out0;
assign v$G29_10300_out0 = v$A4$COMP$B4_7411_out0 || v$G30_1781_out0;
assign v$G41_10879_out0 = v$G38_7298_out0 && v$G40_13367_out0;
assign v$G41_10880_out0 = v$G38_7299_out0 && v$G40_13368_out0;
assign v$G41_10894_out0 = v$G38_7313_out0 && v$G40_13382_out0;
assign v$G41_10895_out0 = v$G38_7314_out0 && v$G40_13383_out0;
assign v$WREN_10997_out0 = v$WREN_2534_out0;
assign v$WREN_10998_out0 = v$WREN_2535_out0;
assign v$SEL5_11625_out0 = v$_7277_out1[4:4];
assign v$TXSet_12652_out0 = v$TXSet_14337_out0;
assign v$TXSet_12653_out0 = v$TXSet_14338_out0;
assign v$G28_13022_out0 = v$A1XNORB1_16052_out0 && v$G25_10941_out0;
assign v$G28_13023_out0 = v$A1XNORB1_16053_out0 && v$G25_10942_out0;
assign v$G28_13037_out0 = v$A1XNORB1_16067_out0 && v$G25_10956_out0;
assign v$G28_13038_out0 = v$A1XNORB1_16068_out0 && v$G25_10957_out0;
assign v$G22_13334_out0 = v$A2XNORB2_4497_out0 && v$G20_9889_out0;
assign v$G22_13335_out0 = v$A2XNORB2_4498_out0 && v$G20_9890_out0;
assign v$G22_13349_out0 = v$A2XNORB2_4512_out0 && v$G20_9904_out0;
assign v$G22_13350_out0 = v$A2XNORB2_4513_out0 && v$G20_9905_out0;
assign v$B1_14220_out0 = v$SEL9_10837_out0;
assign v$B1_14223_out0 = v$SEL9_10840_out0;
assign v$B1_14235_out0 = v$SEL9_10852_out0;
assign v$B1_14238_out0 = v$SEL9_10855_out0;
assign v$SEL6_14244_out0 = v$_7277_out1[5:5];
assign v$B_14426_out0 = v$SEL3_9047_out0;
assign v$B_14427_out0 = v$SEL2_17438_out0;
assign v$B_14430_out0 = v$SEL3_9048_out0;
assign v$B_14431_out0 = v$SEL2_17439_out0;
assign v$B_14446_out0 = v$SEL3_9052_out0;
assign v$B_14447_out0 = v$SEL2_17443_out0;
assign v$B_14450_out0 = v$SEL3_9053_out0;
assign v$B_14451_out0 = v$SEL2_17444_out0;
assign v$Clear_14641_out0 = v$Clear_12750_out0;
assign v$Clear_14642_out0 = v$Clear_12751_out0;
assign v$USELESS_15483_out0 = v$_7277_out0;
assign v$SEL2_15836_out0 = v$_7277_out1[1:1];
assign v$SEL4_16422_out0 = v$_7277_out1[3:3];
assign v$B2_16624_out0 = v$SEL8_12914_out0;
assign v$B2_16627_out0 = v$SEL8_12917_out0;
assign v$B2_16639_out0 = v$SEL8_12929_out0;
assign v$B2_16642_out0 = v$SEL8_12932_out0;
assign v$SEL7_17010_out0 = v$_7277_out1[6:6];
assign v$G3_17692_out0 = ! v$R_1588_out0;
assign v$G3_17693_out0 = ! v$R_1589_out0;
assign v$B3_17850_out0 = v$SEL7_4166_out0;
assign v$B3_17853_out0 = v$SEL7_4169_out0;
assign v$B3_17865_out0 = v$SEL7_4181_out0;
assign v$B3_17868_out0 = v$SEL7_4184_out0;
assign v$G18_18097_out0 = v$WREN_2534_out0 || v$G19_8261_out0;
assign v$G18_18098_out0 = v$WREN_2535_out0 || v$G19_8262_out0;
assign v$R_18338_out0 = v$RXreset_5959_out0;
assign v$R_18349_out0 = v$RXreset_5960_out0;
assign v$SAME_18736_out0 = v$G1_9389_out0;
assign v$SAME_18740_out0 = v$G1_9390_out0;
assign v$G32_398_out0 = v$A1$COMP$B1_12492_out0 || v$A0$COMP$B0_7992_out0;
assign v$G32_413_out0 = v$A1$COMP$B1_12507_out0 || v$A0$COMP$B0_8007_out0;
assign v$_1553_out0 = v$IN_9568_out0[15:15];
assign v$_1554_out0 = v$IN_9572_out0[15:15];
assign v$A2$COMP$B2_1979_out0 = v$G13_4406_out0;
assign v$A2$COMP$B2_1980_out0 = v$G13_4407_out0;
assign v$A2$COMP$B2_1994_out0 = v$G13_4421_out0;
assign v$A2$COMP$B2_1995_out0 = v$G13_4422_out0;
assign v$G21_3522_out0 = ! v$B1_14220_out0;
assign v$G21_3525_out0 = ! v$B1_14223_out0;
assign v$G21_3537_out0 = ! v$B1_14235_out0;
assign v$G21_3540_out0 = ! v$B1_14238_out0;
assign v$G8_3726_out0 = !((v$A3_10702_out0 && !v$B3_17850_out0) || (!v$A3_10702_out0) && v$B3_17850_out0);
assign v$G8_3729_out0 = !((v$A3_10705_out0 && !v$B3_17853_out0) || (!v$A3_10705_out0) && v$B3_17853_out0);
assign v$G8_3741_out0 = !((v$A3_10717_out0 && !v$B3_17865_out0) || (!v$A3_10717_out0) && v$B3_17865_out0);
assign v$G8_3744_out0 = !((v$A3_10720_out0 && !v$B3_17868_out0) || (!v$A3_10720_out0) && v$B3_17868_out0);
assign v$OUT_3922_out0 = v$G29_10300_out0;
assign v$SEL7_4167_out0 = v$B_14426_out0[3:3];
assign v$SEL7_4168_out0 = v$B_14427_out0[3:3];
assign v$SEL7_4170_out0 = v$B_14430_out0[3:3];
assign v$SEL7_4171_out0 = v$B_14431_out0[3:3];
assign v$SEL7_4182_out0 = v$B_14446_out0[3:3];
assign v$SEL7_4183_out0 = v$B_14447_out0[3:3];
assign v$SEL7_4185_out0 = v$B_14450_out0[3:3];
assign v$SEL7_4186_out0 = v$B_14451_out0[3:3];
assign v$G27_4783_out0 = v$A2XNORB2_4497_out0 && v$G28_13022_out0;
assign v$G27_4784_out0 = v$A2XNORB2_4498_out0 && v$G28_13023_out0;
assign v$G27_4798_out0 = v$A2XNORB2_4512_out0 && v$G28_13037_out0;
assign v$G27_4799_out0 = v$A2XNORB2_4513_out0 && v$G28_13038_out0;
assign v$_4802_out0 = v$IN_9568_out0[11:0];
assign v$_4806_out0 = v$IN_9572_out0[11:0];
assign v$G18_4980_out0 = v$A3XNORB3_14723_out0 && v$G22_13334_out0;
assign v$G18_4981_out0 = v$A3XNORB3_14724_out0 && v$G22_13335_out0;
assign v$G18_4995_out0 = v$A3XNORB3_14738_out0 && v$G22_13349_out0;
assign v$G18_4996_out0 = v$A3XNORB3_14739_out0 && v$G22_13350_out0;
assign v$G3_5001_out0 = v$SEL5_11625_out0 && v$SEL6_14244_out0;
assign v$G36_5906_out0 = !((v$B3_17850_out0 && !v$A3_10702_out0) || (!v$B3_17850_out0) && v$A3_10702_out0);
assign v$G36_5909_out0 = !((v$B3_17853_out0 && !v$A3_10705_out0) || (!v$B3_17853_out0) && v$A3_10705_out0);
assign v$G36_5921_out0 = !((v$B3_17865_out0 && !v$A3_10717_out0) || (!v$B3_17865_out0) && v$A3_10717_out0);
assign v$G36_5924_out0 = !((v$B3_17868_out0 && !v$A3_10720_out0) || (!v$B3_17868_out0) && v$A3_10720_out0);
assign v$G4_6417_out0 = v$SEL7_17010_out0 && v$SEL8_1968_out0;
assign v$G6_6549_out0 = ! v$B3_17850_out0;
assign v$G6_6552_out0 = ! v$B3_17853_out0;
assign v$G6_6564_out0 = ! v$B3_17865_out0;
assign v$G6_6567_out0 = ! v$B3_17868_out0;
assign v$_7378_out0 = v$IN_9568_out0[3:0];
assign v$_7379_out0 = v$IN_9572_out0[3:0];
assign v$ShiftEN_7722_out0 = v$G18_18097_out0;
assign v$ShiftEN_7723_out0 = v$G18_18098_out0;
assign v$G17_8178_out0 = !((v$A0_1725_out0 && !v$B0_3645_out0) || (!v$A0_1725_out0) && v$B0_3645_out0);
assign v$G17_8181_out0 = !((v$A0_1728_out0 && !v$B0_3648_out0) || (!v$A0_1728_out0) && v$B0_3648_out0);
assign v$G17_8193_out0 = !((v$A0_1740_out0 && !v$B0_3660_out0) || (!v$A0_1740_out0) && v$B0_3660_out0);
assign v$G17_8196_out0 = !((v$A0_1743_out0 && !v$B0_3663_out0) || (!v$A0_1743_out0) && v$B0_3663_out0);
assign v$G9_8671_out0 = v$TXSet_12652_out0 && v$TXLast_11385_out0;
assign v$G9_8672_out0 = v$TXSet_12653_out0 && v$TXLast_11386_out0;
assign v$G17_8894_out0 = ! v$WREN_10997_out0;
assign v$G17_8895_out0 = ! v$WREN_10998_out0;
assign v$SEL9_10838_out0 = v$B_14426_out0[1:1];
assign v$SEL9_10839_out0 = v$B_14427_out0[1:1];
assign v$SEL9_10841_out0 = v$B_14430_out0[1:1];
assign v$SEL9_10842_out0 = v$B_14431_out0[1:1];
assign v$SEL9_10853_out0 = v$B_14446_out0[1:1];
assign v$SEL9_10854_out0 = v$B_14447_out0[1:1];
assign v$SEL9_10856_out0 = v$B_14450_out0[1:1];
assign v$SEL9_10857_out0 = v$B_14451_out0[1:1];
assign v$G2_11697_out0 = v$SEL3_3126_out0 && v$SEL4_16422_out0;
assign v$G23_12175_out0 = ! v$B0_3645_out0;
assign v$G23_12178_out0 = ! v$B0_3648_out0;
assign v$G23_12190_out0 = ! v$B0_3660_out0;
assign v$G23_12193_out0 = ! v$B0_3663_out0;
assign v$SEL10_12607_out0 = v$B_14426_out0[0:0];
assign v$SEL10_12608_out0 = v$B_14427_out0[0:0];
assign v$SEL10_12610_out0 = v$B_14430_out0[0:0];
assign v$SEL10_12611_out0 = v$B_14431_out0[0:0];
assign v$SEL10_12622_out0 = v$B_14446_out0[0:0];
assign v$SEL10_12623_out0 = v$B_14447_out0[0:0];
assign v$SEL10_12625_out0 = v$B_14450_out0[0:0];
assign v$SEL10_12626_out0 = v$B_14451_out0[0:0];
assign v$SEL8_12915_out0 = v$B_14426_out0[2:2];
assign v$SEL8_12916_out0 = v$B_14427_out0[2:2];
assign v$SEL8_12918_out0 = v$B_14430_out0[2:2];
assign v$SEL8_12919_out0 = v$B_14431_out0[2:2];
assign v$SEL8_12930_out0 = v$B_14446_out0[2:2];
assign v$SEL8_12931_out0 = v$B_14447_out0[2:2];
assign v$SEL8_12933_out0 = v$B_14450_out0[2:2];
assign v$SEL8_12934_out0 = v$B_14451_out0[2:2];
assign v$G1_12984_out0 = v$STATE_16015_out0 && v$G3_17692_out0;
assign v$G1_12985_out0 = v$STATE_16016_out0 && v$G3_17693_out0;
assign v$G33_13099_out0 = !((v$A0_1725_out0 && !v$B0_3645_out0) || (!v$A0_1725_out0) && v$B0_3645_out0);
assign v$G33_13102_out0 = !((v$A0_1728_out0 && !v$B0_3648_out0) || (!v$A0_1728_out0) && v$B0_3648_out0);
assign v$G33_13114_out0 = !((v$A0_1740_out0 && !v$B0_3660_out0) || (!v$A0_1740_out0) && v$B0_3660_out0);
assign v$G33_13117_out0 = !((v$A0_1743_out0 && !v$B0_3663_out0) || (!v$A0_1743_out0) && v$B0_3663_out0);
assign v$_13270_out0 = v$IN_9568_out0[3:0];
assign v$_13273_out0 = v$IN_9572_out0[3:0];
assign v$G15_13643_out0 = !((v$A2_8057_out0 && !v$B2_16624_out0) || (!v$A2_8057_out0) && v$B2_16624_out0);
assign v$G15_13646_out0 = !((v$A2_8060_out0 && !v$B2_16627_out0) || (!v$A2_8060_out0) && v$B2_16627_out0);
assign v$G15_13658_out0 = !((v$A2_8072_out0 && !v$B2_16639_out0) || (!v$A2_8072_out0) && v$B2_16639_out0);
assign v$G15_13661_out0 = !((v$A2_8075_out0 && !v$B2_16642_out0) || (!v$A2_8075_out0) && v$B2_16642_out0);
assign v$G1_14410_out0 = v$SEL1_7005_out0 && v$SEL2_15836_out0;
assign v$G35_14523_out0 = !((v$A2_8057_out0 && !v$B2_16624_out0) || (!v$A2_8057_out0) && v$B2_16624_out0);
assign v$G35_14526_out0 = !((v$A2_8060_out0 && !v$B2_16627_out0) || (!v$A2_8060_out0) && v$B2_16627_out0);
assign v$G35_14538_out0 = !((v$A2_8072_out0 && !v$B2_16639_out0) || (!v$A2_8072_out0) && v$B2_16639_out0);
assign v$G35_14541_out0 = !((v$A2_8075_out0 && !v$B2_16642_out0) || (!v$A2_8075_out0) && v$B2_16642_out0);
assign v$_14601_out0 = v$IN_9568_out0[15:4];
assign v$_14605_out0 = v$IN_9572_out0[15:4];
assign v$_14635_out0 = v$IN_9568_out0[15:4];
assign v$_14639_out0 = v$IN_9572_out0[15:4];
assign v$G31_15515_out0 = v$A2$COMP$B2_1981_out0 || v$G32_401_out0;
assign v$G31_15516_out0 = v$A2$COMP$B2_1982_out0 || v$G32_402_out0;
assign v$G31_15517_out0 = v$A2$COMP$B2_1983_out0 || v$G32_403_out0;
assign v$G31_15519_out0 = v$A2$COMP$B2_1985_out0 || v$G32_405_out0;
assign v$G31_15520_out0 = v$A2$COMP$B2_1986_out0 || v$G32_406_out0;
assign v$G6_15566_out0 = ! v$R_18338_out0;
assign v$G6_15577_out0 = ! v$R_18349_out0;
assign v$G12_16468_out0 = ! v$B2_16624_out0;
assign v$G12_16471_out0 = ! v$B2_16627_out0;
assign v$G12_16483_out0 = ! v$B2_16639_out0;
assign v$G12_16486_out0 = ! v$B2_16642_out0;
assign v$_16749_out0 = v$IN_9568_out0[15:4];
assign v$_16753_out0 = v$IN_9572_out0[15:4];
assign v$G16_16862_out0 = !((v$A1_14339_out0 && !v$B1_14220_out0) || (!v$A1_14339_out0) && v$B1_14220_out0);
assign v$G16_16865_out0 = !((v$A1_14342_out0 && !v$B1_14223_out0) || (!v$A1_14342_out0) && v$B1_14223_out0);
assign v$G16_16877_out0 = !((v$A1_14354_out0 && !v$B1_14235_out0) || (!v$A1_14354_out0) && v$B1_14235_out0);
assign v$G16_16880_out0 = !((v$A1_14357_out0 && !v$B1_14238_out0) || (!v$A1_14357_out0) && v$B1_14238_out0);
assign v$S_16936_out0 = v$TXSet_12652_out0;
assign v$S_16947_out0 = v$TXSet_12653_out0;
assign v$G34_17292_out0 = !((v$A1_14339_out0 && !v$B1_14220_out0) || (!v$A1_14339_out0) && v$B1_14220_out0);
assign v$G34_17295_out0 = !((v$A1_14342_out0 && !v$B1_14223_out0) || (!v$A1_14342_out0) && v$B1_14223_out0);
assign v$G34_17307_out0 = !((v$A1_14354_out0 && !v$B1_14235_out0) || (!v$A1_14354_out0) && v$B1_14235_out0);
assign v$G34_17310_out0 = !((v$A1_14357_out0 && !v$B1_14238_out0) || (!v$A1_14357_out0) && v$B1_14238_out0);
assign v$R_18339_out0 = v$Clear_14641_out0;
assign v$R_18340_out0 = v$Clear_14641_out0;
assign v$R_18341_out0 = v$Clear_14641_out0;
assign v$R_18350_out0 = v$Clear_14642_out0;
assign v$R_18351_out0 = v$Clear_14642_out0;
assign v$R_18352_out0 = v$Clear_14642_out0;
assign v$SAME_18366_out0 = v$SAME_18736_out0;
assign v$SAME_18368_out0 = v$SAME_18740_out0;
assign v$SAME_18733_out0 = v$G41_10879_out0;
assign v$SAME_18734_out0 = v$G41_10880_out0;
assign v$SAME_18753_out0 = v$G41_10894_out0;
assign v$SAME_18754_out0 = v$G41_10895_out0;
assign v$MUX1_416_out0 = v$G17_8894_out0 ? v$FF2_2951_out0 : v$_3486_out0;
assign v$MUX1_417_out0 = v$G17_8895_out0 ? v$FF2_2952_out0 : v$_3487_out0;
assign v$G5_1124_out0 = v$FF2_13046_out0 && v$G6_15566_out0;
assign v$G5_1129_out0 = v$FF2_13057_out0 && v$G6_15577_out0;
assign v$A0XNORB0_1432_out0 = v$G17_8178_out0;
assign v$A0XNORB0_1435_out0 = v$G17_8181_out0;
assign v$A0XNORB0_1447_out0 = v$G17_8193_out0;
assign v$A0XNORB0_1450_out0 = v$G17_8196_out0;
assign v$_1479_out0 = { v$C1_7973_out0,v$_4802_out0 };
assign v$_1483_out0 = { v$C1_7977_out0,v$_4806_out0 };
assign v$MUX8_1496_out0 = v$G17_8894_out0 ? v$C1_12852_out0 : v$_9372_out1;
assign v$MUX8_1497_out0 = v$G17_8895_out0 ? v$C1_12853_out0 : v$_9373_out1;
assign v$G30_1778_out0 = v$A3$COMP$B3_4954_out0 || v$G31_15515_out0;
assign v$G30_1779_out0 = v$A3$COMP$B3_4955_out0 || v$G31_15516_out0;
assign v$G30_1780_out0 = v$A3$COMP$B3_4956_out0 || v$G31_15517_out0;
assign v$G30_1782_out0 = v$A3$COMP$B3_4958_out0 || v$G31_15519_out0;
assign v$G30_1783_out0 = v$A3$COMP$B3_4959_out0 || v$G31_15520_out0;
assign v$MUX3_3395_out0 = v$OUT_3922_out0 ? v$A$EXP_288_out0 : v$B$EXP_16676_out0;
assign v$B0_3646_out0 = v$SEL10_12607_out0;
assign v$B0_3647_out0 = v$SEL10_12608_out0;
assign v$B0_3649_out0 = v$SEL10_12610_out0;
assign v$B0_3650_out0 = v$SEL10_12611_out0;
assign v$B0_3661_out0 = v$SEL10_12622_out0;
assign v$B0_3662_out0 = v$SEL10_12623_out0;
assign v$B0_3664_out0 = v$SEL10_12625_out0;
assign v$B0_3665_out0 = v$SEL10_12626_out0;
assign v$A2XNORB2_4490_out0 = v$G15_13643_out0;
assign v$A2XNORB2_4493_out0 = v$G15_13646_out0;
assign v$A2XNORB2_4505_out0 = v$G15_13658_out0;
assign v$A2XNORB2_4508_out0 = v$G15_13661_out0;
assign v$G5_5797_out0 = v$G1_14410_out0 && v$G2_11697_out0;
assign v$G5_6934_out0 = v$A3_10702_out0 && v$G6_6549_out0;
assign v$G5_6937_out0 = v$A3_10705_out0 && v$G6_6552_out0;
assign v$G5_6949_out0 = v$A3_10717_out0 && v$G6_6564_out0;
assign v$G5_6952_out0 = v$A3_10720_out0 && v$G6_6567_out0;
assign v$G38_7291_out0 = v$G33_13099_out0 && v$G34_17292_out0;
assign v$G38_7294_out0 = v$G33_13102_out0 && v$G34_17295_out0;
assign v$G38_7306_out0 = v$G33_13114_out0 && v$G34_17307_out0;
assign v$G38_7309_out0 = v$G33_13117_out0 && v$G34_17310_out0;
assign v$G2_7576_out0 = v$G1_12984_out0 || v$S_8019_out0;
assign v$G2_7577_out0 = v$G1_12985_out0 || v$S_8020_out0;
assign v$MUX6_9130_out0 = v$G17_8894_out0 ? v$FF7_18120_out0 : v$_8090_out1;
assign v$MUX6_9131_out0 = v$G17_8895_out0 ? v$FF7_18121_out0 : v$_8091_out1;
assign v$_9447_out0 = { v$_16749_out0,v$LSBS_15316_out0 };
assign v$_9451_out0 = { v$_16753_out0,v$LSBS_15317_out0 };
assign v$MUX7_9480_out0 = v$G17_8894_out0 ? v$FF8_8026_out0 : v$_9372_out0;
assign v$MUX7_9481_out0 = v$G17_8895_out0 ? v$FF8_8027_out0 : v$_9373_out0;
assign v$G20_9882_out0 = v$A1_14339_out0 && v$G21_3522_out0;
assign v$G20_9885_out0 = v$A1_14342_out0 && v$G21_3525_out0;
assign v$G20_9897_out0 = v$A1_14354_out0 && v$G21_3537_out0;
assign v$G20_9900_out0 = v$A1_14357_out0 && v$G21_3540_out0;
assign v$_9911_out0 = { v$_1553_out0,v$_1553_out0 };
assign v$_9912_out0 = { v$_1554_out0,v$_1554_out0 };
assign v$LOWER$SAME_10183_out0 = v$SAME_18734_out0;
assign v$LOWER$SAME_10188_out0 = v$SAME_18754_out0;
assign v$G25_10934_out0 = v$A0_1725_out0 && v$G23_12175_out0;
assign v$G25_10937_out0 = v$A0_1728_out0 && v$G23_12178_out0;
assign v$G25_10949_out0 = v$A0_1740_out0 && v$G23_12190_out0;
assign v$G25_10952_out0 = v$A0_1743_out0 && v$G23_12193_out0;
assign v$MUX4_11648_out0 = v$IS$32$BITS_2992_out0 ? v$SAME_18366_out0 : v$SAME_18365_out0;
assign v$MUX4_11649_out0 = v$IS$32$BITS_1282_out0 ? v$SAME_18368_out0 : v$SAME_18367_out0;
assign v$G4_11833_out0 = v$G5_1123_out0 || v$S_16936_out0;
assign v$G4_11838_out0 = v$G5_1128_out0 || v$S_16947_out0;
assign v$A1$COMP$B1_12493_out0 = v$G18_4980_out0;
assign v$A1$COMP$B1_12494_out0 = v$G18_4981_out0;
assign v$A1$COMP$B1_12508_out0 = v$G18_4995_out0;
assign v$A1$COMP$B1_12509_out0 = v$G18_4996_out0;
assign v$MUX2_13287_out0 = v$G17_8894_out0 ? v$FF3_262_out0 : v$_3486_out1;
assign v$MUX2_13288_out0 = v$G17_8895_out0 ? v$FF3_263_out0 : v$_3487_out1;
assign v$_13306_out0 = { v$_14601_out0,v$_13270_out0 };
assign v$_13310_out0 = { v$_14605_out0,v$_13273_out0 };
assign v$G40_13360_out0 = v$G35_14523_out0 && v$G36_5906_out0;
assign v$G40_13363_out0 = v$G35_14526_out0 && v$G36_5909_out0;
assign v$G40_13375_out0 = v$G35_14538_out0 && v$G36_5921_out0;
assign v$G40_13378_out0 = v$G35_14541_out0 && v$G36_5924_out0;
assign v$OUT_13760_out0 = v$OUT_3922_out0;
assign v$B1_14221_out0 = v$SEL9_10838_out0;
assign v$B1_14222_out0 = v$SEL9_10839_out0;
assign v$B1_14224_out0 = v$SEL9_10841_out0;
assign v$B1_14225_out0 = v$SEL9_10842_out0;
assign v$B1_14236_out0 = v$SEL9_10853_out0;
assign v$B1_14237_out0 = v$SEL9_10854_out0;
assign v$B1_14239_out0 = v$SEL9_10856_out0;
assign v$B1_14240_out0 = v$SEL9_10857_out0;
assign v$MUX5_14489_out0 = v$S_10347_out0 ? v$_7378_out0 : v$C1_12825_out0;
assign v$MUX5_14490_out0 = v$S_10348_out0 ? v$_7379_out0 : v$C1_12826_out0;
assign v$A3XNORB3_14716_out0 = v$G8_3726_out0;
assign v$A3XNORB3_14719_out0 = v$G8_3729_out0;
assign v$A3XNORB3_14731_out0 = v$G8_3741_out0;
assign v$A3XNORB3_14734_out0 = v$G8_3744_out0;
assign v$HIGHER$SAME_15022_out0 = v$SAME_18733_out0;
assign v$HIGHER$SAME_15027_out0 = v$SAME_18753_out0;
assign v$G31_15512_out0 = v$A2$COMP$B2_1978_out0 || v$G32_398_out0;
assign v$G31_15527_out0 = v$A2$COMP$B2_1993_out0 || v$G32_413_out0;
assign v$G6_15567_out0 = ! v$R_18339_out0;
assign v$G6_15568_out0 = ! v$R_18340_out0;
assign v$G6_15569_out0 = ! v$R_18341_out0;
assign v$G6_15578_out0 = ! v$R_18350_out0;
assign v$G6_15579_out0 = ! v$R_18351_out0;
assign v$G6_15580_out0 = ! v$R_18352_out0;
assign v$MUX4_15635_out0 = v$G17_8894_out0 ? v$FF5_16338_out0 : v$_14078_out1;
assign v$MUX4_15636_out0 = v$G17_8895_out0 ? v$FF5_16339_out0 : v$_14079_out1;
assign v$G11_15637_out0 = v$A2_8057_out0 && v$G12_16468_out0;
assign v$G11_15640_out0 = v$A2_8060_out0 && v$G12_16471_out0;
assign v$G11_15652_out0 = v$A2_8072_out0 && v$G12_16483_out0;
assign v$G11_15655_out0 = v$A2_8075_out0 && v$G12_16486_out0;
assign v$G24_15691_out0 = v$A3XNORB3_14723_out0 && v$G27_4783_out0;
assign v$G24_15692_out0 = v$A3XNORB3_14724_out0 && v$G27_4784_out0;
assign v$G24_15706_out0 = v$A3XNORB3_14738_out0 && v$G27_4798_out0;
assign v$G24_15707_out0 = v$A3XNORB3_14739_out0 && v$G27_4799_out0;
assign v$A1XNORB1_16045_out0 = v$G16_16862_out0;
assign v$A1XNORB1_16048_out0 = v$G16_16865_out0;
assign v$A1XNORB1_16060_out0 = v$G16_16877_out0;
assign v$A1XNORB1_16063_out0 = v$G16_16880_out0;
assign v$B2_16625_out0 = v$SEL8_12915_out0;
assign v$B2_16626_out0 = v$SEL8_12916_out0;
assign v$B2_16628_out0 = v$SEL8_12918_out0;
assign v$B2_16629_out0 = v$SEL8_12919_out0;
assign v$B2_16640_out0 = v$SEL8_12930_out0;
assign v$B2_16641_out0 = v$SEL8_12931_out0;
assign v$B2_16643_out0 = v$SEL8_12933_out0;
assign v$B2_16644_out0 = v$SEL8_12934_out0;
assign v$S_16938_out0 = v$G9_8671_out0;
assign v$S_16949_out0 = v$G9_8672_out0;
assign v$G6_17398_out0 = v$G3_5001_out0 && v$G4_6417_out0;
assign v$MUX3_17725_out0 = v$G17_8894_out0 ? v$FF4_2347_out0 : v$_14078_out0;
assign v$MUX3_17726_out0 = v$G17_8895_out0 ? v$FF4_2348_out0 : v$_14079_out0;
assign v$B3_17851_out0 = v$SEL7_4167_out0;
assign v$B3_17852_out0 = v$SEL7_4168_out0;
assign v$B3_17854_out0 = v$SEL7_4170_out0;
assign v$B3_17855_out0 = v$SEL7_4171_out0;
assign v$B3_17866_out0 = v$SEL7_4182_out0;
assign v$B3_17867_out0 = v$SEL7_4183_out0;
assign v$B3_17869_out0 = v$SEL7_4185_out0;
assign v$B3_17870_out0 = v$SEL7_4186_out0;
assign v$MUX1_17927_out0 = v$OUT_3922_out0 ? v$B$EXP_16676_out0 : v$A$EXP_288_out0;
assign v$MUX5_18559_out0 = v$G17_8894_out0 ? v$FF6_15324_out0 : v$_8090_out0;
assign v$MUX5_18560_out0 = v$G17_8895_out0 ? v$FF6_15325_out0 : v$_8091_out0;
assign v$G5_1125_out0 = v$FF2_13047_out0 && v$G6_15567_out0;
assign v$G5_1126_out0 = v$FF2_13048_out0 && v$G6_15568_out0;
assign v$G5_1127_out0 = v$FF2_13049_out0 && v$G6_15569_out0;
assign v$G5_1130_out0 = v$FF2_13058_out0 && v$G6_15578_out0;
assign v$G5_1131_out0 = v$FF2_13059_out0 && v$G6_15579_out0;
assign v$G5_1132_out0 = v$FF2_13060_out0 && v$G6_15580_out0;
assign v$G30_1775_out0 = v$A3$COMP$B3_4951_out0 || v$G31_15512_out0;
assign v$G30_1790_out0 = v$A3$COMP$B3_4966_out0 || v$G31_15527_out0;
assign v$G21_3523_out0 = ! v$B1_14221_out0;
assign v$G21_3524_out0 = ! v$B1_14222_out0;
assign v$G21_3526_out0 = ! v$B1_14224_out0;
assign v$G21_3527_out0 = ! v$B1_14225_out0;
assign v$G21_3538_out0 = ! v$B1_14236_out0;
assign v$G21_3539_out0 = ! v$B1_14237_out0;
assign v$G21_3541_out0 = ! v$B1_14239_out0;
assign v$G21_3542_out0 = ! v$B1_14240_out0;
assign v$G8_3727_out0 = !((v$A3_10703_out0 && !v$B3_17851_out0) || (!v$A3_10703_out0) && v$B3_17851_out0);
assign v$G8_3728_out0 = !((v$A3_10704_out0 && !v$B3_17852_out0) || (!v$A3_10704_out0) && v$B3_17852_out0);
assign v$G8_3730_out0 = !((v$A3_10706_out0 && !v$B3_17854_out0) || (!v$A3_10706_out0) && v$B3_17854_out0);
assign v$G8_3731_out0 = !((v$A3_10707_out0 && !v$B3_17855_out0) || (!v$A3_10707_out0) && v$B3_17855_out0);
assign v$G8_3742_out0 = !((v$A3_10718_out0 && !v$B3_17866_out0) || (!v$A3_10718_out0) && v$B3_17866_out0);
assign v$G8_3743_out0 = !((v$A3_10719_out0 && !v$B3_17867_out0) || (!v$A3_10719_out0) && v$B3_17867_out0);
assign v$G8_3745_out0 = !((v$A3_10721_out0 && !v$B3_17869_out0) || (!v$A3_10721_out0) && v$B3_17869_out0);
assign v$G8_3746_out0 = !((v$A3_10722_out0 && !v$B3_17870_out0) || (!v$A3_10722_out0) && v$B3_17870_out0);
assign v$OUT_3920_out0 = v$G30_1779_out0;
assign v$OUT_3921_out0 = v$G30_1780_out0;
assign v$OUT_3924_out0 = v$G30_1782_out0;
assign v$OUT_3925_out0 = v$G30_1783_out0;
assign v$G13_4399_out0 = v$A3XNORB3_14716_out0 && v$G11_15637_out0;
assign v$G13_4402_out0 = v$A3XNORB3_14719_out0 && v$G11_15640_out0;
assign v$G13_4414_out0 = v$A3XNORB3_14731_out0 && v$G11_15652_out0;
assign v$G13_4417_out0 = v$A3XNORB3_14734_out0 && v$G11_15655_out0;
assign v$A3$COMP$B3_4945_out0 = v$G5_6934_out0;
assign v$A3$COMP$B3_4948_out0 = v$G5_6937_out0;
assign v$A3$COMP$B3_4960_out0 = v$G5_6949_out0;
assign v$A3$COMP$B3_4963_out0 = v$G5_6952_out0;
assign v$G36_5907_out0 = !((v$B3_17851_out0 && !v$A3_10703_out0) || (!v$B3_17851_out0) && v$A3_10703_out0);
assign v$G36_5908_out0 = !((v$B3_17852_out0 && !v$A3_10704_out0) || (!v$B3_17852_out0) && v$A3_10704_out0);
assign v$G36_5910_out0 = !((v$B3_17854_out0 && !v$A3_10706_out0) || (!v$B3_17854_out0) && v$A3_10706_out0);
assign v$G36_5911_out0 = !((v$B3_17855_out0 && !v$A3_10707_out0) || (!v$B3_17855_out0) && v$A3_10707_out0);
assign v$G36_5922_out0 = !((v$B3_17866_out0 && !v$A3_10718_out0) || (!v$B3_17866_out0) && v$A3_10718_out0);
assign v$G36_5923_out0 = !((v$B3_17867_out0 && !v$A3_10719_out0) || (!v$B3_17867_out0) && v$A3_10719_out0);
assign v$G36_5925_out0 = !((v$B3_17869_out0 && !v$A3_10721_out0) || (!v$B3_17869_out0) && v$A3_10721_out0);
assign v$G36_5926_out0 = !((v$B3_17870_out0 && !v$A3_10722_out0) || (!v$B3_17870_out0) && v$A3_10722_out0);
assign v$G6_6550_out0 = ! v$B3_17851_out0;
assign v$G6_6551_out0 = ! v$B3_17852_out0;
assign v$G6_6553_out0 = ! v$B3_17854_out0;
assign v$G6_6554_out0 = ! v$B3_17855_out0;
assign v$G6_6565_out0 = ! v$B3_17866_out0;
assign v$G6_6566_out0 = ! v$B3_17867_out0;
assign v$G6_6568_out0 = ! v$B3_17869_out0;
assign v$G6_6569_out0 = ! v$B3_17870_out0;
assign v$_7550_out0 = { v$_9911_out0,v$_9911_out0 };
assign v$_7551_out0 = { v$_9912_out0,v$_9912_out0 };
assign v$XOR1_7593_out0 = v$C1_13578_out0 ^ v$MUX1_17927_out0;
assign v$A0$COMP$B0_7993_out0 = v$G24_15691_out0;
assign v$A0$COMP$B0_7994_out0 = v$G24_15692_out0;
assign v$A0$COMP$B0_8008_out0 = v$G24_15706_out0;
assign v$A0$COMP$B0_8009_out0 = v$G24_15707_out0;
assign v$G17_8179_out0 = !((v$A0_1726_out0 && !v$B0_3646_out0) || (!v$A0_1726_out0) && v$B0_3646_out0);
assign v$G17_8180_out0 = !((v$A0_1727_out0 && !v$B0_3647_out0) || (!v$A0_1727_out0) && v$B0_3647_out0);
assign v$G17_8182_out0 = !((v$A0_1729_out0 && !v$B0_3649_out0) || (!v$A0_1729_out0) && v$B0_3649_out0);
assign v$G17_8183_out0 = !((v$A0_1730_out0 && !v$B0_3650_out0) || (!v$A0_1730_out0) && v$B0_3650_out0);
assign v$G17_8194_out0 = !((v$A0_1741_out0 && !v$B0_3661_out0) || (!v$A0_1741_out0) && v$B0_3661_out0);
assign v$G17_8195_out0 = !((v$A0_1742_out0 && !v$B0_3662_out0) || (!v$A0_1742_out0) && v$B0_3662_out0);
assign v$G17_8197_out0 = !((v$A0_1744_out0 && !v$B0_3664_out0) || (!v$A0_1744_out0) && v$B0_3664_out0);
assign v$G17_8198_out0 = !((v$A0_1745_out0 && !v$B0_3665_out0) || (!v$A0_1745_out0) && v$B0_3665_out0);
assign v$G1_9388_out0 = v$LOWER$SAME_10183_out0 && v$HIGHER$SAME_15022_out0;
assign v$G1_9393_out0 = v$LOWER$SAME_10188_out0 && v$HIGHER$SAME_15027_out0;
assign v$G29_10299_out0 = v$A4$COMP$B4_7410_out0 || v$G30_1778_out0;
assign v$G41_10872_out0 = v$G38_7291_out0 && v$G40_13360_out0;
assign v$G41_10875_out0 = v$G38_7294_out0 && v$G40_13363_out0;
assign v$G41_10887_out0 = v$G38_7306_out0 && v$G40_13375_out0;
assign v$G41_10890_out0 = v$G38_7309_out0 && v$G40_13378_out0;
assign v$G4_11834_out0 = v$G5_1124_out0 || v$S_16937_out0;
assign v$G4_11839_out0 = v$G5_1129_out0 || v$S_16948_out0;
assign v$G23_12176_out0 = ! v$B0_3646_out0;
assign v$G23_12177_out0 = ! v$B0_3647_out0;
assign v$G23_12179_out0 = ! v$B0_3649_out0;
assign v$G23_12180_out0 = ! v$B0_3650_out0;
assign v$G23_12191_out0 = ! v$B0_3661_out0;
assign v$G23_12192_out0 = ! v$B0_3662_out0;
assign v$G23_12194_out0 = ! v$B0_3664_out0;
assign v$G23_12195_out0 = ! v$B0_3665_out0;
assign v$G28_13015_out0 = v$A1XNORB1_16045_out0 && v$G25_10934_out0;
assign v$G28_13018_out0 = v$A1XNORB1_16048_out0 && v$G25_10937_out0;
assign v$G28_13030_out0 = v$A1XNORB1_16060_out0 && v$G25_10949_out0;
assign v$G28_13033_out0 = v$A1XNORB1_16063_out0 && v$G25_10952_out0;
assign v$G33_13100_out0 = !((v$A0_1726_out0 && !v$B0_3646_out0) || (!v$A0_1726_out0) && v$B0_3646_out0);
assign v$G33_13101_out0 = !((v$A0_1727_out0 && !v$B0_3647_out0) || (!v$A0_1727_out0) && v$B0_3647_out0);
assign v$G33_13103_out0 = !((v$A0_1729_out0 && !v$B0_3649_out0) || (!v$A0_1729_out0) && v$B0_3649_out0);
assign v$G33_13104_out0 = !((v$A0_1730_out0 && !v$B0_3650_out0) || (!v$A0_1730_out0) && v$B0_3650_out0);
assign v$G33_13115_out0 = !((v$A0_1741_out0 && !v$B0_3661_out0) || (!v$A0_1741_out0) && v$B0_3661_out0);
assign v$G33_13116_out0 = !((v$A0_1742_out0 && !v$B0_3662_out0) || (!v$A0_1742_out0) && v$B0_3662_out0);
assign v$G33_13118_out0 = !((v$A0_1744_out0 && !v$B0_3664_out0) || (!v$A0_1744_out0) && v$B0_3664_out0);
assign v$G33_13119_out0 = !((v$A0_1745_out0 && !v$B0_3665_out0) || (!v$A0_1745_out0) && v$B0_3665_out0);
assign v$G22_13327_out0 = v$A2XNORB2_4490_out0 && v$G20_9882_out0;
assign v$G22_13330_out0 = v$A2XNORB2_4493_out0 && v$G20_9885_out0;
assign v$G22_13342_out0 = v$A2XNORB2_4505_out0 && v$G20_9897_out0;
assign v$G22_13345_out0 = v$A2XNORB2_4508_out0 && v$G20_9900_out0;
assign v$NEXTSTATE_13537_out0 = v$G2_7576_out0;
assign v$NEXTSTATE_13538_out0 = v$G2_7577_out0;
assign v$G15_13644_out0 = !((v$A2_8058_out0 && !v$B2_16625_out0) || (!v$A2_8058_out0) && v$B2_16625_out0);
assign v$G15_13645_out0 = !((v$A2_8059_out0 && !v$B2_16626_out0) || (!v$A2_8059_out0) && v$B2_16626_out0);
assign v$G15_13647_out0 = !((v$A2_8061_out0 && !v$B2_16628_out0) || (!v$A2_8061_out0) && v$B2_16628_out0);
assign v$G15_13648_out0 = !((v$A2_8062_out0 && !v$B2_16629_out0) || (!v$A2_8062_out0) && v$B2_16629_out0);
assign v$G15_13659_out0 = !((v$A2_8073_out0 && !v$B2_16640_out0) || (!v$A2_8073_out0) && v$B2_16640_out0);
assign v$G15_13660_out0 = !((v$A2_8074_out0 && !v$B2_16641_out0) || (!v$A2_8074_out0) && v$B2_16641_out0);
assign v$G15_13662_out0 = !((v$A2_8076_out0 && !v$B2_16643_out0) || (!v$A2_8076_out0) && v$B2_16643_out0);
assign v$G15_13663_out0 = !((v$A2_8077_out0 && !v$B2_16644_out0) || (!v$A2_8077_out0) && v$B2_16644_out0);
assign v$Q_14146_out0 = v$G4_11833_out0;
assign v$Q_14157_out0 = v$G4_11838_out0;
assign v$G35_14524_out0 = !((v$A2_8058_out0 && !v$B2_16625_out0) || (!v$A2_8058_out0) && v$B2_16625_out0);
assign v$G35_14525_out0 = !((v$A2_8059_out0 && !v$B2_16626_out0) || (!v$A2_8059_out0) && v$B2_16626_out0);
assign v$G35_14527_out0 = !((v$A2_8061_out0 && !v$B2_16628_out0) || (!v$A2_8061_out0) && v$B2_16628_out0);
assign v$G35_14528_out0 = !((v$A2_8062_out0 && !v$B2_16629_out0) || (!v$A2_8062_out0) && v$B2_16629_out0);
assign v$G35_14539_out0 = !((v$A2_8073_out0 && !v$B2_16640_out0) || (!v$A2_8073_out0) && v$B2_16640_out0);
assign v$G35_14540_out0 = !((v$A2_8074_out0 && !v$B2_16641_out0) || (!v$A2_8074_out0) && v$B2_16641_out0);
assign v$G35_14542_out0 = !((v$A2_8076_out0 && !v$B2_16643_out0) || (!v$A2_8076_out0) && v$B2_16643_out0);
assign v$G35_14543_out0 = !((v$A2_8077_out0 && !v$B2_16644_out0) || (!v$A2_8077_out0) && v$B2_16644_out0);
assign v$G7_14806_out0 = v$G5_5797_out0 && v$G6_17398_out0;
assign v$MUX4_15992_out0 = v$EN_16967_out0 ? v$_1479_out0 : v$IN_9568_out0;
assign v$MUX4_15996_out0 = v$EN_16971_out0 ? v$_1483_out0 : v$IN_9572_out0;
assign v$G12_16469_out0 = ! v$B2_16625_out0;
assign v$G12_16470_out0 = ! v$B2_16626_out0;
assign v$G12_16472_out0 = ! v$B2_16628_out0;
assign v$G12_16473_out0 = ! v$B2_16629_out0;
assign v$G12_16484_out0 = ! v$B2_16640_out0;
assign v$G12_16485_out0 = ! v$B2_16641_out0;
assign v$G12_16487_out0 = ! v$B2_16643_out0;
assign v$G12_16488_out0 = ! v$B2_16644_out0;
assign v$EXP$SAME_16546_out0 = v$MUX4_11648_out0;
assign v$EXP$SAME_16547_out0 = v$MUX4_11649_out0;
assign v$G16_16863_out0 = !((v$A1_14340_out0 && !v$B1_14221_out0) || (!v$A1_14340_out0) && v$B1_14221_out0);
assign v$G16_16864_out0 = !((v$A1_14341_out0 && !v$B1_14222_out0) || (!v$A1_14341_out0) && v$B1_14222_out0);
assign v$G16_16866_out0 = !((v$A1_14343_out0 && !v$B1_14224_out0) || (!v$A1_14343_out0) && v$B1_14224_out0);
assign v$G16_16867_out0 = !((v$A1_14344_out0 && !v$B1_14225_out0) || (!v$A1_14344_out0) && v$B1_14225_out0);
assign v$G16_16878_out0 = !((v$A1_14355_out0 && !v$B1_14236_out0) || (!v$A1_14355_out0) && v$B1_14236_out0);
assign v$G16_16879_out0 = !((v$A1_14356_out0 && !v$B1_14237_out0) || (!v$A1_14356_out0) && v$B1_14237_out0);
assign v$G16_16881_out0 = !((v$A1_14358_out0 && !v$B1_14239_out0) || (!v$A1_14358_out0) && v$B1_14239_out0);
assign v$G16_16882_out0 = !((v$A1_14359_out0 && !v$B1_14240_out0) || (!v$A1_14359_out0) && v$B1_14240_out0);
assign v$G34_17293_out0 = !((v$A1_14340_out0 && !v$B1_14221_out0) || (!v$A1_14340_out0) && v$B1_14221_out0);
assign v$G34_17294_out0 = !((v$A1_14341_out0 && !v$B1_14222_out0) || (!v$A1_14341_out0) && v$B1_14222_out0);
assign v$G34_17296_out0 = !((v$A1_14343_out0 && !v$B1_14224_out0) || (!v$A1_14343_out0) && v$B1_14224_out0);
assign v$G34_17297_out0 = !((v$A1_14344_out0 && !v$B1_14225_out0) || (!v$A1_14344_out0) && v$B1_14225_out0);
assign v$G34_17308_out0 = !((v$A1_14355_out0 && !v$B1_14236_out0) || (!v$A1_14355_out0) && v$B1_14236_out0);
assign v$G34_17309_out0 = !((v$A1_14356_out0 && !v$B1_14237_out0) || (!v$A1_14356_out0) && v$B1_14237_out0);
assign v$G34_17311_out0 = !((v$A1_14358_out0 && !v$B1_14239_out0) || (!v$A1_14358_out0) && v$B1_14239_out0);
assign v$G34_17312_out0 = !((v$A1_14359_out0 && !v$B1_14240_out0) || (!v$A1_14359_out0) && v$B1_14240_out0);
assign v$G32_399_out0 = v$A1$COMP$B1_12493_out0 || v$A0$COMP$B0_7993_out0;
assign v$G32_400_out0 = v$A1$COMP$B1_12494_out0 || v$A0$COMP$B0_7994_out0;
assign v$G32_414_out0 = v$A1$COMP$B1_12508_out0 || v$A0$COMP$B0_8008_out0;
assign v$G32_415_out0 = v$A1$COMP$B1_12509_out0 || v$A0$COMP$B0_8009_out0;
assign v$A0XNORB0_1433_out0 = v$G17_8179_out0;
assign v$A0XNORB0_1434_out0 = v$G17_8180_out0;
assign v$A0XNORB0_1436_out0 = v$G17_8182_out0;
assign v$A0XNORB0_1437_out0 = v$G17_8183_out0;
assign v$A0XNORB0_1448_out0 = v$G17_8194_out0;
assign v$A0XNORB0_1449_out0 = v$G17_8195_out0;
assign v$A0XNORB0_1451_out0 = v$G17_8197_out0;
assign v$A0XNORB0_1452_out0 = v$G17_8198_out0;
assign v$A2$COMP$B2_1972_out0 = v$G13_4399_out0;
assign v$A2$COMP$B2_1975_out0 = v$G13_4402_out0;
assign v$A2$COMP$B2_1987_out0 = v$G13_4414_out0;
assign v$A2$COMP$B2_1990_out0 = v$G13_4417_out0;
assign v$MUX6_2847_out0 = v$FF1_13680_out0 ? v$LSBS_15316_out0 : v$_7550_out0;
assign v$MUX6_2848_out0 = v$FF1_13681_out0 ? v$LSBS_15317_out0 : v$_7551_out0;
assign v$HIGHER$OUT_3832_out0 = v$OUT_3920_out0;
assign v$HIGHER$OUT_3833_out0 = v$OUT_3924_out0;
assign v$OUT_3918_out0 = v$G29_10299_out0;
assign v$LOWER$OUT_4224_out0 = v$OUT_3921_out0;
assign v$LOWER$OUT_4225_out0 = v$OUT_3925_out0;
assign v$A2XNORB2_4491_out0 = v$G15_13644_out0;
assign v$A2XNORB2_4492_out0 = v$G15_13645_out0;
assign v$A2XNORB2_4494_out0 = v$G15_13647_out0;
assign v$A2XNORB2_4495_out0 = v$G15_13648_out0;
assign v$A2XNORB2_4506_out0 = v$G15_13659_out0;
assign v$A2XNORB2_4507_out0 = v$G15_13660_out0;
assign v$A2XNORB2_4509_out0 = v$G15_13662_out0;
assign v$A2XNORB2_4510_out0 = v$G15_13663_out0;
assign v$G27_4776_out0 = v$A2XNORB2_4490_out0 && v$G28_13015_out0;
assign v$G27_4779_out0 = v$A2XNORB2_4493_out0 && v$G28_13018_out0;
assign v$G27_4791_out0 = v$A2XNORB2_4505_out0 && v$G28_13030_out0;
assign v$G27_4794_out0 = v$A2XNORB2_4508_out0 && v$G28_13033_out0;
assign v$G18_4973_out0 = v$A3XNORB3_14716_out0 && v$G22_13327_out0;
assign v$G18_4976_out0 = v$A3XNORB3_14719_out0 && v$G22_13330_out0;
assign v$G18_4988_out0 = v$A3XNORB3_14731_out0 && v$G22_13342_out0;
assign v$G18_4991_out0 = v$A3XNORB3_14734_out0 && v$G22_13345_out0;
assign {v$A1_5793_out1,v$A1_5793_out0 } = v$MUX3_3395_out0 + v$XOR1_7593_out0 + v$CIN_18229_out0;
assign v$G5_6935_out0 = v$A3_10703_out0 && v$G6_6550_out0;
assign v$G5_6936_out0 = v$A3_10704_out0 && v$G6_6551_out0;
assign v$G5_6938_out0 = v$A3_10706_out0 && v$G6_6553_out0;
assign v$G5_6939_out0 = v$A3_10707_out0 && v$G6_6554_out0;
assign v$G5_6950_out0 = v$A3_10718_out0 && v$G6_6565_out0;
assign v$G5_6951_out0 = v$A3_10719_out0 && v$G6_6566_out0;
assign v$G5_6953_out0 = v$A3_10721_out0 && v$G6_6568_out0;
assign v$G5_6954_out0 = v$A3_10722_out0 && v$G6_6569_out0;
assign v$G38_7292_out0 = v$G33_13100_out0 && v$G34_17293_out0;
assign v$G38_7293_out0 = v$G33_13101_out0 && v$G34_17294_out0;
assign v$G38_7295_out0 = v$G33_13103_out0 && v$G34_17296_out0;
assign v$G38_7296_out0 = v$G33_13104_out0 && v$G34_17297_out0;
assign v$G38_7307_out0 = v$G33_13115_out0 && v$G34_17308_out0;
assign v$G38_7308_out0 = v$G33_13116_out0 && v$G34_17309_out0;
assign v$G38_7310_out0 = v$G33_13118_out0 && v$G34_17311_out0;
assign v$G38_7311_out0 = v$G33_13119_out0 && v$G34_17312_out0;
assign v$TXFlag_7718_out0 = v$Q_14146_out0;
assign v$TXFlag_7719_out0 = v$Q_14157_out0;
assign v$IGNORE_8283_out0 = v$G7_14806_out0;
assign v$G20_9883_out0 = v$A1_14340_out0 && v$G21_3523_out0;
assign v$G20_9884_out0 = v$A1_14341_out0 && v$G21_3524_out0;
assign v$G20_9886_out0 = v$A1_14343_out0 && v$G21_3526_out0;
assign v$G20_9887_out0 = v$A1_14344_out0 && v$G21_3527_out0;
assign v$G20_9898_out0 = v$A1_14355_out0 && v$G21_3538_out0;
assign v$G20_9899_out0 = v$A1_14356_out0 && v$G21_3539_out0;
assign v$G20_9901_out0 = v$A1_14358_out0 && v$G21_3541_out0;
assign v$G20_9902_out0 = v$A1_14359_out0 && v$G21_3542_out0;
assign v$G29_10298_out0 = v$A4$COMP$B4_7409_out0 || v$G30_1775_out0;
assign v$G29_10301_out0 = v$A4$COMP$B4_7412_out0 || v$G30_1790_out0;
assign v$G25_10935_out0 = v$A0_1726_out0 && v$G23_12176_out0;
assign v$G25_10936_out0 = v$A0_1727_out0 && v$G23_12177_out0;
assign v$G25_10938_out0 = v$A0_1729_out0 && v$G23_12179_out0;
assign v$G25_10939_out0 = v$A0_1730_out0 && v$G23_12180_out0;
assign v$G25_10950_out0 = v$A0_1741_out0 && v$G23_12191_out0;
assign v$G25_10951_out0 = v$A0_1742_out0 && v$G23_12192_out0;
assign v$G25_10953_out0 = v$A0_1744_out0 && v$G23_12194_out0;
assign v$G25_10954_out0 = v$A0_1745_out0 && v$G23_12195_out0;
assign v$G4_11835_out0 = v$G5_1125_out0 || v$S_16938_out0;
assign v$G4_11836_out0 = v$G5_1126_out0 || v$S_16939_out0;
assign v$G4_11837_out0 = v$G5_1127_out0 || v$S_16940_out0;
assign v$G4_11840_out0 = v$G5_1130_out0 || v$S_16949_out0;
assign v$G4_11841_out0 = v$G5_1131_out0 || v$S_16950_out0;
assign v$G4_11842_out0 = v$G5_1132_out0 || v$S_16951_out0;
assign v$MUX2_12040_out0 = v$G3_2607_out0 ? v$_9447_out0 : v$MUX4_15992_out0;
assign v$MUX2_12044_out0 = v$G3_2611_out0 ? v$_9451_out0 : v$MUX4_15996_out0;
assign v$G40_13361_out0 = v$G35_14524_out0 && v$G36_5907_out0;
assign v$G40_13362_out0 = v$G35_14525_out0 && v$G36_5908_out0;
assign v$G40_13364_out0 = v$G35_14527_out0 && v$G36_5910_out0;
assign v$G40_13365_out0 = v$G35_14528_out0 && v$G36_5911_out0;
assign v$G40_13376_out0 = v$G35_14539_out0 && v$G36_5922_out0;
assign v$G40_13377_out0 = v$G35_14540_out0 && v$G36_5923_out0;
assign v$G40_13379_out0 = v$G35_14542_out0 && v$G36_5925_out0;
assign v$G40_13380_out0 = v$G35_14543_out0 && v$G36_5926_out0;
assign v$Q_14147_out0 = v$G4_11834_out0;
assign v$Q_14158_out0 = v$G4_11839_out0;
assign v$A3XNORB3_14717_out0 = v$G8_3727_out0;
assign v$A3XNORB3_14718_out0 = v$G8_3728_out0;
assign v$A3XNORB3_14720_out0 = v$G8_3730_out0;
assign v$A3XNORB3_14721_out0 = v$G8_3731_out0;
assign v$A3XNORB3_14732_out0 = v$G8_3742_out0;
assign v$A3XNORB3_14733_out0 = v$G8_3743_out0;
assign v$A3XNORB3_14735_out0 = v$G8_3745_out0;
assign v$A3XNORB3_14736_out0 = v$G8_3746_out0;
assign v$G11_15638_out0 = v$A2_8058_out0 && v$G12_16469_out0;
assign v$G11_15639_out0 = v$A2_8059_out0 && v$G12_16470_out0;
assign v$G11_15641_out0 = v$A2_8061_out0 && v$G12_16472_out0;
assign v$G11_15642_out0 = v$A2_8062_out0 && v$G12_16473_out0;
assign v$G11_15653_out0 = v$A2_8073_out0 && v$G12_16484_out0;
assign v$G11_15654_out0 = v$A2_8074_out0 && v$G12_16485_out0;
assign v$G11_15656_out0 = v$A2_8076_out0 && v$G12_16487_out0;
assign v$G11_15657_out0 = v$A2_8077_out0 && v$G12_16488_out0;
assign v$A1XNORB1_16046_out0 = v$G16_16863_out0;
assign v$A1XNORB1_16047_out0 = v$G16_16864_out0;
assign v$A1XNORB1_16049_out0 = v$G16_16866_out0;
assign v$A1XNORB1_16050_out0 = v$G16_16867_out0;
assign v$A1XNORB1_16061_out0 = v$G16_16878_out0;
assign v$A1XNORB1_16062_out0 = v$G16_16879_out0;
assign v$A1XNORB1_16064_out0 = v$G16_16881_out0;
assign v$A1XNORB1_16065_out0 = v$G16_16882_out0;
assign v$SAME_18723_out0 = v$G41_10872_out0;
assign v$SAME_18727_out0 = v$G41_10875_out0;
assign v$SAME_18732_out0 = v$G1_9388_out0;
assign v$SAME_18743_out0 = v$G41_10887_out0;
assign v$SAME_18747_out0 = v$G41_10890_out0;
assign v$SAME_18752_out0 = v$G1_9393_out0;
assign v$MUX3_3393_out0 = v$OUT_3918_out0 ? v$A$EXP_286_out0 : v$B$EXP_16674_out0;
assign v$OUT_3914_out0 = v$G29_10298_out0;
assign v$OUT_3934_out0 = v$G29_10301_out0;
assign v$G13_4400_out0 = v$A3XNORB3_14717_out0 && v$G11_15638_out0;
assign v$G13_4401_out0 = v$A3XNORB3_14718_out0 && v$G11_15639_out0;
assign v$G13_4403_out0 = v$A3XNORB3_14720_out0 && v$G11_15641_out0;
assign v$G13_4404_out0 = v$A3XNORB3_14721_out0 && v$G11_15642_out0;
assign v$G13_4415_out0 = v$A3XNORB3_14732_out0 && v$G11_15653_out0;
assign v$G13_4416_out0 = v$A3XNORB3_14733_out0 && v$G11_15654_out0;
assign v$G13_4418_out0 = v$A3XNORB3_14735_out0 && v$G11_15656_out0;
assign v$G13_4419_out0 = v$A3XNORB3_14736_out0 && v$G11_15657_out0;
assign v$A3$COMP$B3_4946_out0 = v$G5_6935_out0;
assign v$A3$COMP$B3_4947_out0 = v$G5_6936_out0;
assign v$A3$COMP$B3_4949_out0 = v$G5_6938_out0;
assign v$A3$COMP$B3_4950_out0 = v$G5_6939_out0;
assign v$A3$COMP$B3_4961_out0 = v$G5_6950_out0;
assign v$A3$COMP$B3_4962_out0 = v$G5_6951_out0;
assign v$A3$COMP$B3_4964_out0 = v$G5_6953_out0;
assign v$A3$COMP$B3_4965_out0 = v$G5_6954_out0;
assign v$G3_8817_out0 = v$HIGHER$SAME_15023_out0 && v$LOWER$OUT_4224_out0;
assign v$G3_8818_out0 = v$HIGHER$SAME_15024_out0 && v$LOWER$OUT_4225_out0;
assign v$DIFF_9091_out0 = v$A1_5793_out0;
assign v$HIGHER$SAME_9132_out0 = v$SAME_18723_out0;
assign v$HIGHER$SAME_9133_out0 = v$SAME_18727_out0;
assign v$HIGHER$SAME_9134_out0 = v$SAME_18743_out0;
assign v$HIGHER$SAME_9135_out0 = v$SAME_18747_out0;
assign v$G41_10873_out0 = v$G38_7292_out0 && v$G40_13361_out0;
assign v$G41_10874_out0 = v$G38_7293_out0 && v$G40_13362_out0;
assign v$G41_10876_out0 = v$G38_7295_out0 && v$G40_13364_out0;
assign v$G41_10877_out0 = v$G38_7296_out0 && v$G40_13365_out0;
assign v$G41_10888_out0 = v$G38_7307_out0 && v$G40_13376_out0;
assign v$G41_10889_out0 = v$G38_7308_out0 && v$G40_13377_out0;
assign v$G41_10891_out0 = v$G38_7310_out0 && v$G40_13379_out0;
assign v$G41_10892_out0 = v$G38_7311_out0 && v$G40_13380_out0;
assign v$_11810_out0 = { v$_14635_out0,v$MUX6_2847_out0 };
assign v$_11814_out0 = { v$_14639_out0,v$MUX6_2848_out0 };
assign v$A1$COMP$B1_12486_out0 = v$G18_4973_out0;
assign v$A1$COMP$B1_12489_out0 = v$G18_4976_out0;
assign v$A1$COMP$B1_12501_out0 = v$G18_4988_out0;
assign v$A1$COMP$B1_12504_out0 = v$G18_4991_out0;
assign v$G28_13016_out0 = v$A1XNORB1_16046_out0 && v$G25_10935_out0;
assign v$G28_13017_out0 = v$A1XNORB1_16047_out0 && v$G25_10936_out0;
assign v$G28_13019_out0 = v$A1XNORB1_16049_out0 && v$G25_10938_out0;
assign v$G28_13020_out0 = v$A1XNORB1_16050_out0 && v$G25_10939_out0;
assign v$G28_13031_out0 = v$A1XNORB1_16061_out0 && v$G25_10950_out0;
assign v$G28_13032_out0 = v$A1XNORB1_16062_out0 && v$G25_10951_out0;
assign v$G28_13034_out0 = v$A1XNORB1_16064_out0 && v$G25_10953_out0;
assign v$G28_13035_out0 = v$A1XNORB1_16065_out0 && v$G25_10954_out0;
assign v$G22_13328_out0 = v$A2XNORB2_4491_out0 && v$G20_9883_out0;
assign v$G22_13329_out0 = v$A2XNORB2_4492_out0 && v$G20_9884_out0;
assign v$G22_13331_out0 = v$A2XNORB2_4494_out0 && v$G20_9886_out0;
assign v$G22_13332_out0 = v$A2XNORB2_4495_out0 && v$G20_9887_out0;
assign v$G22_13343_out0 = v$A2XNORB2_4506_out0 && v$G20_9898_out0;
assign v$G22_13344_out0 = v$A2XNORB2_4507_out0 && v$G20_9899_out0;
assign v$G22_13346_out0 = v$A2XNORB2_4509_out0 && v$G20_9901_out0;
assign v$G22_13347_out0 = v$A2XNORB2_4510_out0 && v$G20_9902_out0;
assign v$OUT_13758_out0 = v$OUT_3918_out0;
assign v$Q_14148_out0 = v$G4_11835_out0;
assign v$Q_14149_out0 = v$G4_11836_out0;
assign v$Q_14150_out0 = v$G4_11837_out0;
assign v$Q_14159_out0 = v$G4_11840_out0;
assign v$Q_14160_out0 = v$G4_11841_out0;
assign v$Q_14161_out0 = v$G4_11842_out0;
assign v$NOT$USED1_14382_out0 = v$A1_5793_out1;
assign v$TXFlag_15247_out0 = v$TXFlag_7718_out0;
assign v$TXFlag_15248_out0 = v$TXFlag_7719_out0;
assign v$G31_15513_out0 = v$A2$COMP$B2_1979_out0 || v$G32_399_out0;
assign v$G31_15514_out0 = v$A2$COMP$B2_1980_out0 || v$G32_400_out0;
assign v$G31_15528_out0 = v$A2$COMP$B2_1994_out0 || v$G32_414_out0;
assign v$G31_15529_out0 = v$A2$COMP$B2_1995_out0 || v$G32_415_out0;
assign v$G24_15684_out0 = v$A3XNORB3_14716_out0 && v$G27_4776_out0;
assign v$G24_15687_out0 = v$A3XNORB3_14719_out0 && v$G27_4779_out0;
assign v$G24_15699_out0 = v$A3XNORB3_14731_out0 && v$G27_4791_out0;
assign v$G24_15702_out0 = v$A3XNORB3_14734_out0 && v$G27_4794_out0;
assign v$RXflag_15841_out0 = v$Q_14147_out0;
assign v$RXflag_15842_out0 = v$Q_14158_out0;
assign v$G6_16809_out0 = ! v$IGNORE_8283_out0;
assign v$MUX1_17925_out0 = v$OUT_3918_out0 ? v$B$EXP_16674_out0 : v$A$EXP_286_out0;
assign v$SAME_18364_out0 = v$SAME_18732_out0;
assign v$SAME_18370_out0 = v$SAME_18752_out0;
assign v$G30_1776_out0 = v$A3$COMP$B3_4952_out0 || v$G31_15513_out0;
assign v$G30_1777_out0 = v$A3$COMP$B3_4953_out0 || v$G31_15514_out0;
assign v$G30_1791_out0 = v$A3$COMP$B3_4967_out0 || v$G31_15528_out0;
assign v$G30_1792_out0 = v$A3$COMP$B3_4968_out0 || v$G31_15529_out0;
assign v$A2$COMP$B2_1973_out0 = v$G13_4400_out0;
assign v$A2$COMP$B2_1974_out0 = v$G13_4401_out0;
assign v$A2$COMP$B2_1976_out0 = v$G13_4403_out0;
assign v$A2$COMP$B2_1977_out0 = v$G13_4404_out0;
assign v$A2$COMP$B2_1988_out0 = v$G13_4415_out0;
assign v$A2$COMP$B2_1989_out0 = v$G13_4416_out0;
assign v$A2$COMP$B2_1991_out0 = v$G13_4418_out0;
assign v$A2$COMP$B2_1992_out0 = v$G13_4419_out0;
assign v$MUX14_2957_out0 = v$IS$32$BIT_10862_out0 ? v$SAME_18364_out0 : v$SAME_18363_out0;
assign v$MUX14_2958_out0 = v$IS$32$BIT_10863_out0 ? v$SAME_18370_out0 : v$SAME_18369_out0;
assign v$MUX3_3391_out0 = v$OUT_3914_out0 ? v$A$EXP_284_out0 : v$B$EXP_16672_out0;
assign v$MUX3_3397_out0 = v$OUT_3934_out0 ? v$A$EXP_290_out0 : v$B$EXP_16678_out0;
assign v$Error_3767_out0 = v$Q_14150_out0;
assign v$Error_3768_out0 = v$Q_14161_out0;
assign v$TXoverflow_4108_out0 = v$Q_14148_out0;
assign v$TXoverflow_4109_out0 = v$Q_14159_out0;
assign v$G27_4777_out0 = v$A2XNORB2_4491_out0 && v$G28_13016_out0;
assign v$G27_4778_out0 = v$A2XNORB2_4492_out0 && v$G28_13017_out0;
assign v$G27_4780_out0 = v$A2XNORB2_4494_out0 && v$G28_13019_out0;
assign v$G27_4781_out0 = v$A2XNORB2_4495_out0 && v$G28_13020_out0;
assign v$G27_4792_out0 = v$A2XNORB2_4506_out0 && v$G28_13031_out0;
assign v$G27_4793_out0 = v$A2XNORB2_4507_out0 && v$G28_13032_out0;
assign v$G27_4795_out0 = v$A2XNORB2_4509_out0 && v$G28_13034_out0;
assign v$G27_4796_out0 = v$A2XNORB2_4510_out0 && v$G28_13035_out0;
assign v$G18_4974_out0 = v$A3XNORB3_14717_out0 && v$G22_13328_out0;
assign v$G18_4975_out0 = v$A3XNORB3_14718_out0 && v$G22_13329_out0;
assign v$G18_4977_out0 = v$A3XNORB3_14720_out0 && v$G22_13331_out0;
assign v$G18_4978_out0 = v$A3XNORB3_14721_out0 && v$G22_13332_out0;
assign v$G18_4989_out0 = v$A3XNORB3_14732_out0 && v$G22_13343_out0;
assign v$G18_4990_out0 = v$A3XNORB3_14733_out0 && v$G22_13344_out0;
assign v$G18_4992_out0 = v$A3XNORB3_14735_out0 && v$G22_13346_out0;
assign v$G18_4993_out0 = v$A3XNORB3_14736_out0 && v$G22_13347_out0;
assign v$MUX1_6679_out0 = v$G4_4031_out0 ? v$_11810_out0 : v$MUX2_12040_out0;
assign v$MUX1_6683_out0 = v$G4_4035_out0 ? v$_11814_out0 : v$MUX2_12044_out0;
assign v$XOR1_7591_out0 = v$C1_13576_out0 ^ v$MUX1_17925_out0;
assign v$A0$COMP$B0_7986_out0 = v$G24_15684_out0;
assign v$A0$COMP$B0_7989_out0 = v$G24_15687_out0;
assign v$A0$COMP$B0_8001_out0 = v$G24_15699_out0;
assign v$A0$COMP$B0_8004_out0 = v$G24_15702_out0;
assign v$RXoverflow_9540_out0 = v$Q_14149_out0;
assign v$RXoverflow_9541_out0 = v$Q_14160_out0;
assign v$RXFLAG_12134_out0 = v$RXflag_15841_out0;
assign v$RXFLAG_12135_out0 = v$RXflag_15842_out0;
assign v$G2_12907_out0 = v$HIGHER$OUT_3832_out0 || v$G3_8817_out0;
assign v$G2_12908_out0 = v$HIGHER$OUT_3833_out0 || v$G3_8818_out0;
assign v$OUT_13756_out0 = v$OUT_3914_out0;
assign v$OUT_13762_out0 = v$OUT_3934_out0;
assign v$TXFLAG_14691_out0 = v$TXFlag_15247_out0;
assign v$TXFLAG_14692_out0 = v$TXFlag_15248_out0;
assign v$_17406_out0 = { v$DIFF_9091_out0,v$C2_13326_out0 };
assign v$G7_17665_out0 = v$G5_2668_out0 && v$G6_16809_out0;
assign v$MUX1_17923_out0 = v$OUT_3914_out0 ? v$B$EXP_16672_out0 : v$A$EXP_284_out0;
assign v$MUX1_17929_out0 = v$OUT_3934_out0 ? v$B$EXP_16678_out0 : v$A$EXP_290_out0;
assign v$SAME_18725_out0 = v$G41_10873_out0;
assign v$SAME_18726_out0 = v$G41_10874_out0;
assign v$SAME_18729_out0 = v$G41_10876_out0;
assign v$SAME_18730_out0 = v$G41_10877_out0;
assign v$SAME_18745_out0 = v$G41_10888_out0;
assign v$SAME_18746_out0 = v$G41_10889_out0;
assign v$SAME_18749_out0 = v$G41_10891_out0;
assign v$SAME_18750_out0 = v$G41_10892_out0;
assign v$G32_392_out0 = v$A1$COMP$B1_12486_out0 || v$A0$COMP$B0_7986_out0;
assign v$G32_395_out0 = v$A1$COMP$B1_12489_out0 || v$A0$COMP$B0_7989_out0;
assign v$G32_407_out0 = v$A1$COMP$B1_12501_out0 || v$A0$COMP$B0_8001_out0;
assign v$G32_410_out0 = v$A1$COMP$B1_12504_out0 || v$A0$COMP$B0_8004_out0;
assign v$EXP$SAME_903_out0 = v$MUX14_2957_out0;
assign v$EXP$SAME_904_out0 = v$MUX14_2958_out0;
assign v$MUX3_1959_out0 = v$G8_1888_out0 ? v$_13306_out0 : v$MUX1_6679_out0;
assign v$MUX3_1963_out0 = v$G8_1892_out0 ? v$_13310_out0 : v$MUX1_6683_out0;
assign v$TXFLAG_3878_out0 = v$TXFLAG_14691_out0;
assign v$TXFLAG_3879_out0 = v$TXFLAG_14692_out0;
assign v$OUT_3916_out0 = v$G30_1776_out0;
assign v$OUT_3917_out0 = v$G30_1777_out0;
assign v$OUT_3919_out0 = v$G2_12907_out0;
assign v$OUT_3923_out0 = v$G2_12908_out0;
assign v$OUT_3936_out0 = v$G30_1791_out0;
assign v$OUT_3937_out0 = v$G30_1792_out0;
assign {v$A1_5791_out1,v$A1_5791_out0 } = v$MUX3_3393_out0 + v$XOR1_7591_out0 + v$CIN_18227_out0;
assign v$XOR1_7589_out0 = v$C1_13574_out0 ^ v$MUX1_17923_out0;
assign v$XOR1_7595_out0 = v$C1_13580_out0 ^ v$MUX1_17929_out0;
assign v$_9917_out0 = { v$RXoverflow_9540_out0,v$Error_3767_out0 };
assign v$_9918_out0 = { v$RXoverflow_9541_out0,v$Error_3768_out0 };
assign v$LOWER$SAME_10181_out0 = v$SAME_18726_out0;
assign v$LOWER$SAME_10182_out0 = v$SAME_18730_out0;
assign v$LOWER$SAME_10186_out0 = v$SAME_18746_out0;
assign v$LOWER$SAME_10187_out0 = v$SAME_18750_out0;
assign v$A1$COMP$B1_12487_out0 = v$G18_4974_out0;
assign v$A1$COMP$B1_12488_out0 = v$G18_4975_out0;
assign v$A1$COMP$B1_12490_out0 = v$G18_4977_out0;
assign v$A1$COMP$B1_12491_out0 = v$G18_4978_out0;
assign v$A1$COMP$B1_12502_out0 = v$G18_4989_out0;
assign v$A1$COMP$B1_12503_out0 = v$G18_4990_out0;
assign v$A1$COMP$B1_12505_out0 = v$G18_4992_out0;
assign v$A1$COMP$B1_12506_out0 = v$G18_4993_out0;
assign v$RXFLAG_15003_out0 = v$RXFLAG_12134_out0;
assign v$RXFLAG_15004_out0 = v$RXFLAG_12135_out0;
assign v$HIGHER$SAME_15020_out0 = v$SAME_18725_out0;
assign v$HIGHER$SAME_15021_out0 = v$SAME_18729_out0;
assign v$HIGHER$SAME_15025_out0 = v$SAME_18745_out0;
assign v$HIGHER$SAME_15026_out0 = v$SAME_18749_out0;
assign v$_15298_out0 = { v$TXFlag_7718_out0,v$TXoverflow_4108_out0 };
assign v$_15299_out0 = { v$TXFlag_7719_out0,v$TXoverflow_4109_out0 };
assign v$G24_15685_out0 = v$A3XNORB3_14717_out0 && v$G27_4777_out0;
assign v$G24_15686_out0 = v$A3XNORB3_14718_out0 && v$G27_4778_out0;
assign v$G24_15688_out0 = v$A3XNORB3_14720_out0 && v$G27_4780_out0;
assign v$G24_15689_out0 = v$A3XNORB3_14721_out0 && v$G27_4781_out0;
assign v$G24_15700_out0 = v$A3XNORB3_14732_out0 && v$G27_4792_out0;
assign v$G24_15701_out0 = v$A3XNORB3_14733_out0 && v$G27_4793_out0;
assign v$G24_15703_out0 = v$A3XNORB3_14735_out0 && v$G27_4795_out0;
assign v$G24_15704_out0 = v$A3XNORB3_14736_out0 && v$G27_4796_out0;
assign v$RAMWEN_17961_out0 = v$G7_17665_out0;
assign v$F_1969_out0 = v$TXFLAG_3878_out0;
assign v$F_1970_out0 = v$TXFLAG_3879_out0;
assign v$OUT_3178_out0 = v$MUX3_1959_out0;
assign v$OUT_3182_out0 = v$MUX3_1963_out0;
assign v$MUX3_3394_out0 = v$OUT_3919_out0 ? v$A$EXP_287_out0 : v$B$EXP_16675_out0;
assign v$MUX3_3396_out0 = v$OUT_3923_out0 ? v$A$EXP_289_out0 : v$B$EXP_16677_out0;
assign v$HIGHER$OUT_3831_out0 = v$OUT_3916_out0;
assign v$HIGHER$OUT_3836_out0 = v$OUT_3936_out0;
assign v$LOWER$OUT_4223_out0 = v$OUT_3917_out0;
assign v$LOWER$OUT_4228_out0 = v$OUT_3937_out0;
assign {v$A1_5789_out1,v$A1_5789_out0 } = v$MUX3_3391_out0 + v$XOR1_7589_out0 + v$CIN_18225_out0;
assign {v$A1_5795_out1,v$A1_5795_out0 } = v$MUX3_3397_out0 + v$XOR1_7595_out0 + v$CIN_18231_out0;
assign v$A0$COMP$B0_7987_out0 = v$G24_15685_out0;
assign v$A0$COMP$B0_7988_out0 = v$G24_15686_out0;
assign v$A0$COMP$B0_7990_out0 = v$G24_15688_out0;
assign v$A0$COMP$B0_7991_out0 = v$G24_15689_out0;
assign v$A0$COMP$B0_8002_out0 = v$G24_15700_out0;
assign v$A0$COMP$B0_8003_out0 = v$G24_15701_out0;
assign v$A0$COMP$B0_8005_out0 = v$G24_15703_out0;
assign v$A0$COMP$B0_8006_out0 = v$G24_15704_out0;
assign v$DIFF_9089_out0 = v$A1_5791_out0;
assign v$G1_9386_out0 = v$LOWER$SAME_10181_out0 && v$HIGHER$SAME_15020_out0;
assign v$G1_9387_out0 = v$LOWER$SAME_10182_out0 && v$HIGHER$SAME_15021_out0;
assign v$G1_9391_out0 = v$LOWER$SAME_10186_out0 && v$HIGHER$SAME_15025_out0;
assign v$G1_9392_out0 = v$LOWER$SAME_10187_out0 && v$HIGHER$SAME_15026_out0;
assign v$OUT_13759_out0 = v$OUT_3919_out0;
assign v$OUT_13761_out0 = v$OUT_3923_out0;
assign v$NOT$USED1_14380_out0 = v$A1_5791_out1;
assign v$G31_15506_out0 = v$A2$COMP$B2_1972_out0 || v$G32_392_out0;
assign v$G31_15509_out0 = v$A2$COMP$B2_1975_out0 || v$G32_395_out0;
assign v$G31_15521_out0 = v$A2$COMP$B2_1987_out0 || v$G32_407_out0;
assign v$G31_15524_out0 = v$A2$COMP$B2_1990_out0 || v$G32_410_out0;
assign v$MUX1_17926_out0 = v$OUT_3919_out0 ? v$B$EXP_16675_out0 : v$A$EXP_287_out0;
assign v$MUX1_17928_out0 = v$OUT_3923_out0 ? v$B$EXP_16677_out0 : v$A$EXP_289_out0;
assign v$_18544_out0 = { v$RXflag_15841_out0,v$_9917_out0 };
assign v$_18545_out0 = { v$RXflag_15842_out0,v$_9918_out0 };
assign v$G32_393_out0 = v$A1$COMP$B1_12487_out0 || v$A0$COMP$B0_7987_out0;
assign v$G32_394_out0 = v$A1$COMP$B1_12488_out0 || v$A0$COMP$B0_7988_out0;
assign v$G32_396_out0 = v$A1$COMP$B1_12490_out0 || v$A0$COMP$B0_7990_out0;
assign v$G32_397_out0 = v$A1$COMP$B1_12491_out0 || v$A0$COMP$B0_7991_out0;
assign v$G32_408_out0 = v$A1$COMP$B1_12502_out0 || v$A0$COMP$B0_8002_out0;
assign v$G32_409_out0 = v$A1$COMP$B1_12503_out0 || v$A0$COMP$B0_8003_out0;
assign v$G32_411_out0 = v$A1$COMP$B1_12505_out0 || v$A0$COMP$B0_8005_out0;
assign v$G32_412_out0 = v$A1$COMP$B1_12506_out0 || v$A0$COMP$B0_8006_out0;
assign v$G30_1769_out0 = v$A3$COMP$B3_4945_out0 || v$G31_15506_out0;
assign v$G30_1772_out0 = v$A3$COMP$B3_4948_out0 || v$G31_15509_out0;
assign v$G30_1784_out0 = v$A3$COMP$B3_4960_out0 || v$G31_15521_out0;
assign v$G30_1787_out0 = v$A3$COMP$B3_4963_out0 || v$G31_15524_out0;
assign v$G51_3464_out0 = v$NQ1_11038_out0 && v$F_1969_out0;
assign v$G51_3465_out0 = v$NQ1_11039_out0 && v$F_1970_out0;
assign v$G28_3765_out0 = ! v$F_1969_out0;
assign v$G28_3766_out0 = ! v$F_1970_out0;
assign v$IN_4363_out0 = v$OUT_3178_out0;
assign v$IN_4367_out0 = v$OUT_3182_out0;
assign v$_6341_out0 = { v$_15298_out0,v$_18544_out0 };
assign v$_6342_out0 = { v$_15299_out0,v$_18545_out0 };
assign v$XOR1_7592_out0 = v$C1_13577_out0 ^ v$MUX1_17926_out0;
assign v$XOR1_7594_out0 = v$C1_13579_out0 ^ v$MUX1_17928_out0;
assign v$G3_8816_out0 = v$HIGHER$SAME_15022_out0 && v$LOWER$OUT_4223_out0;
assign v$G3_8821_out0 = v$HIGHER$SAME_15027_out0 && v$LOWER$OUT_4228_out0;
assign v$DIFF_9087_out0 = v$A1_5789_out0;
assign v$DIFF_9093_out0 = v$A1_5795_out0;
assign v$NOT$USED1_14378_out0 = v$A1_5789_out1;
assign v$NOT$USED1_14384_out0 = v$A1_5795_out1;
assign v$MUX5_15500_out0 = v$IS$32$BITS_2992_out0 ? v$OUT_13759_out0 : v$OUT_13758_out0;
assign v$MUX5_15501_out0 = v$IS$32$BITS_1282_out0 ? v$OUT_13761_out0 : v$OUT_13760_out0;
assign v$_17405_out0 = { v$DIFF_9089_out0,v$C2_13325_out0 };
assign v$SAME_18724_out0 = v$G1_9386_out0;
assign v$SAME_18728_out0 = v$G1_9387_out0;
assign v$SAME_18744_out0 = v$G1_9391_out0;
assign v$SAME_18748_out0 = v$G1_9392_out0;
assign v$LOWER$SAME_3793_out0 = v$SAME_18724_out0;
assign v$LOWER$SAME_3794_out0 = v$SAME_18728_out0;
assign v$LOWER$SAME_3795_out0 = v$SAME_18744_out0;
assign v$LOWER$SAME_3796_out0 = v$SAME_18748_out0;
assign v$OUT_3906_out0 = v$G30_1769_out0;
assign v$OUT_3910_out0 = v$G30_1772_out0;
assign v$OUT_3926_out0 = v$G30_1784_out0;
assign v$OUT_3930_out0 = v$G30_1787_out0;
assign {v$A1_5792_out1,v$A1_5792_out0 } = v$MUX3_3394_out0 + v$XOR1_7592_out0 + v$CIN_18228_out0;
assign {v$A1_5794_out1,v$A1_5794_out0 } = v$MUX3_3396_out0 + v$XOR1_7594_out0 + v$CIN_18230_out0;
assign v$_7610_out0 = { v$DIFF_9087_out0,v$C4_6625_out0 };
assign v$_7611_out0 = { v$DIFF_9093_out0,v$C4_6626_out0 };
assign v$A$EXP$LARGER_9441_out0 = v$MUX5_15500_out0;
assign v$A$EXP$LARGER_9442_out0 = v$MUX5_15501_out0;
assign v$IN_9569_out0 = v$IN_4363_out0;
assign v$IN_9573_out0 = v$IN_4367_out0;
assign v$G49_11052_out0 = v$G50_17323_out0 || v$G51_3464_out0;
assign v$G49_11053_out0 = v$G50_17324_out0 || v$G51_3465_out0;
assign v$G2_12906_out0 = v$HIGHER$OUT_3831_out0 || v$G3_8816_out0;
assign v$G2_12911_out0 = v$HIGHER$OUT_3836_out0 || v$G3_8821_out0;
assign v$NF_14564_out0 = v$G28_3765_out0;
assign v$NF_14565_out0 = v$G28_3766_out0;
assign v$G31_15507_out0 = v$A2$COMP$B2_1973_out0 || v$G32_393_out0;
assign v$G31_15508_out0 = v$A2$COMP$B2_1974_out0 || v$G32_394_out0;
assign v$G31_15510_out0 = v$A2$COMP$B2_1976_out0 || v$G32_396_out0;
assign v$G31_15511_out0 = v$A2$COMP$B2_1977_out0 || v$G32_397_out0;
assign v$G31_15522_out0 = v$A2$COMP$B2_1988_out0 || v$G32_408_out0;
assign v$G31_15523_out0 = v$A2$COMP$B2_1989_out0 || v$G32_409_out0;
assign v$G31_15525_out0 = v$A2$COMP$B2_1991_out0 || v$G32_411_out0;
assign v$G31_15526_out0 = v$A2$COMP$B2_1992_out0 || v$G32_412_out0;
assign v$_16169_out0 = { v$_6341_out0,v$C1_16842_out0 };
assign v$_16170_out0 = { v$_6342_out0,v$C1_16843_out0 };
assign v$G30_1770_out0 = v$A3$COMP$B3_4946_out0 || v$G31_15507_out0;
assign v$G30_1771_out0 = v$A3$COMP$B3_4947_out0 || v$G31_15508_out0;
assign v$G30_1773_out0 = v$A3$COMP$B3_4949_out0 || v$G31_15510_out0;
assign v$G30_1774_out0 = v$A3$COMP$B3_4950_out0 || v$G31_15511_out0;
assign v$G30_1785_out0 = v$A3$COMP$B3_4961_out0 || v$G31_15522_out0;
assign v$G30_1786_out0 = v$A3$COMP$B3_4962_out0 || v$G31_15523_out0;
assign v$G30_1788_out0 = v$A3$COMP$B3_4964_out0 || v$G31_15525_out0;
assign v$G30_1789_out0 = v$A3$COMP$B3_4965_out0 || v$G31_15526_out0;
assign v$G2_1894_out0 = v$EXP$SAME_16546_out0 || v$A$EXP$LARGER_9441_out0;
assign v$G2_1895_out0 = v$EXP$SAME_16547_out0 || v$A$EXP$LARGER_9442_out0;
assign v$Status_3791_out0 = v$_16169_out0;
assign v$Status_3792_out0 = v$_16170_out0;
assign v$OUT_3915_out0 = v$G2_12906_out0;
assign v$OUT_3935_out0 = v$G2_12911_out0;
assign v$_4803_out0 = v$IN_9569_out0[7:0];
assign v$_4807_out0 = v$IN_9573_out0[7:0];
assign v$_7476_out0 = v$IN_9569_out0[15:15];
assign v$_7477_out0 = v$IN_9573_out0[15:15];
assign v$HIGHER$OUT_7785_out0 = v$OUT_3906_out0;
assign v$HIGHER$OUT_7786_out0 = v$OUT_3910_out0;
assign v$HIGHER$OUT_7787_out0 = v$OUT_3926_out0;
assign v$HIGHER$OUT_7788_out0 = v$OUT_3930_out0;
assign v$DIFF_9090_out0 = v$A1_5792_out0;
assign v$DIFF_9092_out0 = v$A1_5794_out0;
assign v$_13271_out0 = v$IN_9569_out0[7:0];
assign v$_13274_out0 = v$IN_9573_out0[7:0];
assign v$_14093_out0 = v$IN_9569_out0[7:0];
assign v$_14094_out0 = v$IN_9573_out0[7:0];
assign v$NOT$USED1_14381_out0 = v$A1_5792_out1;
assign v$NOT$USED1_14383_out0 = v$A1_5794_out1;
assign v$_14602_out0 = v$IN_9569_out0[15:8];
assign v$_14606_out0 = v$IN_9573_out0[15:8];
assign v$_14636_out0 = v$IN_9569_out0[15:8];
assign v$_14640_out0 = v$IN_9573_out0[15:8];
assign v$IS$A$LARGER_14661_out0 = v$A$EXP$LARGER_9441_out0;
assign v$IS$A$LARGER_14662_out0 = v$A$EXP$LARGER_9442_out0;
assign v$G4_15340_out0 = v$EXP$SAME_16546_out0 || v$A$EXP$LARGER_9441_out0;
assign v$G4_15341_out0 = v$EXP$SAME_16547_out0 || v$A$EXP$LARGER_9442_out0;
assign v$_16750_out0 = v$IN_9569_out0[15:8];
assign v$_16754_out0 = v$IN_9573_out0[15:8];
assign v$G1_17446_out0 = v$LOWER$SAME_3793_out0 && v$HIGHER$SAME_9132_out0;
assign v$G1_17447_out0 = v$LOWER$SAME_3794_out0 && v$HIGHER$SAME_9133_out0;
assign v$G1_17448_out0 = v$LOWER$SAME_3795_out0 && v$HIGHER$SAME_9134_out0;
assign v$G1_17449_out0 = v$LOWER$SAME_3796_out0 && v$HIGHER$SAME_9135_out0;
assign v$G48_18516_out0 = v$NQ0_15621_out0 && v$G49_11052_out0;
assign v$G48_18517_out0 = v$NQ0_15622_out0 && v$G49_11053_out0;
assign v$_1480_out0 = { v$C1_7974_out0,v$_4803_out0 };
assign v$_1484_out0 = { v$C1_7978_out0,v$_4807_out0 };
assign v$MUX2_1609_out0 = v$IS$A$LARGER_14661_out0 ? v$SEL4_2279_out0 : v$SEL3_11894_out0;
assign v$MUX2_1610_out0 = v$IS$A$LARGER_14662_out0 ? v$SEL4_2280_out0 : v$SEL3_11895_out0;
assign v$MUX1_1933_out0 = v$IS$A$LARGER_14661_out0 ? v$SEL1_15748_out0 : v$SEL2_11011_out0;
assign v$MUX1_1934_out0 = v$IS$A$LARGER_14662_out0 ? v$SEL1_15749_out0 : v$SEL2_11012_out0;
assign v$MUX3_3392_out0 = v$OUT_3915_out0 ? v$A$EXP_285_out0 : v$B$EXP_16673_out0;
assign v$MUX3_3398_out0 = v$OUT_3935_out0 ? v$A$EXP_291_out0 : v$B$EXP_16679_out0;
assign v$OUT_3908_out0 = v$G30_1770_out0;
assign v$OUT_3909_out0 = v$G30_1771_out0;
assign v$OUT_3912_out0 = v$G30_1773_out0;
assign v$OUT_3913_out0 = v$G30_1774_out0;
assign v$OUT_3928_out0 = v$G30_1785_out0;
assign v$OUT_3929_out0 = v$G30_1786_out0;
assign v$OUT_3932_out0 = v$G30_1788_out0;
assign v$OUT_3933_out0 = v$G30_1789_out0;
assign v$MUX1_4041_out0 = v$G2_1894_out0 ? v$B_6548_out0 : v$A_2293_out0;
assign v$MUX1_4042_out0 = v$G2_1895_out0 ? v$B_12138_out0 : v$A_16090_out0;
assign v$MUX6_7948_out0 = v$IS$32$BITS_2992_out0 ? v$DIFF_9090_out0 : v$_17405_out0;
assign v$MUX6_7949_out0 = v$IS$32$BITS_1282_out0 ? v$DIFF_9092_out0 : v$_17406_out0;
assign v$STATUS_8810_out0 = v$Status_3791_out0;
assign v$STATUS_8811_out0 = v$Status_3792_out0;
assign v$SAME_8919_out0 = v$G1_17446_out0;
assign v$SAME_8920_out0 = v$G1_17447_out0;
assign v$SAME_8921_out0 = v$G1_17448_out0;
assign v$SAME_8922_out0 = v$G1_17449_out0;
assign v$_9448_out0 = { v$_16750_out0,v$LSBS_7937_out0 };
assign v$_9452_out0 = { v$_16754_out0,v$LSBS_7938_out0 };
assign v$_13307_out0 = { v$_14602_out0,v$_13271_out0 };
assign v$_13311_out0 = { v$_14606_out0,v$_13274_out0 };
assign v$MUX6_13706_out0 = v$S_17947_out0 ? v$_14093_out0 : v$C1_13448_out0;
assign v$MUX6_13707_out0 = v$S_17948_out0 ? v$_14094_out0 : v$C1_13449_out0;
assign v$OUT_13757_out0 = v$OUT_3915_out0;
assign v$OUT_13763_out0 = v$OUT_3935_out0;
assign v$MUX2_15190_out0 = v$G2_1894_out0 ? v$A_2293_out0 : v$B_6548_out0;
assign v$MUX2_15191_out0 = v$G2_1895_out0 ? v$A_16090_out0 : v$B_12138_out0;
assign v$MUX10_16829_out0 = v$G4_15340_out0 ? v$A_2293_out0 : v$B_6548_out0;
assign v$MUX10_16830_out0 = v$G4_15341_out0 ? v$A_16090_out0 : v$B_12138_out0;
assign v$G5_17879_out0 = v$G6_3163_out0 || v$G48_18516_out0;
assign v$G5_17880_out0 = v$G6_3164_out0 || v$G48_18517_out0;
assign v$MUX1_17924_out0 = v$OUT_3915_out0 ? v$B$EXP_16673_out0 : v$A$EXP_285_out0;
assign v$MUX1_17930_out0 = v$OUT_3935_out0 ? v$B$EXP_16679_out0 : v$A$EXP_291_out0;
assign v$MUX9_17941_out0 = v$G4_15340_out0 ? v$B_6548_out0 : v$A_2293_out0;
assign v$MUX9_17942_out0 = v$G4_15341_out0 ? v$B_12138_out0 : v$A_16090_out0;
assign v$_17969_out0 = { v$_7476_out0,v$_7476_out0 };
assign v$_17970_out0 = { v$_7477_out0,v$_7477_out0 };
assign v$SEL10_3010_out0 = v$MUX9_17941_out0[14:10];
assign v$SEL10_3011_out0 = v$MUX9_17942_out0[14:10];
assign v$SEL9_3773_out0 = v$MUX10_16829_out0[14:10];
assign v$SEL9_3774_out0 = v$MUX10_16830_out0[14:10];
assign v$HIGHER$OUT_3829_out0 = v$OUT_3908_out0;
assign v$HIGHER$OUT_3830_out0 = v$OUT_3912_out0;
assign v$HIGHER$OUT_3834_out0 = v$OUT_3928_out0;
assign v$HIGHER$OUT_3835_out0 = v$OUT_3932_out0;
assign v$LOWER$OUT_4221_out0 = v$OUT_3909_out0;
assign v$LOWER$OUT_4222_out0 = v$OUT_3913_out0;
assign v$LOWER$OUT_4226_out0 = v$OUT_3929_out0;
assign v$LOWER$OUT_4227_out0 = v$OUT_3933_out0;
assign v$MUX2_4852_out0 = v$IS$32$BIT_10862_out0 ? v$OUT_13757_out0 : v$OUT_13756_out0;
assign v$MUX2_4853_out0 = v$IS$32$BIT_10863_out0 ? v$OUT_13763_out0 : v$OUT_13762_out0;
assign v$XOR1_7590_out0 = v$C1_13575_out0 ^ v$MUX1_17924_out0;
assign v$XOR1_7596_out0 = v$C1_13581_out0 ^ v$MUX1_17930_out0;
assign v$MUX1_7642_out0 = v$G47_1531_out0 ? v$C1_1471_out0 : v$G5_17879_out0;
assign v$MUX1_7643_out0 = v$G47_1532_out0 ? v$C1_1472_out0 : v$G5_17880_out0;
assign v$SAME$H_8915_out0 = v$SAME_8919_out0;
assign v$SAME$H_8916_out0 = v$SAME_8921_out0;
assign v$_11015_out0 = { v$MUX2_1609_out0,v$C2_3628_out0 };
assign v$_11016_out0 = { v$MUX2_1610_out0,v$C2_3629_out0 };
assign v$SEL4_12199_out0 = v$MUX2_15190_out0[14:7];
assign v$SEL4_12200_out0 = v$MUX2_15191_out0[14:7];
assign v$EXP$DIFF_12470_out0 = v$MUX6_7948_out0;
assign v$EXP$DIFF_12471_out0 = v$MUX6_7949_out0;
assign v$_14091_out0 = { v$MUX1_1933_out0,v$C1_4356_out0 };
assign v$_14092_out0 = { v$MUX1_1934_out0,v$C1_4357_out0 };
assign v$MUX4_15993_out0 = v$EN_16968_out0 ? v$_1480_out0 : v$IN_9569_out0;
assign v$MUX4_15997_out0 = v$EN_16972_out0 ? v$_1484_out0 : v$IN_9573_out0;
assign v$SAME$L_16440_out0 = v$SAME_8920_out0;
assign v$SAME$L_16441_out0 = v$SAME_8922_out0;
assign v$_17409_out0 = { v$_17969_out0,v$_17969_out0 };
assign v$_17410_out0 = { v$_17970_out0,v$_17970_out0 };
assign v$MUX2_17760_out0 = v$FF2_9418_out0 ? v$STATUS_8810_out0 : v$RXBYTE_9628_out0;
assign v$MUX2_17761_out0 = v$FF2_9419_out0 ? v$STATUS_8811_out0 : v$RXBYTE_9629_out0;
assign v$SEL3_17817_out0 = v$MUX1_4041_out0[14:7];
assign v$SEL3_17818_out0 = v$MUX1_4042_out0[14:7];
assign v$SMALLER$EXP_2941_out0 = v$SEL10_3010_out0;
assign v$SMALLER$EXP_2942_out0 = v$SEL3_17817_out0;
assign v$SMALLER$EXP_2943_out0 = v$SEL10_3011_out0;
assign v$SMALLER$EXP_2944_out0 = v$SEL3_17818_out0;
assign {v$A1_5790_out1,v$A1_5790_out0 } = v$MUX3_3392_out0 + v$XOR1_7590_out0 + v$CIN_18226_out0;
assign {v$A1_5796_out1,v$A1_5796_out0 } = v$MUX3_3398_out0 + v$XOR1_7596_out0 + v$CIN_18232_out0;
assign v$_6913_out0 = { v$MUX2_17760_out0,v$C1_14812_out0 };
assign v$_6914_out0 = { v$MUX2_17761_out0,v$C1_14813_out0 };
assign v$G3_8814_out0 = v$HIGHER$SAME_15020_out0 && v$LOWER$OUT_4221_out0;
assign v$G3_8815_out0 = v$HIGHER$SAME_15021_out0 && v$LOWER$OUT_4222_out0;
assign v$G3_8819_out0 = v$HIGHER$SAME_15025_out0 && v$LOWER$OUT_4226_out0;
assign v$G3_8820_out0 = v$HIGHER$SAME_15026_out0 && v$LOWER$OUT_4227_out0;
assign v$LARGER$EXP_10274_out0 = v$SEL9_3773_out0;
assign v$LARGER$EXP_10275_out0 = v$SEL4_12199_out0;
assign v$LARGER$EXP_10276_out0 = v$SEL9_3774_out0;
assign v$LARGER$EXP_10277_out0 = v$SEL4_12200_out0;
assign v$MUX2_12041_out0 = v$G3_2608_out0 ? v$_9448_out0 : v$MUX4_15993_out0;
assign v$MUX2_12045_out0 = v$G3_2612_out0 ? v$_9452_out0 : v$MUX4_15997_out0;
assign v$IN_13168_out0 = v$_11015_out0;
assign v$IN_13169_out0 = v$_11016_out0;
assign v$_14313_out0 = { v$_17409_out0,v$_17409_out0 };
assign v$_14314_out0 = { v$_17410_out0,v$_17410_out0 };
assign v$EXP$DIFF_14330_out0 = v$EXP$DIFF_12470_out0;
assign v$EXP$DIFF_14331_out0 = v$EXP$DIFF_12471_out0;
assign v$SEL5_16175_out0 = v$_14091_out0[23:13];
assign v$SEL5_16176_out0 = v$_14092_out0[23:13];
assign v$Q0P_16773_out0 = v$MUX1_7642_out0;
assign v$Q0P_16774_out0 = v$MUX1_7643_out0;
assign v$DIFF_17503_out0 = v$EXP$DIFF_12470_out0;
assign v$DIFF_17504_out0 = v$EXP$DIFF_12470_out0;
assign v$DIFF_17505_out0 = v$EXP$DIFF_12471_out0;
assign v$DIFF_17506_out0 = v$EXP$DIFF_12471_out0;
assign v$A$EXP$LARGER_18245_out0 = v$MUX2_4852_out0;
assign v$A$EXP$LARGER_18246_out0 = v$MUX2_4853_out0;
assign v$G4_18277_out0 = v$SAME$L_16440_out0 && v$SAME$H_8915_out0;
assign v$G4_18278_out0 = v$SAME$L_16441_out0 && v$SAME$H_8916_out0;
assign v$MUX1_1996_out0 = v$FF1_11054_out0 ? v$_6913_out0 : v$RAMDOUT_16779_out0;
assign v$MUX1_1997_out0 = v$FF1_11055_out0 ? v$_6914_out0 : v$RAMDOUT_16780_out0;
assign v$IN_5169_out0 = v$IN_13168_out0;
assign v$IN_5180_out0 = v$IN_13169_out0;
assign v$SAME_6264_out0 = v$G4_18277_out0;
assign v$SAME_6265_out0 = v$G4_18278_out0;
assign v$DIFF_9088_out0 = v$A1_5790_out0;
assign v$DIFF_9094_out0 = v$A1_5796_out0;
assign v$_10038_out0 = { v$C4_2451_out0,v$SEL5_16175_out0 };
assign v$_10039_out0 = { v$C4_2452_out0,v$SEL5_16176_out0 };
assign v$G2_12904_out0 = v$HIGHER$OUT_3829_out0 || v$G3_8814_out0;
assign v$G2_12905_out0 = v$HIGHER$OUT_3830_out0 || v$G3_8815_out0;
assign v$G2_12909_out0 = v$HIGHER$OUT_3834_out0 || v$G3_8819_out0;
assign v$G2_12910_out0 = v$HIGHER$OUT_3835_out0 || v$G3_8820_out0;
assign v$MUX5_13175_out0 = v$FF1_8223_out0 ? v$LSBS_7937_out0 : v$_14313_out0;
assign v$MUX5_13176_out0 = v$FF1_8224_out0 ? v$LSBS_7938_out0 : v$_14314_out0;
assign v$N_14070_out0 = v$DIFF_17503_out0;
assign v$N_14071_out0 = v$DIFF_17504_out0;
assign v$N_14072_out0 = v$DIFF_17505_out0;
assign v$N_14073_out0 = v$DIFF_17506_out0;
assign v$NOT$USED1_14379_out0 = v$A1_5790_out1;
assign v$NOT$USED1_14385_out0 = v$A1_5796_out1;
assign v$_16135_out0 = { v$Q0P_16773_out0,v$Q1P_5742_out0 };
assign v$_16136_out0 = { v$Q0P_16774_out0,v$Q1P_5743_out0 };
assign v$EXP$DIFF_17679_out0 = v$EXP$DIFF_14330_out0;
assign v$EXP$DIFF_17680_out0 = v$EXP$DIFF_14331_out0;
assign v$MANTISA$SAME_2436_out0 = v$SAME_6264_out0;
assign v$MANTISA$SAME_2437_out0 = v$SAME_6265_out0;
assign v$MUX3_3107_out0 = v$IS$32$BITS_4148_out0 ? v$_14091_out0 : v$_10038_out0;
assign v$MUX3_3108_out0 = v$IS$32$BITS_4149_out0 ? v$_14092_out0 : v$_10039_out0;
assign v$RAMDOutOut_3187_out0 = v$MUX1_1996_out0;
assign v$RAMDOutOut_3188_out0 = v$MUX1_1997_out0;
assign v$IN_3861_out0 = v$IN_5169_out0;
assign v$IN_3865_out0 = v$IN_5180_out0;
assign v$OUT_3907_out0 = v$G2_12904_out0;
assign v$OUT_3911_out0 = v$G2_12905_out0;
assign v$OUT_3927_out0 = v$G2_12909_out0;
assign v$OUT_3931_out0 = v$G2_12910_out0;
assign v$SEL26_4837_out0 = v$N_14070_out0[7:5];
assign v$SEL26_4838_out0 = v$N_14071_out0[7:5];
assign v$SEL26_4839_out0 = v$N_14072_out0[7:5];
assign v$SEL26_4840_out0 = v$N_14073_out0[7:5];
assign v$SHIFT$AMOUNT_7390_out0 = v$EXP$DIFF_17679_out0;
assign v$SHIFT$AMOUNT_7391_out0 = v$EXP$DIFF_17680_out0;
assign v$_9432_out0 = { v$_16135_out0,v$_2669_out0 };
assign v$_9433_out0 = { v$_16136_out0,v$_2670_out0 };
assign v$MUX13_10363_out0 = v$IS$32$BIT_10862_out0 ? v$DIFF_9088_out0 : v$_7610_out0;
assign v$MUX13_10364_out0 = v$IS$32$BIT_10863_out0 ? v$DIFF_9094_out0 : v$_7611_out0;
assign v$_11811_out0 = { v$_14636_out0,v$MUX5_13175_out0 };
assign v$_11815_out0 = { v$_14640_out0,v$MUX5_13176_out0 };
assign v$SEL25_13454_out0 = v$N_14070_out0[4:0];
assign v$SEL25_13455_out0 = v$N_14071_out0[4:0];
assign v$SEL25_13456_out0 = v$N_14072_out0[4:0];
assign v$SEL25_13457_out0 = v$N_14073_out0[4:0];
assign v$SEL3_1140_out0 = v$SHIFT$AMOUNT_7390_out0[2:2];
assign v$SEL3_1141_out0 = v$SHIFT$AMOUNT_7391_out0[2:2];
assign v$SEL1_2272_out0 = v$SHIFT$AMOUNT_7390_out0[0:0];
assign v$SEL1_2273_out0 = v$SHIFT$AMOUNT_7391_out0[0:0];
assign v$OP1_4100_out0 = v$MUX3_3107_out0;
assign v$OP1_4101_out0 = v$MUX3_3108_out0;
assign v$SEL4_4940_out0 = v$SHIFT$AMOUNT_7390_out0[3:3];
assign v$SEL4_4941_out0 = v$SHIFT$AMOUNT_7391_out0[3:3];
assign v$SEL7_6348_out0 = v$SHIFT$AMOUNT_7390_out0[5:5];
assign v$SEL7_6349_out0 = v$SHIFT$AMOUNT_7391_out0[5:5];
assign v$LOWER$OUT_6422_out0 = v$OUT_3907_out0;
assign v$LOWER$OUT_6423_out0 = v$OUT_3911_out0;
assign v$LOWER$OUT_6424_out0 = v$OUT_3927_out0;
assign v$LOWER$OUT_6425_out0 = v$OUT_3931_out0;
assign v$MUX1_6680_out0 = v$G4_4032_out0 ? v$_11811_out0 : v$MUX2_12041_out0;
assign v$MUX1_6684_out0 = v$G4_4036_out0 ? v$_11815_out0 : v$MUX2_12045_out0;
assign v$SEL1_8717_out0 = v$IN_3861_out0[23:1];
assign v$SEL1_8728_out0 = v$IN_3865_out0[23:1];
assign v$SEL5_12218_out0 = v$SHIFT$AMOUNT_7390_out0[4:4];
assign v$SEL5_12219_out0 = v$SHIFT$AMOUNT_7391_out0[4:4];
assign v$DIFF_12660_out0 = v$MUX13_10363_out0;
assign v$DIFF_12661_out0 = v$MUX13_10364_out0;
assign v$SEL6_13782_out0 = v$SHIFT$AMOUNT_7390_out0[6:6];
assign v$SEL6_13783_out0 = v$SHIFT$AMOUNT_7391_out0[6:6];
assign v$SEL1_15408_out0 = v$IN_3861_out0[22:0];
assign v$SEL1_15419_out0 = v$IN_3865_out0[22:0];
assign v$N_16246_out0 = v$SEL25_13454_out0;
assign v$N_16247_out0 = v$SEL25_13455_out0;
assign v$N_16248_out0 = v$SEL25_13456_out0;
assign v$N_16249_out0 = v$SEL25_13457_out0;
assign v$SEL8_16573_out0 = v$SHIFT$AMOUNT_7390_out0[7:7];
assign v$SEL8_16574_out0 = v$SHIFT$AMOUNT_7391_out0[7:7];
assign v$NUPPER_17364_out0 = v$SEL26_4837_out0;
assign v$NUPPER_17365_out0 = v$SEL26_4838_out0;
assign v$NUPPER_17366_out0 = v$SEL26_4839_out0;
assign v$NUPPER_17367_out0 = v$SEL26_4840_out0;
assign v$UART$DOUT_17461_out0 = v$RAMDOutOut_3187_out0;
assign v$UART$DOUT_17462_out0 = v$RAMDOutOut_3188_out0;
assign v$SEL2_18358_out0 = v$SHIFT$AMOUNT_7390_out0[1:1];
assign v$SEL2_18359_out0 = v$SHIFT$AMOUNT_7391_out0[1:1];
assign v$DIFF_292_out0 = v$DIFF_12660_out0;
assign v$DIFF_293_out0 = v$DIFF_12661_out0;
assign v$EN_1338_out0 = v$SEL5_12218_out0;
assign v$EN_1339_out0 = v$SEL4_4940_out0;
assign v$EN_1341_out0 = v$SEL5_12219_out0;
assign v$EN_1342_out0 = v$SEL4_4941_out0;
assign v$EQ3_1816_out0 = v$N_16246_out0 == 5'h2;
assign v$EQ3_1817_out0 = v$N_16247_out0 == 5'h2;
assign v$EQ3_1818_out0 = v$N_16248_out0 == 5'h2;
assign v$EQ3_1819_out0 = v$N_16249_out0 == 5'h2;
assign v$MUX3_1960_out0 = v$G8_1889_out0 ? v$_13307_out0 : v$MUX1_6680_out0;
assign v$MUX3_1964_out0 = v$G8_1893_out0 ? v$_13311_out0 : v$MUX1_6684_out0;
assign v$EQ24_2536_out0 = v$N_16246_out0 == 5'h17;
assign v$EQ24_2537_out0 = v$N_16247_out0 == 5'h17;
assign v$EQ24_2538_out0 = v$N_16248_out0 == 5'h17;
assign v$EQ24_2539_out0 = v$N_16249_out0 == 5'h17;
assign v$EQ22_2836_out0 = v$N_16246_out0 == 5'h15;
assign v$EQ22_2837_out0 = v$N_16247_out0 == 5'h15;
assign v$EQ22_2838_out0 = v$N_16248_out0 == 5'h15;
assign v$EQ22_2839_out0 = v$N_16249_out0 == 5'h15;
assign v$EQ23_3194_out0 = v$N_16246_out0 == 5'h16;
assign v$EQ23_3195_out0 = v$N_16247_out0 == 5'h16;
assign v$EQ23_3196_out0 = v$N_16248_out0 == 5'h16;
assign v$EQ23_3197_out0 = v$N_16249_out0 == 5'h16;
assign v$EQ5_3315_out0 = v$N_16246_out0 == 5'h4;
assign v$EQ5_3316_out0 = v$N_16247_out0 == 5'h4;
assign v$EQ5_3317_out0 = v$N_16248_out0 == 5'h4;
assign v$EQ5_3318_out0 = v$N_16249_out0 == 5'h4;
assign v$EQ21_3324_out0 = v$N_16246_out0 == 5'h14;
assign v$EQ21_3325_out0 = v$N_16247_out0 == 5'h14;
assign v$EQ21_3326_out0 = v$N_16248_out0 == 5'h14;
assign v$EQ21_3327_out0 = v$N_16249_out0 == 5'h14;
assign v$A_3463_out0 = v$OP1_4100_out0;
assign v$EQ7_4085_out0 = v$N_16246_out0 == 5'h6;
assign v$EQ7_4086_out0 = v$N_16247_out0 == 5'h6;
assign v$EQ7_4087_out0 = v$N_16248_out0 == 5'h6;
assign v$EQ7_4088_out0 = v$N_16249_out0 == 5'h6;
assign v$_4267_out0 = { v$C2_125_out0,v$SEL1_15408_out0 };
assign v$_4278_out0 = { v$C2_136_out0,v$SEL1_15419_out0 };
assign v$EN_4755_out0 = v$SEL3_1140_out0;
assign v$EN_4757_out0 = v$SEL3_1141_out0;
assign v$EN_5214_out0 = v$SEL1_2272_out0;
assign v$EN_5216_out0 = v$SEL1_2273_out0;
assign v$EQ14_5401_out0 = v$N_16246_out0 == 5'hd;
assign v$EQ14_5402_out0 = v$N_16247_out0 == 5'hd;
assign v$EQ14_5403_out0 = v$N_16248_out0 == 5'hd;
assign v$EQ14_5404_out0 = v$N_16249_out0 == 5'hd;
assign v$A_5418_out0 = v$OP1_4101_out0;
assign v$EQ6_5425_out0 = v$N_16246_out0 == 5'h5;
assign v$EQ6_5426_out0 = v$N_16247_out0 == 5'h5;
assign v$EQ6_5427_out0 = v$N_16248_out0 == 5'h5;
assign v$EQ6_5428_out0 = v$N_16249_out0 == 5'h5;
assign v$EQ19_5442_out0 = v$N_16246_out0 == 5'h12;
assign v$EQ19_5443_out0 = v$N_16247_out0 == 5'h12;
assign v$EQ19_5444_out0 = v$N_16248_out0 == 5'h12;
assign v$EQ19_5445_out0 = v$N_16249_out0 == 5'h12;
assign v$EQ17_5879_out0 = v$N_16246_out0 == 5'h10;
assign v$EQ17_5880_out0 = v$N_16247_out0 == 5'h10;
assign v$EQ17_5881_out0 = v$N_16248_out0 == 5'h10;
assign v$EQ17_5882_out0 = v$N_16249_out0 == 5'h10;
assign v$EQ10_5892_out0 = v$N_16246_out0 == 5'h8;
assign v$EQ10_5893_out0 = v$N_16247_out0 == 5'h8;
assign v$EQ10_5894_out0 = v$N_16248_out0 == 5'h8;
assign v$EQ10_5895_out0 = v$N_16249_out0 == 5'h8;
assign v$EQ11_6143_out0 = v$N_16246_out0 == 5'ha;
assign v$EQ11_6144_out0 = v$N_16247_out0 == 5'ha;
assign v$EQ11_6145_out0 = v$N_16248_out0 == 5'ha;
assign v$EQ11_6146_out0 = v$N_16249_out0 == 5'ha;
assign v$SEL28_7327_out0 = v$NUPPER_17364_out0[1:1];
assign v$SEL28_7328_out0 = v$NUPPER_17365_out0[1:1];
assign v$SEL28_7329_out0 = v$NUPPER_17366_out0[1:1];
assign v$SEL28_7330_out0 = v$NUPPER_17367_out0[1:1];
assign v$EN_7877_out0 = v$SEL2_18358_out0;
assign v$EN_7879_out0 = v$SEL2_18359_out0;
assign v$RAMDOUT_7917_out0 = v$UART$DOUT_17461_out0;
assign v$RAMDOUT_7918_out0 = v$UART$DOUT_17462_out0;
assign v$EQ16_8286_out0 = v$N_16246_out0 == 5'hf;
assign v$EQ16_8287_out0 = v$N_16247_out0 == 5'hf;
assign v$EQ16_8288_out0 = v$N_16248_out0 == 5'hf;
assign v$EQ16_8289_out0 = v$N_16249_out0 == 5'hf;
assign v$_9002_out0 = { v$SEL1_8717_out0,v$C1_5983_out0 };
assign v$_9013_out0 = { v$SEL1_8728_out0,v$C1_5994_out0 };
assign v$EQ13_9515_out0 = v$N_16246_out0 == 5'hc;
assign v$EQ13_9516_out0 = v$N_16247_out0 == 5'hc;
assign v$EQ13_9517_out0 = v$N_16248_out0 == 5'hc;
assign v$EQ13_9518_out0 = v$N_16249_out0 == 5'hc;
assign v$EQ20_9946_out0 = v$N_16246_out0 == 5'h13;
assign v$EQ20_9947_out0 = v$N_16247_out0 == 5'h13;
assign v$EQ20_9948_out0 = v$N_16248_out0 == 5'h13;
assign v$EQ20_9949_out0 = v$N_16249_out0 == 5'h13;
assign v$EQ18_12806_out0 = v$N_16246_out0 == 5'h11;
assign v$EQ18_12807_out0 = v$N_16247_out0 == 5'h11;
assign v$EQ18_12808_out0 = v$N_16248_out0 == 5'h11;
assign v$EQ18_12809_out0 = v$N_16249_out0 == 5'h11;
assign v$EQ1_13414_out0 = v$N_16246_out0 == 5'h0;
assign v$EQ1_13415_out0 = v$N_16247_out0 == 5'h0;
assign v$EQ1_13416_out0 = v$N_16248_out0 == 5'h0;
assign v$EQ1_13417_out0 = v$N_16249_out0 == 5'h0;
assign v$EQ9_13775_out0 = v$N_16246_out0 == 5'h9;
assign v$EQ9_13776_out0 = v$N_16247_out0 == 5'h9;
assign v$EQ9_13777_out0 = v$N_16248_out0 == 5'h9;
assign v$EQ9_13778_out0 = v$N_16249_out0 == 5'h9;
assign v$EQ12_13838_out0 = v$N_16246_out0 == 5'hb;
assign v$EQ12_13839_out0 = v$N_16247_out0 == 5'hb;
assign v$EQ12_13840_out0 = v$N_16248_out0 == 5'hb;
assign v$EQ12_13841_out0 = v$N_16249_out0 == 5'hb;
assign v$EQ2_14208_out0 = v$N_16246_out0 == 5'h1;
assign v$EQ2_14209_out0 = v$N_16247_out0 == 5'h1;
assign v$EQ2_14210_out0 = v$N_16248_out0 == 5'h1;
assign v$EQ2_14211_out0 = v$N_16249_out0 == 5'h1;
assign v$EQ8_14414_out0 = v$N_16246_out0 == 5'h7;
assign v$EQ8_14415_out0 = v$N_16247_out0 == 5'h7;
assign v$EQ8_14416_out0 = v$N_16248_out0 == 5'h7;
assign v$EQ8_14417_out0 = v$N_16249_out0 == 5'h7;
assign v$EQ15_15965_out0 = v$N_16246_out0 == 5'he;
assign v$EQ15_15966_out0 = v$N_16247_out0 == 5'he;
assign v$EQ15_15967_out0 = v$N_16248_out0 == 5'he;
assign v$EQ15_15968_out0 = v$N_16249_out0 == 5'he;
assign v$G1_16032_out0 = v$SEL7_6348_out0 || v$SEL6_13782_out0;
assign v$G1_16033_out0 = v$SEL7_6349_out0 || v$SEL6_13783_out0;
assign v$SEL27_16304_out0 = v$NUPPER_17364_out0[0:0];
assign v$SEL27_16305_out0 = v$NUPPER_17365_out0[0:0];
assign v$SEL27_16306_out0 = v$NUPPER_17366_out0[0:0];
assign v$SEL27_16307_out0 = v$NUPPER_17367_out0[0:0];
assign v$SEL29_16594_out0 = v$NUPPER_17364_out0[2:2];
assign v$SEL29_16595_out0 = v$NUPPER_17365_out0[2:2];
assign v$SEL29_16596_out0 = v$NUPPER_17366_out0[2:2];
assign v$SEL29_16597_out0 = v$NUPPER_17367_out0[2:2];
assign v$G2_18239_out0 = v$HIGHER$SAME_9132_out0 && v$LOWER$OUT_6422_out0;
assign v$G2_18240_out0 = v$HIGHER$SAME_9133_out0 && v$LOWER$OUT_6423_out0;
assign v$G2_18241_out0 = v$HIGHER$SAME_9134_out0 && v$LOWER$OUT_6424_out0;
assign v$G2_18242_out0 = v$HIGHER$SAME_9135_out0 && v$LOWER$OUT_6425_out0;
assign v$EQ4_18599_out0 = v$N_16246_out0 == 5'h3;
assign v$EQ4_18600_out0 = v$N_16247_out0 == 5'h3;
assign v$EQ4_18601_out0 = v$N_16248_out0 == 5'h3;
assign v$EQ4_18602_out0 = v$N_16249_out0 == 5'h3;
assign v$RAMDOUT_68_out0 = v$RAMDOUT_7917_out0;
assign v$RAMDOUT_69_out0 = v$RAMDOUT_7918_out0;
assign v$MUX1_2371_out0 = v$LEFT$SHIT_3063_out0 ? v$_4267_out0 : v$_9002_out0;
assign v$MUX1_2382_out0 = v$LEFT$SHIT_3074_out0 ? v$_4278_out0 : v$_9013_out0;
assign v$DIFF_2820_out0 = v$DIFF_292_out0;
assign v$DIFF_2821_out0 = v$DIFF_293_out0;
assign v$OUT_3179_out0 = v$MUX3_1960_out0;
assign v$OUT_3183_out0 = v$MUX3_1964_out0;
assign v$G1_8792_out0 = v$SEL27_16304_out0 || v$SEL28_7327_out0;
assign v$G1_8793_out0 = v$SEL27_16305_out0 || v$SEL28_7328_out0;
assign v$G1_8794_out0 = v$SEL27_16306_out0 || v$SEL28_7329_out0;
assign v$G1_8795_out0 = v$SEL27_16307_out0 || v$SEL28_7330_out0;
assign v$G3_13061_out0 = v$HIGHER$OUT_7785_out0 || v$G2_18239_out0;
assign v$G3_13062_out0 = v$HIGHER$OUT_7786_out0 || v$G2_18240_out0;
assign v$G3_13063_out0 = v$HIGHER$OUT_7787_out0 || v$G2_18241_out0;
assign v$G3_13064_out0 = v$HIGHER$OUT_7788_out0 || v$G2_18242_out0;
assign v$A_14255_out0 = v$A_3463_out0;
assign v$A_14801_out0 = v$A_5418_out0;
assign v$G2_17414_out0 = v$G1_16032_out0 || v$SEL8_16573_out0;
assign v$G2_17415_out0 = v$G1_16033_out0 || v$SEL8_16574_out0;
assign v$MULTIPLIER_3669_out0 = v$A_14801_out0;
assign v$MULTIPLIER_3671_out0 = v$A_14801_out0;
assign v$MULTIPLIER_3672_out0 = v$A_14801_out0;
assign v$MULTIPLIER_3673_out0 = v$A_14801_out0;
assign v$MULTIPLIER_3674_out0 = v$A_14801_out0;
assign v$MULTIPLIER_3675_out0 = v$A_14801_out0;
assign v$MULTIPLIER_3676_out0 = v$A_14801_out0;
assign v$MULTIPLIER_3677_out0 = v$A_14801_out0;
assign v$MULTIPLIER_3678_out0 = v$A_14801_out0;
assign v$MULTIPLIER_3679_out0 = v$A_14801_out0;
assign v$MULTIPLIER_3680_out0 = v$A_14801_out0;
assign v$RAMDOUT_5423_out0 = v$RAMDOUT_68_out0;
assign v$RAMDOUT_5424_out0 = v$RAMDOUT_69_out0;
assign v$MULTIPLIER_6355_out0 = v$A_14801_out0;
assign v$SHIFT$AMOUNT_7387_out0 = v$DIFF_2820_out0;
assign v$SHIFT$AMOUNT_7388_out0 = v$DIFF_2820_out0;
assign v$SHIFT$AMOUNT_7392_out0 = v$DIFF_2821_out0;
assign v$SHIFT$AMOUNT_7393_out0 = v$DIFF_2821_out0;
assign v$OUT_8937_out0 = v$G3_13061_out0;
assign v$OUT_8938_out0 = v$G3_13062_out0;
assign v$OUT_8939_out0 = v$G3_13063_out0;
assign v$OUT_8940_out0 = v$G3_13064_out0;
assign v$SEL5_10328_out0 = v$A_14255_out0[23:1];
assign v$G2_11902_out0 = v$G1_8792_out0 || v$SEL29_16594_out0;
assign v$G2_11903_out0 = v$G1_8793_out0 || v$SEL29_16595_out0;
assign v$G2_11904_out0 = v$G1_8794_out0 || v$SEL29_16596_out0;
assign v$G2_11905_out0 = v$G1_8795_out0 || v$SEL29_16597_out0;
assign v$OUT_14505_out0 = v$OUT_3179_out0;
assign v$OUT_14506_out0 = v$OUT_3183_out0;
assign v$MUX2_18577_out0 = v$EN_5214_out0 ? v$MUX1_2371_out0 : v$IN_3861_out0;
assign v$MUX2_18579_out0 = v$EN_5216_out0 ? v$MUX1_2382_out0 : v$IN_3865_out0;
assign v$SEL3_1137_out0 = v$SHIFT$AMOUNT_7387_out0[2:2];
assign v$SEL3_1138_out0 = v$SHIFT$AMOUNT_7388_out0[2:2];
assign v$SEL3_1142_out0 = v$SHIFT$AMOUNT_7392_out0[2:2];
assign v$SEL3_1143_out0 = v$SHIFT$AMOUNT_7393_out0[2:2];
assign v$_1158_out0 = { v$SEL5_10328_out0,v$C6_8836_out0 };
assign v$SEL1_2269_out0 = v$SHIFT$AMOUNT_7387_out0[0:0];
assign v$SEL1_2270_out0 = v$SHIFT$AMOUNT_7388_out0[0:0];
assign v$SEL1_2274_out0 = v$SHIFT$AMOUNT_7392_out0[0:0];
assign v$SEL1_2275_out0 = v$SHIFT$AMOUNT_7393_out0[0:0];
assign v$G3_4724_out0 = v$OUT_8938_out0 && v$SAME$H_8915_out0;
assign v$G3_4725_out0 = v$OUT_8940_out0 && v$SAME$H_8916_out0;
assign v$SEL4_4937_out0 = v$SHIFT$AMOUNT_7387_out0[3:3];
assign v$SEL4_4938_out0 = v$SHIFT$AMOUNT_7388_out0[3:3];
assign v$SEL4_4942_out0 = v$SHIFT$AMOUNT_7392_out0[3:3];
assign v$SEL4_4943_out0 = v$SHIFT$AMOUNT_7393_out0[3:3];
assign v$SEL7_6345_out0 = v$SHIFT$AMOUNT_7387_out0[5:5];
assign v$SEL7_6346_out0 = v$SHIFT$AMOUNT_7388_out0[5:5];
assign v$SEL7_6350_out0 = v$SHIFT$AMOUNT_7392_out0[5:5];
assign v$SEL7_6351_out0 = v$SHIFT$AMOUNT_7393_out0[5:5];
assign v$OP2_10191_out0 = v$OUT_14505_out0;
assign v$OP2_10192_out0 = v$OUT_14506_out0;
assign v$OP2_10374_out0 = v$MULTIPLIER_3669_out0;
assign v$OP2_10375_out0 = v$MULTIPLIER_6355_out0;
assign v$OP2_10376_out0 = v$MULTIPLIER_3671_out0;
assign v$OP2_10377_out0 = v$MULTIPLIER_3672_out0;
assign v$OP2_10378_out0 = v$MULTIPLIER_3673_out0;
assign v$OP2_10379_out0 = v$MULTIPLIER_3674_out0;
assign v$OP2_10380_out0 = v$MULTIPLIER_3675_out0;
assign v$OP2_10381_out0 = v$MULTIPLIER_3676_out0;
assign v$OP2_10382_out0 = v$MULTIPLIER_3677_out0;
assign v$OP2_10383_out0 = v$MULTIPLIER_3678_out0;
assign v$OP2_10384_out0 = v$MULTIPLIER_3679_out0;
assign v$OP2_10385_out0 = v$MULTIPLIER_3680_out0;
assign v$MUX2_11980_out0 = v$G24_17931_out0 ? v$RAMDOUT_5423_out0 : v$RMN_6155_out0;
assign v$MUX2_11981_out0 = v$G24_17932_out0 ? v$RAMDOUT_5424_out0 : v$RMN_6156_out0;
assign v$SEL5_12215_out0 = v$SHIFT$AMOUNT_7387_out0[4:4];
assign v$SEL5_12216_out0 = v$SHIFT$AMOUNT_7388_out0[4:4];
assign v$SEL5_12220_out0 = v$SHIFT$AMOUNT_7392_out0[4:4];
assign v$SEL5_12221_out0 = v$SHIFT$AMOUNT_7393_out0[4:4];
assign v$SEL6_13779_out0 = v$SHIFT$AMOUNT_7387_out0[6:6];
assign v$SEL6_13780_out0 = v$SHIFT$AMOUNT_7388_out0[6:6];
assign v$SEL6_13784_out0 = v$SHIFT$AMOUNT_7392_out0[6:6];
assign v$SEL6_13785_out0 = v$SHIFT$AMOUNT_7393_out0[6:6];
assign v$OUT_14923_out0 = v$MUX2_18577_out0;
assign v$OUT_14934_out0 = v$MUX2_18579_out0;
assign v$SEL8_16570_out0 = v$SHIFT$AMOUNT_7387_out0[7:7];
assign v$SEL8_16571_out0 = v$SHIFT$AMOUNT_7388_out0[7:7];
assign v$SEL8_16575_out0 = v$SHIFT$AMOUNT_7392_out0[7:7];
assign v$SEL8_16576_out0 = v$SHIFT$AMOUNT_7393_out0[7:7];
assign v$SEL2_18355_out0 = v$SHIFT$AMOUNT_7387_out0[1:1];
assign v$SEL2_18356_out0 = v$SHIFT$AMOUNT_7388_out0[1:1];
assign v$SEL2_18360_out0 = v$SHIFT$AMOUNT_7392_out0[1:1];
assign v$SEL2_18361_out0 = v$SHIFT$AMOUNT_7393_out0[1:1];
assign v$EN_1331_out0 = v$SEL5_12215_out0;
assign v$EN_1332_out0 = v$SEL4_4937_out0;
assign v$EN_1333_out0 = v$SEL5_12216_out0;
assign v$EN_1334_out0 = v$SEL4_4938_out0;
assign v$EN_1345_out0 = v$SEL5_12220_out0;
assign v$EN_1346_out0 = v$SEL4_4942_out0;
assign v$EN_1347_out0 = v$SEL5_12221_out0;
assign v$EN_1348_out0 = v$SEL4_4943_out0;
assign v$EN_4751_out0 = v$SEL3_1137_out0;
assign v$EN_4752_out0 = v$SEL3_1138_out0;
assign v$EN_4760_out0 = v$SEL3_1142_out0;
assign v$EN_4761_out0 = v$SEL3_1143_out0;
assign v$IN_5171_out0 = v$OUT_14923_out0;
assign v$IN_5182_out0 = v$OUT_14934_out0;
assign v$EN_5210_out0 = v$SEL1_2269_out0;
assign v$EN_5211_out0 = v$SEL1_2270_out0;
assign v$EN_5223_out0 = v$SEL1_2274_out0;
assign v$EN_5224_out0 = v$SEL1_2275_out0;
assign v$EN_7873_out0 = v$SEL2_18355_out0;
assign v$EN_7874_out0 = v$SEL2_18356_out0;
assign v$EN_7882_out0 = v$SEL2_18360_out0;
assign v$EN_7883_out0 = v$SEL2_18361_out0;
assign v$OP2_15055_out0 = v$OP2_10191_out0;
assign v$OP2_15056_out0 = v$OP2_10192_out0;
assign v$G1_15586_out0 = v$G3_4724_out0 || v$OUT_8937_out0;
assign v$G1_15587_out0 = v$G3_4725_out0 || v$OUT_8939_out0;
assign v$G1_16029_out0 = v$SEL7_6345_out0 || v$SEL6_13779_out0;
assign v$G1_16030_out0 = v$SEL7_6346_out0 || v$SEL6_13780_out0;
assign v$G1_16034_out0 = v$SEL7_6350_out0 || v$SEL6_13784_out0;
assign v$G1_16035_out0 = v$SEL7_6351_out0 || v$SEL6_13785_out0;
assign v$REGDIN_18379_out0 = v$MUX2_11980_out0;
assign v$REGDIN_18380_out0 = v$MUX2_11981_out0;
assign v$OUT_3840_out0 = v$G1_15586_out0;
assign v$OUT_3841_out0 = v$G1_15587_out0;
assign v$OP2_7579_out0 = v$OP2_15055_out0;
assign v$OP2_7580_out0 = v$OP2_15056_out0;
assign v$IN_11785_out0 = v$IN_5171_out0;
assign v$IN_11787_out0 = v$IN_5182_out0;
assign v$REGDIN_16498_out0 = v$REGDIN_18379_out0;
assign v$REGDIN_16499_out0 = v$REGDIN_18380_out0;
assign v$G2_17411_out0 = v$G1_16029_out0 || v$SEL8_16570_out0;
assign v$G2_17412_out0 = v$G1_16030_out0 || v$SEL8_16571_out0;
assign v$G2_17416_out0 = v$G1_16034_out0 || v$SEL8_16575_out0;
assign v$G2_17417_out0 = v$G1_16035_out0 || v$SEL8_16576_out0;
assign v$SEL1_8719_out0 = v$IN_11785_out0[23:2];
assign v$SEL1_8730_out0 = v$IN_11787_out0[23:2];
assign v$XOR1_9542_out0 = v$OP2_7579_out0 ^ v$MUX1_17728_out0;
assign v$XOR1_9543_out0 = v$OP2_7580_out0 ^ v$MUX1_17729_out0;
assign v$B_11720_out0 = v$OP2_7579_out0;
assign v$B_11721_out0 = v$OP2_7580_out0;
assign v$SEL1_15410_out0 = v$IN_11785_out0[21:0];
assign v$SEL1_15421_out0 = v$IN_11787_out0[21:0];
assign v$A$MANTISA$LARGER_16027_out0 = v$OUT_3840_out0;
assign v$A$MANTISA$LARGER_16028_out0 = v$OUT_3841_out0;
assign v$_4269_out0 = { v$C2_127_out0,v$SEL1_15410_out0 };
assign v$_4280_out0 = { v$C2_138_out0,v$SEL1_15421_out0 };
assign v$_9004_out0 = { v$SEL1_8719_out0,v$C1_5985_out0 };
assign v$_9015_out0 = { v$SEL1_8730_out0,v$C1_5996_out0 };
assign {v$A1_9430_out1,v$A1_9430_out0 } = v$OP1_5416_out0 + v$XOR1_9542_out0 + v$MUX2_12234_out0;
assign {v$A1_9431_out1,v$A1_9431_out0 } = v$OP1_5417_out0 + v$XOR1_9543_out0 + v$MUX2_12235_out0;
assign v$B_10007_out0 = v$B_11720_out0;
assign v$B_10008_out0 = v$B_11721_out0;
assign v$G7_18641_out0 = v$A$MANTISA$LARGER_16027_out0 && v$EXP$SAME_903_out0;
assign v$G7_18642_out0 = v$A$MANTISA$LARGER_16028_out0 && v$EXP$SAME_904_out0;
assign v$MUX1_2373_out0 = v$LEFT$SHIT_3065_out0 ? v$_4269_out0 : v$_9004_out0;
assign v$MUX1_2384_out0 = v$LEFT$SHIT_3076_out0 ? v$_4280_out0 : v$_9015_out0;
assign v$ADDEROUT_3504_out0 = v$A1_9430_out0;
assign v$ADDEROUT_3505_out0 = v$A1_9431_out0;
assign v$_5232_out0 = v$B_10007_out0[7:4];
assign v$_5233_out0 = v$B_10008_out0[7:4];
assign v$_6343_out0 = v$B_10007_out0[11:8];
assign v$_6344_out0 = v$B_10008_out0[11:8];
assign v$G9_16920_out0 = v$A$EXP$LARGER_18245_out0 || v$G7_18641_out0;
assign v$G9_16921_out0 = v$A$EXP$LARGER_18246_out0 || v$G7_18642_out0;
assign v$_18249_out0 = v$B_10007_out0[15:12];
assign v$_18250_out0 = v$B_10008_out0[15:12];
assign v$_18607_out0 = v$B_10007_out0[3:0];
assign v$_18608_out0 = v$B_10008_out0[3:0];
assign v$_54_out0 = v$_18607_out0[1:0];
assign v$_54_out1 = v$_18607_out0[3:2];
assign v$_55_out0 = v$_18608_out0[1:0];
assign v$_55_out1 = v$_18608_out0[3:2];
assign v$_229_out0 = v$_5232_out0[1:0];
assign v$_229_out1 = v$_5232_out0[3:2];
assign v$_230_out0 = v$_5233_out0[1:0];
assign v$_230_out1 = v$_5233_out0[3:2];
assign v$_1473_out0 = v$_18249_out0[1:0];
assign v$_1473_out1 = v$_18249_out0[3:2];
assign v$_1474_out0 = v$_18250_out0[1:0];
assign v$_1474_out1 = v$_18250_out0[3:2];
assign v$MUX2_2479_out0 = v$EN_7877_out0 ? v$MUX1_2373_out0 : v$IN_11785_out0;
assign v$MUX2_2481_out0 = v$EN_7879_out0 ? v$MUX1_2384_out0 : v$IN_11787_out0;
assign v$_7467_out0 = v$_6343_out0[1:0];
assign v$_7467_out1 = v$_6343_out0[3:2];
assign v$_7468_out0 = v$_6344_out0[1:0];
assign v$_7468_out1 = v$_6344_out0[3:2];
assign v$IS$A$LARGER_16832_out0 = v$G9_16920_out0;
assign v$IS$A$LARGER_16833_out0 = v$G9_16921_out0;
assign v$G8_246_out0 = v$IS$A$LARGER_16832_out0 || v$IS$SUB_4443_out0;
assign v$G8_247_out0 = v$IS$A$LARGER_16833_out0 || v$IS$SUB_4444_out0;
assign v$MUX11_1204_out0 = v$IS$A$LARGER_16832_out0 ? v$SEL5_313_out0 : v$G1_15142_out0;
assign v$MUX11_1205_out0 = v$IS$A$LARGER_16833_out0 ? v$SEL5_314_out0 : v$G1_15143_out0;
assign v$_5040_out0 = v$_54_out1[0:0];
assign v$_5040_out1 = v$_54_out1[1:1];
assign v$_5041_out0 = v$_55_out1[0:0];
assign v$_5041_out1 = v$_55_out1[1:1];
assign v$MUX15_7008_out0 = v$IS$A$LARGER_16832_out0 ? v$A_3242_out0 : v$B_17746_out0;
assign v$MUX15_7009_out0 = v$IS$A$LARGER_16833_out0 ? v$A_3243_out0 : v$B_17747_out0;
assign v$IS$A$LARGER_7072_out0 = v$IS$A$LARGER_16832_out0;
assign v$IS$A$LARGER_7073_out0 = v$IS$A$LARGER_16833_out0;
assign v$_7395_out0 = v$_229_out1[0:0];
assign v$_7395_out1 = v$_229_out1[1:1];
assign v$_7396_out0 = v$_230_out1[0:0];
assign v$_7396_out1 = v$_230_out1[1:1];
assign v$_9070_out0 = v$_229_out0[0:0];
assign v$_9070_out1 = v$_229_out0[1:1];
assign v$_9071_out0 = v$_230_out0[0:0];
assign v$_9071_out1 = v$_230_out0[1:1];
assign v$_9110_out0 = v$_7467_out0[0:0];
assign v$_9110_out1 = v$_7467_out0[1:1];
assign v$_9111_out0 = v$_7468_out0[0:0];
assign v$_9111_out1 = v$_7468_out0[1:1];
assign v$_14645_out0 = v$_54_out0[0:0];
assign v$_14645_out1 = v$_54_out0[1:1];
assign v$_14646_out0 = v$_55_out0[0:0];
assign v$_14646_out1 = v$_55_out0[1:1];
assign v$OUT_14925_out0 = v$MUX2_2479_out0;
assign v$OUT_14936_out0 = v$MUX2_2481_out0;
assign v$_15188_out0 = v$_1473_out0[0:0];
assign v$_15188_out1 = v$_1473_out0[1:1];
assign v$_15189_out0 = v$_1474_out0[0:0];
assign v$_15189_out1 = v$_1474_out0[1:1];
assign v$_15320_out0 = v$_1473_out1[0:0];
assign v$_15320_out1 = v$_1473_out1[1:1];
assign v$_15321_out0 = v$_1474_out1[0:0];
assign v$_15321_out1 = v$_1474_out1[1:1];
assign v$G2_15542_out0 = v$IS$A$LARGER_16832_out0 && v$IS$SUB_4443_out0;
assign v$G2_15543_out0 = v$IS$A$LARGER_16833_out0 && v$IS$SUB_4444_out0;
assign v$_16137_out0 = v$_7467_out1[0:0];
assign v$_16137_out1 = v$_7467_out1[1:1];
assign v$_16138_out0 = v$_7468_out1[0:0];
assign v$_16138_out1 = v$_7468_out1[1:1];
assign v$MUX16_18527_out0 = v$IS$A$LARGER_16832_out0 ? v$A_3242_out0 : v$B_17746_out0;
assign v$MUX16_18528_out0 = v$IS$A$LARGER_16833_out0 ? v$A_3243_out0 : v$B_17747_out0;
assign v$G14_1673_out0 = v$_16550_out1 && v$_15188_out1;
assign v$G14_1674_out0 = v$_16551_out1 && v$_15189_out1;
assign v$G13_1689_out0 = v$_16550_out0 && v$_15188_out0;
assign v$G13_1690_out0 = v$_16551_out0 && v$_15189_out0;
assign v$G5_2235_out0 = v$_4019_out0 && v$_9070_out0;
assign v$G5_2236_out0 = v$_4020_out0 && v$_9071_out0;
assign v$G6_2247_out0 = v$_4019_out1 && v$_9070_out1;
assign v$G6_2248_out0 = v$_4020_out1 && v$_9071_out1;
assign v$G9_3441_out0 = v$_330_out0 && v$_9110_out0;
assign v$G9_3442_out0 = v$_331_out0 && v$_9111_out0;
assign v$A$IS$OP1_5005_out0 = v$G8_246_out0;
assign v$A$IS$OP1_5006_out0 = v$G8_247_out0;
assign v$IN_5170_out0 = v$OUT_14925_out0;
assign v$IN_5181_out0 = v$OUT_14936_out0;
assign v$SEL17_5388_out0 = v$MUX16_18527_out0[14:7];
assign v$SEL17_5389_out0 = v$MUX16_18528_out0[14:7];
assign v$G11_8202_out0 = v$_4892_out0 && v$_16137_out0;
assign v$G11_8203_out0 = v$_4893_out0 && v$_16138_out0;
assign v$G2_9078_out0 = v$_11056_out1 && v$_14645_out1;
assign v$G2_9079_out0 = v$_11057_out1 && v$_14646_out1;
assign v$G8_9083_out0 = v$_10244_out1 && v$_7395_out1;
assign v$G8_9084_out0 = v$_10245_out1 && v$_7396_out1;
assign v$IS$A$LARGER_10444_out0 = v$IS$A$LARGER_7072_out0;
assign v$IS$A$LARGER_10445_out0 = v$IS$A$LARGER_7073_out0;
assign v$G4_11870_out0 = v$G2_15542_out0 && v$G5_15791_out0;
assign v$G4_11871_out0 = v$G2_15543_out0 && v$G5_15792_out0;
assign v$SUBTRACTION$SIGN_11872_out0 = v$MUX11_1204_out0;
assign v$SUBTRACTION$SIGN_11873_out0 = v$MUX11_1205_out0;
assign v$G1_12124_out0 = v$_11056_out0 && v$_14645_out0;
assign v$G1_12125_out0 = v$_11057_out0 && v$_14646_out0;
assign v$G7_12203_out0 = v$_10244_out0 && v$_7395_out0;
assign v$G7_12204_out0 = v$_10245_out0 && v$_7396_out0;
assign v$G3_12948_out0 = v$_5405_out0 && v$_5040_out0;
assign v$G3_12949_out0 = v$_5406_out0 && v$_5041_out0;
assign v$G12_13795_out0 = v$_4892_out1 && v$_16137_out1;
assign v$G12_13796_out0 = v$_4893_out1 && v$_16138_out1;
assign v$G4_14501_out0 = v$_5405_out1 && v$_5040_out1;
assign v$G4_14502_out0 = v$_5406_out1 && v$_5041_out1;
assign v$G15_14582_out0 = v$_3118_out0 && v$_15320_out0;
assign v$G15_14583_out0 = v$_3119_out0 && v$_15321_out0;
assign v$SEL3_17773_out0 = v$MUX15_7008_out0[14:7];
assign v$SEL3_17774_out0 = v$MUX15_7009_out0[14:7];
assign v$SEL18_18251_out0 = v$MUX16_18527_out0[14:10];
assign v$SEL18_18252_out0 = v$MUX16_18528_out0[14:10];
assign v$G10_18485_out0 = v$_330_out1 && v$_9110_out1;
assign v$G10_18486_out0 = v$_331_out1 && v$_9111_out1;
assign v$G16_18781_out0 = v$_3118_out1 && v$_15320_out1;
assign v$G16_18782_out0 = v$_3119_out1 && v$_15321_out1;
assign v$MUX9_2458_out0 = v$A$IS$OP1_5005_out0 ? v$B$MANTISA_15588_out0 : v$A$MANTISA_3756_out0;
assign v$MUX9_2459_out0 = v$A$IS$OP1_5006_out0 ? v$B$MANTISA_15589_out0 : v$A$MANTISA_3757_out0;
assign v$_3145_out0 = { v$G15_14582_out0,v$G16_18781_out0 };
assign v$_3146_out0 = { v$G15_14583_out0,v$G16_18782_out0 };
assign v$_9457_out0 = { v$G7_12203_out0,v$G8_9083_out0 };
assign v$_9458_out0 = { v$G7_12204_out0,v$G8_9084_out0 };
assign v$_10974_out0 = { v$G3_12948_out0,v$G4_14501_out0 };
assign v$_10975_out0 = { v$G3_12949_out0,v$G4_14502_out0 };
assign v$SINGLE$PRECISION$EXPONENT_11046_out0 = v$SEL3_17773_out0;
assign v$SINGLE$PRECISION$EXPONENT_11047_out0 = v$SEL3_17774_out0;
assign v$MUX3_12800_out0 = v$A$IS$OP1_5005_out0 ? v$A$MANTISA_3756_out0 : v$B$MANTISA_15588_out0;
assign v$MUX3_12801_out0 = v$A$IS$OP1_5006_out0 ? v$A$MANTISA_3757_out0 : v$B$MANTISA_15589_out0;
assign v$EXPONENT_13686_out0 = v$SEL17_5388_out0;
assign v$EXPONENT_13687_out0 = v$SEL17_5389_out0;
assign v$_14166_out0 = { v$G1_12124_out0,v$G2_9078_out0 };
assign v$_14167_out0 = { v$G1_12125_out0,v$G2_9079_out0 };
assign v$_14212_out0 = { v$G5_2235_out0,v$G6_2247_out0 };
assign v$_14213_out0 = { v$G5_2236_out0,v$G6_2248_out0 };
assign v$IN_15607_out0 = v$IN_5170_out0;
assign v$IN_15609_out0 = v$IN_5181_out0;
assign v$G1_15782_out0 = ! v$IS$A$LARGER_10444_out0;
assign v$G1_15783_out0 = ! v$IS$A$LARGER_10445_out0;
assign v$_16000_out0 = { v$G11_8202_out0,v$G12_13795_out0 };
assign v$_16001_out0 = { v$G11_8203_out0,v$G12_13796_out0 };
assign v$EXPONENT_16011_out0 = v$SEL18_18251_out0;
assign v$EXPONENT_16012_out0 = v$SEL18_18252_out0;
assign v$_16775_out0 = { v$G9_3441_out0,v$G10_18485_out0 };
assign v$_16776_out0 = { v$G9_3442_out0,v$G10_18486_out0 };
assign v$MUX4_17721_out0 = v$G4_11870_out0 ? v$A_3242_out0 : v$B_17746_out0;
assign v$MUX4_17722_out0 = v$G4_11871_out0 ? v$A_3243_out0 : v$B_17747_out0;
assign v$_18565_out0 = { v$G13_1689_out0,v$G14_1673_out0 };
assign v$_18566_out0 = { v$G13_1690_out0,v$G14_1674_out0 };
assign v$_258_out0 = { v$_18565_out0,v$_3145_out0 };
assign v$_259_out0 = { v$_18566_out0,v$_3146_out0 };
assign v$EXPONENT_1358_out0 = v$SINGLE$PRECISION$EXPONENT_11046_out0;
assign v$EXPONENT_1359_out0 = v$SINGLE$PRECISION$EXPONENT_11047_out0;
assign v$_3706_out0 = { v$_16775_out0,v$_16000_out0 };
assign v$_3707_out0 = { v$_16776_out0,v$_16001_out0 };
assign v$SEL1_8718_out0 = v$IN_15607_out0[23:4];
assign v$SEL1_8729_out0 = v$IN_15609_out0[23:4];
assign v$OP1$MANTISA_9121_out0 = v$MUX3_12800_out0;
assign v$OP1$MANTISA_9122_out0 = v$MUX3_12801_out0;
assign v$SEL1_9465_out0 = v$MUX4_17721_out0[14:10];
assign v$SEL1_9466_out0 = v$MUX4_17722_out0[14:10];
assign v$OP2$MANTISA_9544_out0 = v$MUX9_2458_out0;
assign v$OP2$MANTISA_9545_out0 = v$MUX9_2459_out0;
assign v$_13013_out0 = { v$_14212_out0,v$_9457_out0 };
assign v$_13014_out0 = { v$_14213_out0,v$_9458_out0 };
assign v$SEL1_15409_out0 = v$IN_15607_out0[19:0];
assign v$SEL1_15420_out0 = v$IN_15609_out0[19:0];
assign v$G2_16502_out0 = v$IS$SUB_13067_out0 && v$G1_15782_out0;
assign v$G2_16503_out0 = v$IS$SUB_13068_out0 && v$G1_15783_out0;
assign v$_16886_out0 = { v$_14166_out0,v$_10974_out0 };
assign v$_16887_out0 = { v$_14167_out0,v$_10975_out0 };
assign v$C0_204_out0 = v$_16886_out0;
assign v$C0_205_out0 = v$_16887_out0;
assign v$OP2$MANTISA_2656_out0 = v$OP2$MANTISA_9544_out0;
assign v$OP2$MANTISA_2657_out0 = v$OP2$MANTISA_9545_out0;
assign v$C12_3282_out0 = v$_258_out0;
assign v$C12_3283_out0 = v$_259_out0;
assign v$OP1$MANTISA_3789_out0 = v$OP1$MANTISA_9121_out0;
assign v$OP1$MANTISA_3790_out0 = v$OP1$MANTISA_9122_out0;
assign v$_4268_out0 = { v$C2_126_out0,v$SEL1_15409_out0 };
assign v$_4279_out0 = { v$C2_137_out0,v$SEL1_15420_out0 };
assign v$NEED$SHIFT$OP1_4821_out0 = v$G2_16502_out0;
assign v$NEED$SHIFT$OP1_4822_out0 = v$G2_16503_out0;
assign v$HALF$PRECISION$EXPONENT_6382_out0 = v$SEL1_9465_out0;
assign v$HALF$PRECISION$EXPONENT_6383_out0 = v$SEL1_9466_out0;
assign v$C8_8325_out0 = v$_3706_out0;
assign v$C8_8326_out0 = v$_3707_out0;
assign v$_9003_out0 = { v$SEL1_8718_out0,v$C1_5984_out0 };
assign v$_9014_out0 = { v$SEL1_8729_out0,v$C1_5995_out0 };
assign v$C4_10778_out0 = v$_13013_out0;
assign v$C4_10779_out0 = v$_13014_out0;
assign v$MUX1_2372_out0 = v$LEFT$SHIT_3064_out0 ? v$_4268_out0 : v$_9003_out0;
assign v$MUX1_2383_out0 = v$LEFT$SHIT_3075_out0 ? v$_4279_out0 : v$_9014_out0;
assign v$OP2$MANTISA_3510_out0 = v$OP2$MANTISA_2656_out0;
assign v$OP2$MANTISA_3511_out0 = v$OP2$MANTISA_2657_out0;
assign v$_3687_out0 = { v$C0_204_out0,v$C4_10778_out0 };
assign v$_3688_out0 = { v$C0_205_out0,v$C4_10779_out0 };
assign v$_9043_out0 = { v$C8_8325_out0,v$C12_3282_out0 };
assign v$_9044_out0 = { v$C8_8326_out0,v$C12_3283_out0 };
assign v$OP1$MANTISA_11806_out0 = v$OP1$MANTISA_3789_out0;
assign v$OP1$MANTISA_11807_out0 = v$OP1$MANTISA_3790_out0;
assign v$EXPONENT_16395_out0 = v$HALF$PRECISION$EXPONENT_6382_out0;
assign v$EXPONENT_16396_out0 = v$HALF$PRECISION$EXPONENT_6383_out0;
assign v$IN_13165_out0 = v$OP2$MANTISA_3510_out0;
assign v$IN_13166_out0 = v$OP1$MANTISA_11806_out0;
assign v$IN_13170_out0 = v$OP2$MANTISA_3511_out0;
assign v$IN_13171_out0 = v$OP1$MANTISA_11807_out0;
assign v$MUX2_15238_out0 = v$EN_4755_out0 ? v$MUX1_2372_out0 : v$IN_15607_out0;
assign v$MUX2_15240_out0 = v$EN_4757_out0 ? v$MUX1_2383_out0 : v$IN_15609_out0;
assign v$_16369_out0 = { v$_3687_out0,v$_9043_out0 };
assign v$_16370_out0 = { v$_3688_out0,v$_9044_out0 };
assign v$IN_5149_out0 = v$IN_13165_out0;
assign v$IN_5154_out0 = v$IN_13166_out0;
assign v$IN_5197_out0 = v$IN_13170_out0;
assign v$IN_5202_out0 = v$IN_13171_out0;
assign v$OUT_14924_out0 = v$MUX2_15238_out0;
assign v$OUT_14935_out0 = v$MUX2_15240_out0;
assign v$C_18106_out0 = v$_16369_out0;
assign v$C_18107_out0 = v$_16370_out0;
assign v$IN_3856_out0 = v$IN_5149_out0;
assign v$IN_3857_out0 = v$IN_5154_out0;
assign v$IN_3872_out0 = v$IN_5197_out0;
assign v$IN_3873_out0 = v$IN_5202_out0;
assign v$IN_5168_out0 = v$OUT_14924_out0;
assign v$IN_5179_out0 = v$OUT_14935_out0;
assign v$ANDOUT_7376_out0 = v$C_18106_out0;
assign v$ANDOUT_7377_out0 = v$C_18107_out0;
assign v$MUX3_3880_out0 = v$G6_5944_out0 ? v$ANDOUT_7376_out0 : v$ADDEROUT_3504_out0;
assign v$MUX3_3881_out0 = v$G6_5945_out0 ? v$ANDOUT_7377_out0 : v$ADDEROUT_3505_out0;
assign v$IN_5026_out0 = v$IN_5168_out0;
assign v$IN_5029_out0 = v$IN_5179_out0;
assign v$SEL1_8697_out0 = v$IN_3856_out0[23:1];
assign v$SEL1_8702_out0 = v$IN_3857_out0[23:1];
assign v$SEL1_8745_out0 = v$IN_3872_out0[23:1];
assign v$SEL1_8750_out0 = v$IN_3873_out0[23:1];
assign v$SEL1_15388_out0 = v$IN_3856_out0[22:0];
assign v$SEL1_15393_out0 = v$IN_3857_out0[22:0];
assign v$SEL1_15436_out0 = v$IN_3872_out0[22:0];
assign v$SEL1_15441_out0 = v$IN_3873_out0[22:0];
assign v$_4247_out0 = { v$C2_105_out0,v$SEL1_15388_out0 };
assign v$_4252_out0 = { v$C2_110_out0,v$SEL1_15393_out0 };
assign v$_4295_out0 = { v$C2_153_out0,v$SEL1_15436_out0 };
assign v$_4300_out0 = { v$C2_158_out0,v$SEL1_15441_out0 };
assign v$MUX4_5935_out0 = v$EQ1_2516_out0 ? v$OP2_7579_out0 : v$MUX3_3880_out0;
assign v$MUX4_5936_out0 = v$EQ1_2517_out0 ? v$OP2_7580_out0 : v$MUX3_3881_out0;
assign v$SEL1_8716_out0 = v$IN_5026_out0[23:8];
assign v$SEL1_8727_out0 = v$IN_5029_out0[23:8];
assign v$_8982_out0 = { v$SEL1_8697_out0,v$C1_5963_out0 };
assign v$_8987_out0 = { v$SEL1_8702_out0,v$C1_5968_out0 };
assign v$_9030_out0 = { v$SEL1_8745_out0,v$C1_6011_out0 };
assign v$_9035_out0 = { v$SEL1_8750_out0,v$C1_6016_out0 };
assign v$SEL1_15407_out0 = v$IN_5026_out0[15:0];
assign v$SEL1_15418_out0 = v$IN_5029_out0[15:0];
assign v$MUX1_2351_out0 = v$LEFT$SHIT_3043_out0 ? v$_4247_out0 : v$_8982_out0;
assign v$MUX1_2356_out0 = v$LEFT$SHIT_3048_out0 ? v$_4252_out0 : v$_8987_out0;
assign v$MUX1_2399_out0 = v$LEFT$SHIT_3091_out0 ? v$_4295_out0 : v$_9030_out0;
assign v$MUX1_2404_out0 = v$LEFT$SHIT_3096_out0 ? v$_4300_out0 : v$_9035_out0;
assign v$_4266_out0 = { v$C2_124_out0,v$SEL1_15407_out0 };
assign v$_4277_out0 = { v$C2_135_out0,v$SEL1_15418_out0 };
assign v$_9001_out0 = { v$SEL1_8716_out0,v$C1_5982_out0 };
assign v$_9012_out0 = { v$SEL1_8727_out0,v$C1_5993_out0 };
assign v$ALUOUT_18072_out0 = v$MUX4_5935_out0;
assign v$ALUOUT_18073_out0 = v$MUX4_5936_out0;
assign v$MUX1_2370_out0 = v$LEFT$SHIT_3062_out0 ? v$_4266_out0 : v$_9001_out0;
assign v$MUX1_2381_out0 = v$LEFT$SHIT_3073_out0 ? v$_4277_out0 : v$_9012_out0;
assign v$ALUOUT_6922_out0 = v$ALUOUT_18072_out0;
assign v$ALUOUT_6923_out0 = v$ALUOUT_18073_out0;
assign v$MUX2_18573_out0 = v$EN_5210_out0 ? v$MUX1_2351_out0 : v$IN_3856_out0;
assign v$MUX2_18574_out0 = v$EN_5211_out0 ? v$MUX1_2356_out0 : v$IN_3857_out0;
assign v$MUX2_18586_out0 = v$EN_5223_out0 ? v$MUX1_2399_out0 : v$IN_3872_out0;
assign v$MUX2_18587_out0 = v$EN_5224_out0 ? v$MUX1_2404_out0 : v$IN_3873_out0;
assign v$MUX4_45_out0 = v$IR2$15_7435_out0 ? v$ALUOUT_6922_out0 : v$REGDIN_16498_out0;
assign v$MUX4_46_out0 = v$IR2$15_7436_out0 ? v$ALUOUT_6923_out0 : v$REGDIN_16499_out0;
assign v$MUX2_2500_out0 = v$EN_1339_out0 ? v$MUX1_2370_out0 : v$IN_5026_out0;
assign v$MUX2_2503_out0 = v$EN_1342_out0 ? v$MUX1_2381_out0 : v$IN_5029_out0;
assign v$OUT_14903_out0 = v$MUX2_18573_out0;
assign v$OUT_14908_out0 = v$MUX2_18574_out0;
assign v$OUT_14951_out0 = v$MUX2_18586_out0;
assign v$OUT_14956_out0 = v$MUX2_18587_out0;
assign v$ALUOUT_16542_out0 = v$ALUOUT_6922_out0;
assign v$ALUOUT_16543_out0 = v$ALUOUT_6923_out0;
assign v$IN_5151_out0 = v$OUT_14903_out0;
assign v$IN_5156_out0 = v$OUT_14908_out0;
assign v$IN_5199_out0 = v$OUT_14951_out0;
assign v$IN_5204_out0 = v$OUT_14956_out0;
assign v$ALUOUT_10219_out0 = v$ALUOUT_16542_out0;
assign v$ALUOUT_10220_out0 = v$ALUOUT_16543_out0;
assign v$OUT_14922_out0 = v$MUX2_2500_out0;
assign v$OUT_14933_out0 = v$MUX2_2503_out0;
assign v$IN_5167_out0 = v$OUT_14922_out0;
assign v$IN_5178_out0 = v$OUT_14933_out0;
assign v$_8774_out0 = v$ALUOUT_10219_out0[15:15];
assign v$_8775_out0 = v$ALUOUT_10220_out0[15:15];
assign v$IN_11781_out0 = v$IN_5151_out0;
assign v$IN_11782_out0 = v$IN_5156_out0;
assign v$IN_11790_out0 = v$IN_5199_out0;
assign v$IN_11791_out0 = v$IN_5204_out0;
assign v$EQ1_16270_out0 = v$ALUOUT_10219_out0 == 16'h0;
assign v$EQ1_16271_out0 = v$ALUOUT_10220_out0 == 16'h0;
assign v$IN_5025_out0 = v$IN_5167_out0;
assign v$IN_5028_out0 = v$IN_5178_out0;
assign v$SEL1_8699_out0 = v$IN_11781_out0[23:2];
assign v$SEL1_8704_out0 = v$IN_11782_out0[23:2];
assign v$SEL1_8747_out0 = v$IN_11790_out0[23:2];
assign v$SEL1_8752_out0 = v$IN_11791_out0[23:2];
assign v$G18_13600_out0 = v$_8774_out0 && v$IR2$VALID_13250_out0;
assign v$G18_13601_out0 = v$_8775_out0 && v$IR2$VALID_13251_out0;
assign v$G17_13831_out0 = v$EQ1_16270_out0 && v$IR2$VALID_13250_out0;
assign v$G17_13832_out0 = v$EQ1_16271_out0 && v$IR2$VALID_13251_out0;
assign v$SEL1_15390_out0 = v$IN_11781_out0[21:0];
assign v$SEL1_15395_out0 = v$IN_11782_out0[21:0];
assign v$SEL1_15438_out0 = v$IN_11790_out0[21:0];
assign v$SEL1_15443_out0 = v$IN_11791_out0[21:0];
assign v$MUX3_1428_out0 = v$G18_13600_out0 ? v$G18_13600_out0 : v$REG2_11798_out0;
assign v$MUX3_1429_out0 = v$G18_13601_out0 ? v$G18_13601_out0 : v$REG2_11799_out0;
assign v$_4249_out0 = { v$C2_107_out0,v$SEL1_15390_out0 };
assign v$_4254_out0 = { v$C2_112_out0,v$SEL1_15395_out0 };
assign v$_4297_out0 = { v$C2_155_out0,v$SEL1_15438_out0 };
assign v$_4302_out0 = { v$C2_160_out0,v$SEL1_15443_out0 };
assign v$SEL1_8715_out0 = v$IN_5025_out0[23:16];
assign v$SEL1_8726_out0 = v$IN_5028_out0[23:16];
assign v$_8984_out0 = { v$SEL1_8699_out0,v$C1_5965_out0 };
assign v$_8989_out0 = { v$SEL1_8704_out0,v$C1_5970_out0 };
assign v$_9032_out0 = { v$SEL1_8747_out0,v$C1_6013_out0 };
assign v$_9037_out0 = { v$SEL1_8752_out0,v$C1_6018_out0 };
assign v$MUX4_12637_out0 = v$G17_13831_out0 ? v$G17_13831_out0 : v$REG3_17753_out0;
assign v$MUX4_12638_out0 = v$G17_13832_out0 ? v$G17_13832_out0 : v$REG3_17754_out0;
assign v$SEL1_15406_out0 = v$IN_5025_out0[7:0];
assign v$SEL1_15417_out0 = v$IN_5028_out0[7:0];
assign v$MUX1_2353_out0 = v$LEFT$SHIT_3045_out0 ? v$_4249_out0 : v$_8984_out0;
assign v$MUX1_2358_out0 = v$LEFT$SHIT_3050_out0 ? v$_4254_out0 : v$_8989_out0;
assign v$MUX1_2401_out0 = v$LEFT$SHIT_3093_out0 ? v$_4297_out0 : v$_9032_out0;
assign v$MUX1_2406_out0 = v$LEFT$SHIT_3098_out0 ? v$_4302_out0 : v$_9037_out0;
assign v$EQ_3708_out0 = v$MUX4_12637_out0;
assign v$EQ_3709_out0 = v$MUX4_12638_out0;
assign v$_4265_out0 = { v$C2_123_out0,v$SEL1_15406_out0 };
assign v$_4276_out0 = { v$C2_134_out0,v$SEL1_15417_out0 };
assign v$_9000_out0 = { v$SEL1_8715_out0,v$C1_5981_out0 };
assign v$_9011_out0 = { v$SEL1_8726_out0,v$C1_5992_out0 };
assign v$MI_12128_out0 = v$MUX3_1428_out0;
assign v$MI_12129_out0 = v$MUX3_1429_out0;
assign v$EQ_431_out0 = v$EQ_3708_out0;
assign v$EQ_432_out0 = v$EQ_3709_out0;
assign v$MUX1_2369_out0 = v$LEFT$SHIT_3061_out0 ? v$_4265_out0 : v$_9000_out0;
assign v$MUX1_2380_out0 = v$LEFT$SHIT_3072_out0 ? v$_4276_out0 : v$_9011_out0;
assign v$MUX2_2475_out0 = v$EN_7873_out0 ? v$MUX1_2353_out0 : v$IN_11781_out0;
assign v$MUX2_2476_out0 = v$EN_7874_out0 ? v$MUX1_2358_out0 : v$IN_11782_out0;
assign v$MUX2_2484_out0 = v$EN_7882_out0 ? v$MUX1_2401_out0 : v$IN_11790_out0;
assign v$MUX2_2485_out0 = v$EN_7883_out0 ? v$MUX1_2406_out0 : v$IN_11791_out0;
assign v$MI_6238_out0 = v$MI_12128_out0;
assign v$MI_6239_out0 = v$MI_12129_out0;
assign v$MI_2416_out0 = v$MI_6238_out0;
assign v$MI_2417_out0 = v$MI_6239_out0;
assign v$MUX2_2499_out0 = v$EN_1338_out0 ? v$MUX1_2369_out0 : v$IN_5025_out0;
assign v$MUX2_2502_out0 = v$EN_1341_out0 ? v$MUX1_2380_out0 : v$IN_5028_out0;
assign v$EQ_6151_out0 = v$EQ_431_out0;
assign v$EQ_6152_out0 = v$EQ_432_out0;
assign v$OUT_14905_out0 = v$MUX2_2475_out0;
assign v$OUT_14910_out0 = v$MUX2_2476_out0;
assign v$OUT_14953_out0 = v$MUX2_2484_out0;
assign v$OUT_14958_out0 = v$MUX2_2485_out0;
assign v$EQ_3478_out0 = v$EQ_6151_out0;
assign v$EQ_3479_out0 = v$EQ_6152_out0;
assign v$IN_5150_out0 = v$OUT_14905_out0;
assign v$IN_5155_out0 = v$OUT_14910_out0;
assign v$IN_5198_out0 = v$OUT_14953_out0;
assign v$IN_5203_out0 = v$OUT_14958_out0;
assign v$MI_8450_out0 = v$MI_2416_out0;
assign v$MI_8451_out0 = v$MI_2417_out0;
assign v$OUT_14921_out0 = v$MUX2_2499_out0;
assign v$OUT_14932_out0 = v$MUX2_2502_out0;
assign v$MUX1_11633_out0 = v$G2_17414_out0 ? v$C1_4457_out0 : v$OUT_14921_out0;
assign v$MUX1_11634_out0 = v$G2_17415_out0 ? v$C1_4458_out0 : v$OUT_14932_out0;
assign v$MI_12466_out0 = v$MI_8450_out0;
assign v$MI_12467_out0 = v$MI_8451_out0;
assign v$EQ_13422_out0 = v$EQ_3478_out0;
assign v$EQ_13423_out0 = v$EQ_3479_out0;
assign v$IN_15603_out0 = v$IN_5150_out0;
assign v$IN_15604_out0 = v$IN_5155_out0;
assign v$IN_15612_out0 = v$IN_5198_out0;
assign v$IN_15613_out0 = v$IN_5203_out0;
assign v$SEL1_8698_out0 = v$IN_15603_out0[23:4];
assign v$SEL1_8703_out0 = v$IN_15604_out0[23:4];
assign v$SEL1_8746_out0 = v$IN_15612_out0[23:4];
assign v$SEL1_8751_out0 = v$IN_15613_out0[23:4];
assign v$OUT_10014_out0 = v$MUX1_11633_out0;
assign v$OUT_10015_out0 = v$MUX1_11634_out0;
assign v$MI_11878_out0 = v$MI_12466_out0;
assign v$MI_11879_out0 = v$MI_12467_out0;
assign v$EQ_14576_out0 = v$EQ_13422_out0;
assign v$EQ_14577_out0 = v$EQ_13423_out0;
assign v$SEL1_15389_out0 = v$IN_15603_out0[19:0];
assign v$SEL1_15394_out0 = v$IN_15604_out0[19:0];
assign v$SEL1_15437_out0 = v$IN_15612_out0[19:0];
assign v$SEL1_15442_out0 = v$IN_15613_out0[19:0];
assign v$G20_2594_out0 = v$G22_15342_out0 || v$EQ_14576_out0;
assign v$G20_2595_out0 = v$G22_15343_out0 || v$EQ_14577_out0;
assign v$OP2_4162_out0 = v$OUT_10014_out0;
assign v$OP2_4163_out0 = v$OUT_10015_out0;
assign v$_4248_out0 = { v$C2_106_out0,v$SEL1_15389_out0 };
assign v$_4253_out0 = { v$C2_111_out0,v$SEL1_15394_out0 };
assign v$_4296_out0 = { v$C2_154_out0,v$SEL1_15437_out0 };
assign v$_4301_out0 = { v$C2_159_out0,v$SEL1_15442_out0 };
assign v$_8983_out0 = { v$SEL1_8698_out0,v$C1_5964_out0 };
assign v$_8988_out0 = { v$SEL1_8703_out0,v$C1_5969_out0 };
assign v$_9031_out0 = { v$SEL1_8746_out0,v$C1_6012_out0 };
assign v$_9036_out0 = { v$SEL1_8751_out0,v$C1_6017_out0 };
assign v$G25_12754_out0 = v$JEQ_1675_out0 && v$EQ_14576_out0;
assign v$G25_12755_out0 = v$JEQ_1676_out0 && v$EQ_14577_out0;
assign v$G19_13997_out0 = v$JMI_13149_out0 && v$MI_11878_out0;
assign v$G19_13998_out0 = v$JMI_13150_out0 && v$MI_11879_out0;
assign v$G24_672_out0 = v$JLS_16442_out0 && v$G20_2594_out0;
assign v$G24_673_out0 = v$JLS_16443_out0 && v$G20_2595_out0;
assign v$MUX1_2352_out0 = v$LEFT$SHIT_3044_out0 ? v$_4248_out0 : v$_8983_out0;
assign v$MUX1_2357_out0 = v$LEFT$SHIT_3049_out0 ? v$_4253_out0 : v$_8988_out0;
assign v$MUX1_2400_out0 = v$LEFT$SHIT_3092_out0 ? v$_4296_out0 : v$_9031_out0;
assign v$MUX1_2405_out0 = v$LEFT$SHIT_3097_out0 ? v$_4301_out0 : v$_9036_out0;
assign v$B_8359_out0 = v$OP2_4163_out0;
assign v$B_13561_out0 = v$OP2_4162_out0;
assign v$G21_15312_out0 = v$G19_13997_out0 || v$G25_12754_out0;
assign v$G21_15313_out0 = v$G19_13998_out0 || v$G25_12755_out0;
assign v$B_81_out0 = v$B_13561_out0;
assign v$B_1965_out0 = v$B_8359_out0;
assign v$G15_5478_out0 = v$JMP_4337_out0 || v$G21_15312_out0;
assign v$G15_5479_out0 = v$JMP_4338_out0 || v$G21_15313_out0;
assign v$MUX2_15234_out0 = v$EN_4751_out0 ? v$MUX1_2352_out0 : v$IN_15603_out0;
assign v$MUX2_15235_out0 = v$EN_4752_out0 ? v$MUX1_2357_out0 : v$IN_15604_out0;
assign v$MUX2_15243_out0 = v$EN_4760_out0 ? v$MUX1_2400_out0 : v$IN_15612_out0;
assign v$MUX2_15244_out0 = v$EN_4761_out0 ? v$MUX1_2405_out0 : v$IN_15613_out0;
assign v$SEL7_1223_out0 = v$B_1965_out0[0:0];
assign v$MUX1_2888_out0 = v$START_4238_out0 ? v$B_81_out0 : v$B$SHIFTED_13792_out0;
assign v$OP2_3670_out0 = v$B_1965_out0;
assign v$OP2_6354_out0 = v$B_1965_out0;
assign v$OP2_6356_out0 = v$B_1965_out0;
assign v$OP2_6357_out0 = v$B_1965_out0;
assign v$OP2_6358_out0 = v$B_1965_out0;
assign v$OP2_6359_out0 = v$B_1965_out0;
assign v$OP2_6360_out0 = v$B_1965_out0;
assign v$OP2_6361_out0 = v$B_1965_out0;
assign v$OP2_6362_out0 = v$B_1965_out0;
assign v$OP2_6363_out0 = v$B_1965_out0;
assign v$OP2_6364_out0 = v$B_1965_out0;
assign v$OP2_6365_out0 = v$B_1965_out0;
assign v$MUX4_8103_out0 = v$START_4238_out0 ? v$B_81_out0 : v$B$SHIFTED_13792_out0;
assign v$OUT_14904_out0 = v$MUX2_15234_out0;
assign v$OUT_14909_out0 = v$MUX2_15235_out0;
assign v$OUT_14952_out0 = v$MUX2_15243_out0;
assign v$OUT_14957_out0 = v$MUX2_15244_out0;
assign v$G23_17687_out0 = v$G15_5478_out0 || v$G17_5460_out0;
assign v$G23_17688_out0 = v$G15_5479_out0 || v$G17_5461_out0;
assign v$G16_1314_out0 = v$G23_17687_out0 || v$G24_672_out0;
assign v$G16_1315_out0 = v$G23_17688_out0 || v$G24_673_out0;
assign v$IN_5148_out0 = v$OUT_14904_out0;
assign v$IN_5153_out0 = v$OUT_14909_out0;
assign v$IN_5177_out0 = v$MUX4_8103_out0;
assign v$IN_5196_out0 = v$OUT_14952_out0;
assign v$IN_5201_out0 = v$OUT_14957_out0;
assign v$MUX3_7636_out0 = v$SEL7_1223_out0 ? v$A_14801_out0 : v$C2_7814_out0;
assign v$SEL1_11087_out0 = v$OP2_6354_out0[12:12];
assign v$SEL1_11088_out0 = v$OP2_3670_out0[1:1];
assign v$SEL1_11089_out0 = v$OP2_6356_out0[8:8];
assign v$SEL1_11090_out0 = v$OP2_6357_out0[10:10];
assign v$SEL1_11091_out0 = v$OP2_6358_out0[9:9];
assign v$SEL1_11092_out0 = v$OP2_6359_out0[11:11];
assign v$SEL1_11093_out0 = v$OP2_6360_out0[7:7];
assign v$SEL1_11094_out0 = v$OP2_6361_out0[2:2];
assign v$SEL1_11095_out0 = v$OP2_6362_out0[6:6];
assign v$SEL1_11096_out0 = v$OP2_6363_out0[3:3];
assign v$SEL1_11097_out0 = v$OP2_6364_out0[4:4];
assign v$SEL1_11098_out0 = v$OP2_6365_out0[5:5];
assign v$SEL2_11607_out0 = v$OP2_3670_out0[13:13];
assign v$SEL2_11608_out0 = v$OP2_6356_out0[20:20];
assign v$SEL2_11609_out0 = v$OP2_6357_out0[22:22];
assign v$SEL2_11610_out0 = v$OP2_6358_out0[21:21];
assign v$SEL2_11611_out0 = v$OP2_6359_out0[23:23];
assign v$SEL2_11612_out0 = v$OP2_6360_out0[19:19];
assign v$SEL2_11613_out0 = v$OP2_6361_out0[14:14];
assign v$SEL2_11614_out0 = v$OP2_6362_out0[18:18];
assign v$SEL2_11615_out0 = v$OP2_6363_out0[15:15];
assign v$SEL2_11616_out0 = v$OP2_6364_out0[16:16];
assign v$SEL2_11617_out0 = v$OP2_6365_out0[17:17];
assign v$OP2_12455_out0 = v$MUX1_2888_out0;
assign v$SEL1_1280_out0 = v$OP2_12455_out0[0:0];
assign v$MULTIPLYING$BIT_2849_out0 = v$SEL1_11087_out0;
assign v$IN_3864_out0 = v$IN_5177_out0;
assign v$IN_5019_out0 = v$IN_5148_out0;
assign v$IN_5021_out0 = v$IN_5153_out0;
assign v$IN_5033_out0 = v$IN_5196_out0;
assign v$IN_5035_out0 = v$IN_5201_out0;
assign v$TAKEJUMP_10799_out0 = v$G16_1314_out0;
assign v$TAKEJUMP_10800_out0 = v$G16_1315_out0;
assign v$MUX1_16952_out0 = v$EXEC1_7960_out0 ? v$SEL1_11088_out0 : v$SEL2_11607_out0;
assign v$MUX1_16953_out0 = v$EXEC1_7961_out0 ? v$SEL1_11089_out0 : v$SEL2_11608_out0;
assign v$MUX1_16954_out0 = v$EXEC1_7962_out0 ? v$SEL1_11090_out0 : v$SEL2_11609_out0;
assign v$MUX1_16955_out0 = v$EXEC1_7963_out0 ? v$SEL1_11091_out0 : v$SEL2_11610_out0;
assign v$MUX1_16956_out0 = v$EXEC1_7964_out0 ? v$SEL1_11092_out0 : v$SEL2_11611_out0;
assign v$MUX1_16957_out0 = v$EXEC1_7965_out0 ? v$SEL1_11093_out0 : v$SEL2_11612_out0;
assign v$MUX1_16958_out0 = v$EXEC1_7966_out0 ? v$SEL1_11094_out0 : v$SEL2_11613_out0;
assign v$MUX1_16959_out0 = v$EXEC1_7967_out0 ? v$SEL1_11095_out0 : v$SEL2_11614_out0;
assign v$MUX1_16960_out0 = v$EXEC1_7968_out0 ? v$SEL1_11096_out0 : v$SEL2_11615_out0;
assign v$MUX1_16961_out0 = v$EXEC1_7969_out0 ? v$SEL1_11097_out0 : v$SEL2_11616_out0;
assign v$MUX1_16962_out0 = v$EXEC1_7970_out0 ? v$SEL1_11098_out0 : v$SEL2_11617_out0;
assign v$MUX2_18043_out0 = v$EXEC1_18513_out0 ? v$MUX3_7636_out0 : v$SEL6_5757_out0;
assign v$SEL3_18659_out0 = v$OP2_12455_out0[0:0];
assign v$SEL5_1581_out0 = v$MUX2_18043_out0[0:0];
assign v$MULTIPLYING$BIT_2850_out0 = v$MUX1_16952_out0;
assign v$MULTIPLYING$BIT_2851_out0 = v$MUX1_16953_out0;
assign v$MULTIPLYING$BIT_2852_out0 = v$MUX1_16954_out0;
assign v$MULTIPLYING$BIT_2853_out0 = v$MUX1_16955_out0;
assign v$MULTIPLYING$BIT_2854_out0 = v$MUX1_16956_out0;
assign v$MULTIPLYING$BIT_2855_out0 = v$MUX1_16957_out0;
assign v$MULTIPLYING$BIT_2856_out0 = v$MUX1_16958_out0;
assign v$MULTIPLYING$BIT_2857_out0 = v$MUX1_16959_out0;
assign v$MULTIPLYING$BIT_2858_out0 = v$MUX1_16960_out0;
assign v$MULTIPLYING$BIT_2859_out0 = v$MUX1_16961_out0;
assign v$MULTIPLYING$BIT_2860_out0 = v$MUX1_16962_out0;
assign v$MUX1_8338_out0 = v$MULTIPLYING$BIT_2849_out0 ? v$OP2_10374_out0 : v$C5_3961_out0;
assign v$SEL1_8696_out0 = v$IN_5019_out0[23:8];
assign v$SEL1_8701_out0 = v$IN_5021_out0[23:8];
assign v$SEL1_8725_out0 = v$IN_3864_out0[23:1];
assign v$SEL1_8744_out0 = v$IN_5033_out0[23:8];
assign v$SEL1_8749_out0 = v$IN_5035_out0[23:8];
assign v$MUX5_10310_out0 = v$SEL3_18659_out0 ? v$_1158_out0 : v$C4_17973_out0;
assign v$MUX2_12458_out0 = v$SEL1_1280_out0 ? v$A_14255_out0 : v$C3_18437_out0;
assign v$G26_13641_out0 = v$G29_7851_out0 || v$TAKEJUMP_10799_out0;
assign v$G26_13642_out0 = v$G29_7852_out0 || v$TAKEJUMP_10800_out0;
assign v$OP1_14186_out0 = v$MUX2_18043_out0;
assign v$SEL1_15387_out0 = v$IN_5019_out0[15:0];
assign v$SEL1_15392_out0 = v$IN_5021_out0[15:0];
assign v$SEL1_15416_out0 = v$IN_3864_out0[22:0];
assign v$SEL1_15435_out0 = v$IN_5033_out0[15:0];
assign v$SEL1_15440_out0 = v$IN_5035_out0[15:0];
assign v$OP1_3380_out0 = v$OP1_14186_out0;
assign v$_4246_out0 = { v$C2_104_out0,v$SEL1_15387_out0 };
assign v$_4251_out0 = { v$C2_109_out0,v$SEL1_15392_out0 };
assign v$_4275_out0 = { v$C2_133_out0,v$SEL1_15416_out0 };
assign v$_4294_out0 = { v$C2_152_out0,v$SEL1_15435_out0 };
assign v$_4299_out0 = { v$C2_157_out0,v$SEL1_15440_out0 };
assign v$MUX1_8339_out0 = v$MULTIPLYING$BIT_2850_out0 ? v$OP2_10375_out0 : v$C5_3962_out0;
assign v$MUX1_8340_out0 = v$MULTIPLYING$BIT_2851_out0 ? v$OP2_10376_out0 : v$C5_3963_out0;
assign v$MUX1_8341_out0 = v$MULTIPLYING$BIT_2852_out0 ? v$OP2_10377_out0 : v$C5_3964_out0;
assign v$MUX1_8342_out0 = v$MULTIPLYING$BIT_2853_out0 ? v$OP2_10378_out0 : v$C5_3965_out0;
assign v$MUX1_8343_out0 = v$MULTIPLYING$BIT_2854_out0 ? v$OP2_10379_out0 : v$C5_3966_out0;
assign v$MUX1_8344_out0 = v$MULTIPLYING$BIT_2855_out0 ? v$OP2_10380_out0 : v$C5_3967_out0;
assign v$MUX1_8345_out0 = v$MULTIPLYING$BIT_2856_out0 ? v$OP2_10381_out0 : v$C5_3968_out0;
assign v$MUX1_8346_out0 = v$MULTIPLYING$BIT_2857_out0 ? v$OP2_10382_out0 : v$C5_3969_out0;
assign v$MUX1_8347_out0 = v$MULTIPLYING$BIT_2858_out0 ? v$OP2_10383_out0 : v$C5_3970_out0;
assign v$MUX1_8348_out0 = v$MULTIPLYING$BIT_2859_out0 ? v$OP2_10384_out0 : v$C5_3971_out0;
assign v$MUX1_8349_out0 = v$MULTIPLYING$BIT_2860_out0 ? v$OP2_10385_out0 : v$C5_3972_out0;
assign v$B2_8417_out0 = v$MUX2_12458_out0;
assign v$_8981_out0 = { v$SEL1_8696_out0,v$C1_5962_out0 };
assign v$_8986_out0 = { v$SEL1_8701_out0,v$C1_5967_out0 };
assign v$_9010_out0 = { v$SEL1_8725_out0,v$C1_5991_out0 };
assign v$_9029_out0 = { v$SEL1_8744_out0,v$C1_6010_out0 };
assign v$_9034_out0 = { v$SEL1_8749_out0,v$C1_6015_out0 };
assign v$MUX8_12286_out0 = v$G26_13641_out0 ? v$MUX5_16988_out0 : v$PCINTERRUPT_17807_out0;
assign v$MUX8_12287_out0 = v$G26_13642_out0 ? v$MUX5_16989_out0 : v$PCINTERRUPT_17808_out0;
assign v$SUM$0_12330_out0 = v$SEL5_1581_out0;
assign v$MUX3_17902_out0 = v$START_4238_out0 ? v$MUX5_10310_out0 : v$RESULT_5062_out0;
assign v$MUX1_2350_out0 = v$LEFT$SHIT_3042_out0 ? v$_4246_out0 : v$_8981_out0;
assign v$MUX1_2355_out0 = v$LEFT$SHIT_3047_out0 ? v$_4251_out0 : v$_8986_out0;
assign v$MUX1_2379_out0 = v$LEFT$SHIT_3071_out0 ? v$_4275_out0 : v$_9010_out0;
assign v$MUX1_2398_out0 = v$LEFT$SHIT_3090_out0 ? v$_4294_out0 : v$_9029_out0;
assign v$MUX1_2403_out0 = v$LEFT$SHIT_3095_out0 ? v$_4299_out0 : v$_9034_out0;
assign v$MUX2_3722_out0 = v$ININTERRUPT_1133_out0 ? v$MUX8_12286_out0 : v$PCNORMAL_12768_out0;
assign v$MUX2_3723_out0 = v$ININTERRUPT_1134_out0 ? v$MUX8_12287_out0 : v$PCNORMAL_12769_out0;
assign v$_3987_out0 = v$B2_8417_out0[11:0];
assign v$_3987_out1 = v$B2_8417_out0[23:12];
assign v$A1_13597_out0 = v$MUX3_17902_out0;
assign v$SEL8_17652_out0 = v$OP1_3380_out0[23:1];
assign v$_1220_out0 = v$_3987_out1[5:0];
assign v$_1220_out1 = v$_3987_out1[11:6];
assign v$_1525_out0 = v$_3987_out0[5:0];
assign v$_1525_out1 = v$_3987_out0[11:6];
assign v$MUX4_1574_out0 = v$TAKEJUMP_10799_out0 ? v$N_18295_out0 : v$MUX2_3722_out0;
assign v$MUX4_1575_out0 = v$TAKEJUMP_10800_out0 ? v$N_18296_out0 : v$MUX2_3723_out0;
assign v$MUX2_2493_out0 = v$EN_1332_out0 ? v$MUX1_2350_out0 : v$IN_5019_out0;
assign v$MUX2_2495_out0 = v$EN_1334_out0 ? v$MUX1_2355_out0 : v$IN_5021_out0;
assign v$MUX2_2507_out0 = v$EN_1346_out0 ? v$MUX1_2398_out0 : v$IN_5033_out0;
assign v$MUX2_2509_out0 = v$EN_1348_out0 ? v$MUX1_2403_out0 : v$IN_5035_out0;
assign v$_7541_out0 = v$A1_13597_out0[11:0];
assign v$_7541_out1 = v$A1_13597_out0[23:12];
assign v$MUX2_14829_out0 = v$EN_3877_out0 ? v$MUX1_2379_out0 : v$IN_3864_out0;
assign v$_17994_out0 = { v$SEL8_17652_out0,v$CIN_16813_out0 };
assign v$PC_3147_out0 = v$MUX4_1574_out0;
assign v$PC_3148_out0 = v$MUX4_1575_out0;
assign v$_9935_out0 = v$_1220_out1[2:0];
assign v$_9935_out1 = v$_1220_out1[5:3];
assign v$_12989_out0 = v$_1525_out1[2:0];
assign v$_12989_out1 = v$_1525_out1[5:3];
assign v$_13743_out0 = v$_1525_out0[2:0];
assign v$_13743_out1 = v$_1525_out0[5:3];
assign v$OUT_14902_out0 = v$MUX2_2493_out0;
assign v$OUT_14907_out0 = v$MUX2_2495_out0;
assign v$OUT_14931_out0 = v$MUX2_14829_out0;
assign v$OUT_14950_out0 = v$MUX2_2507_out0;
assign v$OUT_14955_out0 = v$MUX2_2509_out0;
assign {v$A1_15215_out1,v$A1_15215_out0 } = v$_17994_out0 + v$MUX1_8339_out0 + v$C6_11351_out0;
assign v$_16113_out0 = v$_7541_out0[5:0];
assign v$_16113_out1 = v$_7541_out0[11:6];
assign v$_17030_out0 = v$_7541_out1[5:0];
assign v$_17030_out1 = v$_7541_out1[11:6];
assign v$_17734_out0 = v$_1220_out0[2:0];
assign v$_17734_out1 = v$_1220_out0[5:3];
assign v$NEXTINSTRUCTIONADDRESS_18408_out0 = v$MUX4_1574_out0;
assign v$NEXTINSTRUCTIONADDRESS_18409_out0 = v$MUX4_1575_out0;
assign v$_1865_out0 = v$_17030_out1[2:0];
assign v$_1865_out1 = v$_17030_out1[5:3];
assign v$_2924_out0 = v$_13743_out0[0:0];
assign v$_2924_out1 = v$_13743_out0[2:2];
assign v$IN_5147_out0 = v$OUT_14902_out0;
assign v$IN_5152_out0 = v$OUT_14907_out0;
assign v$IN_5195_out0 = v$OUT_14950_out0;
assign v$IN_5200_out0 = v$OUT_14955_out0;
assign v$PCNEXT_6654_out0 = v$NEXTINSTRUCTIONADDRESS_18408_out0;
assign v$PCNEXT_6655_out0 = v$NEXTINSTRUCTIONADDRESS_18409_out0;
assign v$_7770_out0 = v$_17734_out0[0:0];
assign v$_7770_out1 = v$_17734_out0[2:2];
assign v$COUT_8112_out0 = v$A1_15215_out1;
assign v$_9064_out0 = v$_9935_out1[0:0];
assign v$_9064_out1 = v$_9935_out1[2:2];
assign v$_10050_out0 = v$_17030_out0[2:0];
assign v$_10050_out1 = v$_17030_out0[5:3];
assign v$_10774_out0 = v$_12989_out1[0:0];
assign v$_10774_out1 = v$_12989_out1[2:2];
assign v$_13772_out0 = v$_16113_out0[2:0];
assign v$_13772_out1 = v$_16113_out0[5:3];
assign {v$A1_14820_out1,v$A1_14820_out0 } = v$PC_3147_out0 + v$C1_15940_out0 + v$EN_9080_out0;
assign {v$A1_14821_out1,v$A1_14821_out0 } = v$PC_3148_out0 + v$C1_15941_out0 + v$EN_9081_out0;
assign v$_15150_out0 = v$_9935_out0[0:0];
assign v$_15150_out1 = v$_9935_out0[2:2];
assign v$SUM_15167_out0 = v$A1_15215_out0;
assign v$_16267_out0 = v$_17734_out1[0:0];
assign v$_16267_out1 = v$_17734_out1[2:2];
assign v$_16742_out0 = v$_13743_out1[0:0];
assign v$_16742_out1 = v$_13743_out1[2:2];
assign v$_18190_out0 = v$_12989_out0[0:0];
assign v$_18190_out1 = v$_12989_out0[2:2];
assign v$_18422_out0 = v$_16113_out1[2:0];
assign v$_18422_out1 = v$_16113_out1[5:3];
assign v$_1304_out0 = v$_18422_out0[0:0];
assign v$_1304_out1 = v$_18422_out0[2:2];
assign v$_1355_out0 = v$_13772_out1[0:0];
assign v$_1355_out1 = v$_13772_out1[2:2];
assign v$_1856_out0 = v$_1865_out1[0:0];
assign v$_1856_out1 = v$_1865_out1[2:2];
assign v$PC$NEXT0_1935_out0 = v$PCNEXT_6654_out0;
assign v$B12_1952_out0 = v$_7770_out0;
assign v$B0_3202_out0 = v$_2924_out0;
assign v$SUM_3467_out0 = v$SUM_15167_out0;
assign v$PC$NEXT1_3497_out0 = v$PCNEXT_6655_out0;
assign v$B9_4067_out0 = v$_10774_out0;
assign v$IN_5018_out0 = v$IN_5147_out0;
assign v$IN_5020_out0 = v$IN_5152_out0;
assign v$IN_5032_out0 = v$IN_5195_out0;
assign v$IN_5034_out0 = v$IN_5200_out0;
assign v$IGNORE_5408_out0 = v$A1_14820_out1;
assign v$IGNORE_5409_out0 = v$A1_14821_out1;
assign v$_6900_out0 = v$_18190_out1[0:0];
assign v$_6900_out1 = v$_18190_out1[1:1];
assign v$_6979_out0 = v$_16742_out1[0:0];
assign v$_6979_out1 = v$_16742_out1[1:1];
assign v$_7069_out0 = v$_13772_out0[0:0];
assign v$_7069_out1 = v$_13772_out0[2:2];
assign v$_9383_out0 = v$_9064_out1[0:0];
assign v$_9383_out1 = v$_9064_out1[1:1];
assign v$B3_9473_out0 = v$_16742_out0;
assign v$_9499_out0 = v$_10774_out1[0:0];
assign v$_9499_out1 = v$_10774_out1[1:1];
assign v$B15_10023_out0 = v$_16267_out0;
assign v$_10448_out0 = v$_10050_out0[0:0];
assign v$_10448_out1 = v$_10050_out0[2:2];
assign v$COUT_10729_out0 = v$COUT_8112_out0;
assign v$B18_10869_out0 = v$_15150_out0;
assign v$_10912_out0 = v$_18422_out1[0:0];
assign v$_10912_out1 = v$_18422_out1[2:2];
assign v$_11024_out0 = v$_2924_out1[0:0];
assign v$_11024_out1 = v$_2924_out1[1:1];
assign v$_11101_out0 = v$_1865_out0[0:0];
assign v$_11101_out1 = v$_1865_out0[2:2];
assign v$_13182_out0 = v$_16267_out1[0:0];
assign v$_13182_out1 = v$_16267_out1[1:1];
assign v$B6_13300_out0 = v$_18190_out0;
assign v$SUM_13667_out0 = v$A1_14820_out0;
assign v$SUM_13668_out0 = v$A1_14821_out0;
assign v$_16132_out0 = v$_10050_out1[0:0];
assign v$_16132_out1 = v$_10050_out1[2:2];
assign v$_16591_out0 = v$_15150_out1[0:0];
assign v$_16591_out1 = v$_15150_out1[1:1];
assign v$_17327_out0 = v$_7770_out1[0:0];
assign v$_17327_out1 = v$_7770_out1[1:1];
assign v$B21_18084_out0 = v$_9064_out0;
assign v$A6_310_out0 = v$_1304_out0;
assign v$B23_1285_out0 = v$_9383_out1;
assign v$A21_2600_out0 = v$_1856_out0;
assign v$B_2744_out0 = v$B6_13300_out0;
assign v$B_2745_out0 = v$B3_9473_out0;
assign v$B_2746_out0 = v$B21_18084_out0;
assign v$B_2747_out0 = v$B9_4067_out0;
assign v$B_2748_out0 = v$B15_10023_out0;
assign v$B_2752_out0 = v$B12_1952_out0;
assign v$B_2756_out0 = v$B0_3202_out0;
assign v$B_2761_out0 = v$B18_10869_out0;
assign v$B2_3115_out0 = v$_11024_out1;
assign v$A12_3140_out0 = v$_10448_out0;
assign v$A9_3437_out0 = v$_10912_out0;
assign v$SEL1_3515_out0 = v$SUM_3467_out0[0:0];
assign v$CIN_3893_out0 = v$COUT_10729_out0;
assign v$B20_3945_out0 = v$_16591_out1;
assign v$B14_4004_out0 = v$_17327_out1;
assign v$A0_4310_out0 = v$_7069_out0;
assign v$_5950_out0 = v$_16132_out1[0:0];
assign v$_5950_out1 = v$_16132_out1[1:1];
assign v$_7360_out0 = v$_1355_out1[0:0];
assign v$_7360_out1 = v$_1355_out1[1:1];
assign v$B1_8125_out0 = v$_11024_out0;
assign v$B13_8677_out0 = v$_17327_out0;
assign v$SEL1_8695_out0 = v$IN_5018_out0[23:16];
assign v$SEL1_8700_out0 = v$IN_5020_out0[23:16];
assign v$SEL1_8743_out0 = v$IN_5032_out0[23:16];
assign v$SEL1_8748_out0 = v$IN_5034_out0[23:16];
assign v$B11_9118_out0 = v$_9499_out1;
assign v$B10_9879_out0 = v$_9499_out0;
assign v$_10286_out0 = v$_1856_out1[0:0];
assign v$_10286_out1 = v$_1856_out1[1:1];
assign v$B22_10807_out0 = v$_9383_out0;
assign v$_11620_out0 = v$_7069_out1[0:0];
assign v$_11620_out1 = v$_7069_out1[1:1];
assign v$B8_13140_out0 = v$_6900_out1;
assign v$OP1_14192_out0 = v$SUM_3467_out0;
assign v$A3_14609_out0 = v$_1355_out0;
assign v$B4_14665_out0 = v$_6979_out0;
assign v$ADDRESS_15194_out0 = v$PC$NEXT0_1935_out0;
assign v$ADDRESS_15195_out0 = v$PC$NEXT1_3497_out0;
assign v$SEL1_15386_out0 = v$IN_5018_out0[7:0];
assign v$SEL1_15391_out0 = v$IN_5020_out0[7:0];
assign v$SEL1_15434_out0 = v$IN_5032_out0[7:0];
assign v$SEL1_15439_out0 = v$IN_5034_out0[7:0];
assign v$B17_15537_out0 = v$_13182_out1;
assign v$_15743_out0 = v$_1304_out1[0:0];
assign v$_15743_out1 = v$_1304_out1[1:1];
assign v$_16184_out0 = v$_10448_out1[0:0];
assign v$_16184_out1 = v$_10448_out1[1:1];
assign v$B16_16416_out0 = v$_13182_out0;
assign v$_16706_out0 = v$_11101_out1[0:0];
assign v$_16706_out1 = v$_11101_out1[1:1];
assign v$B19_16791_out0 = v$_16591_out0;
assign v$B7_17042_out0 = v$_6900_out0;
assign v$A15_17320_out0 = v$_16132_out0;
assign v$A18_17697_out0 = v$_11101_out0;
assign v$_17757_out0 = v$_10912_out1[0:0];
assign v$_17757_out1 = v$_10912_out1[1:1];
assign v$B5_18376_out0 = v$_6979_out1;
assign v$A14_678_out0 = v$_16184_out1;
assign v$A19_1215_out0 = v$_16706_out0;
assign v$A10_1550_out0 = v$_17757_out0;
assign v$A1_1712_out0 = v$_11620_out0;
assign v$B_2749_out0 = v$B7_17042_out0;
assign v$B_2750_out0 = v$B1_8125_out0;
assign v$B_2751_out0 = v$B14_4004_out0;
assign v$B_2753_out0 = v$B8_13140_out0;
assign v$B_2754_out0 = v$B17_15537_out0;
assign v$B_2755_out0 = v$B23_1285_out0;
assign v$B_2757_out0 = v$B13_8677_out0;
assign v$B_2758_out0 = v$B4_14665_out0;
assign v$B_2759_out0 = v$B19_16791_out0;
assign v$B_2760_out0 = v$B22_10807_out0;
assign v$B_2762_out0 = v$B10_9879_out0;
assign v$B_2763_out0 = v$B20_3945_out0;
assign v$B_2764_out0 = v$B2_3115_out0;
assign v$B_2765_out0 = v$B11_9118_out0;
assign v$B_2766_out0 = v$B5_18376_out0;
assign v$B_2767_out0 = v$B16_16416_out0;
assign v$OP1_3386_out0 = v$OP1_14192_out0;
assign v$_4245_out0 = { v$C2_103_out0,v$SEL1_15386_out0 };
assign v$_4250_out0 = { v$C2_108_out0,v$SEL1_15391_out0 };
assign v$_4293_out0 = { v$C2_151_out0,v$SEL1_15434_out0 };
assign v$_4298_out0 = { v$C2_156_out0,v$SEL1_15439_out0 };
assign v$A22_4426_out0 = v$_10286_out0;
assign v$A20_4438_out0 = v$_16706_out1;
assign v$A23_5065_out0 = v$_10286_out1;
assign v$A5_6667_out0 = v$_7360_out1;
assign v$A_7149_out0 = v$A6_310_out0;
assign v$A_7150_out0 = v$A3_14609_out0;
assign v$A_7151_out0 = v$A21_2600_out0;
assign v$A_7152_out0 = v$A9_3437_out0;
assign v$A_7153_out0 = v$A15_17320_out0;
assign v$A_7157_out0 = v$A12_3140_out0;
assign v$A_7161_out0 = v$A0_4310_out0;
assign v$A_7166_out0 = v$A18_17697_out0;
assign v$_8980_out0 = { v$SEL1_8695_out0,v$C1_5961_out0 };
assign v$_8985_out0 = { v$SEL1_8700_out0,v$C1_5966_out0 };
assign v$_9028_out0 = { v$SEL1_8743_out0,v$C1_6009_out0 };
assign v$_9033_out0 = { v$SEL1_8748_out0,v$C1_6014_out0 };
assign v$A11_9964_out0 = v$_17757_out1;
assign v$SUM$1_10360_out0 = v$SEL1_3515_out0;
assign {v$A1A_11662_out1,v$A1A_11662_out0 } = v$A0_4310_out0 + v$B0_3202_out0 + v$C1_4466_out0;
assign v$A16_13616_out0 = v$_5950_out0;
assign v$A13_13864_out0 = v$_16184_out0;
assign v$A7_15309_out0 = v$_15743_out0;
assign v$A17_16724_out0 = v$_5950_out1;
assign v$CIN_16819_out0 = v$CIN_3893_out0;
assign v$A4_17500_out0 = v$_7360_out0;
assign v$A8_18092_out0 = v$_15743_out1;
assign v$A2_18268_out0 = v$_11620_out1;
assign v$MUX1_2349_out0 = v$LEFT$SHIT_3041_out0 ? v$_4245_out0 : v$_8980_out0;
assign v$MUX1_2354_out0 = v$LEFT$SHIT_3046_out0 ? v$_4250_out0 : v$_8985_out0;
assign v$MUX1_2397_out0 = v$LEFT$SHIT_3089_out0 ? v$_4293_out0 : v$_9028_out0;
assign v$MUX1_2402_out0 = v$LEFT$SHIT_3094_out0 ? v$_4298_out0 : v$_9033_out0;
assign v$G2_5309_out0 = ((v$A_7149_out0 && !v$B_2744_out0) || (!v$A_7149_out0) && v$B_2744_out0);
assign v$G2_5310_out0 = ((v$A_7150_out0 && !v$B_2745_out0) || (!v$A_7150_out0) && v$B_2745_out0);
assign v$G2_5311_out0 = ((v$A_7151_out0 && !v$B_2746_out0) || (!v$A_7151_out0) && v$B_2746_out0);
assign v$G2_5312_out0 = ((v$A_7152_out0 && !v$B_2747_out0) || (!v$A_7152_out0) && v$B_2747_out0);
assign v$G2_5313_out0 = ((v$A_7153_out0 && !v$B_2748_out0) || (!v$A_7153_out0) && v$B_2748_out0);
assign v$G2_5317_out0 = ((v$A_7157_out0 && !v$B_2752_out0) || (!v$A_7157_out0) && v$B_2752_out0);
assign v$G2_5321_out0 = ((v$A_7161_out0 && !v$B_2756_out0) || (!v$A_7161_out0) && v$B_2756_out0);
assign v$G2_5326_out0 = ((v$A_7166_out0 && !v$B_2761_out0) || (!v$A_7166_out0) && v$B_2761_out0);
assign v$A_7154_out0 = v$A7_15309_out0;
assign v$A_7155_out0 = v$A1_1712_out0;
assign v$A_7156_out0 = v$A14_678_out0;
assign v$A_7158_out0 = v$A8_18092_out0;
assign v$A_7159_out0 = v$A17_16724_out0;
assign v$A_7160_out0 = v$A23_5065_out0;
assign v$A_7162_out0 = v$A13_13864_out0;
assign v$A_7163_out0 = v$A4_17500_out0;
assign v$A_7164_out0 = v$A19_1215_out0;
assign v$A_7165_out0 = v$A22_4426_out0;
assign v$A_7167_out0 = v$A10_1550_out0;
assign v$A_7168_out0 = v$A20_4438_out0;
assign v$A_7169_out0 = v$A2_18268_out0;
assign v$A_7170_out0 = v$A11_9964_out0;
assign v$A_7171_out0 = v$A5_6667_out0;
assign v$A_7172_out0 = v$A16_13616_out0;
assign v$G1_12383_out0 = v$A_7149_out0 && v$B_2744_out0;
assign v$G1_12384_out0 = v$A_7150_out0 && v$B_2745_out0;
assign v$G1_12385_out0 = v$A_7151_out0 && v$B_2746_out0;
assign v$G1_12386_out0 = v$A_7152_out0 && v$B_2747_out0;
assign v$G1_12387_out0 = v$A_7153_out0 && v$B_2748_out0;
assign v$G1_12391_out0 = v$A_7157_out0 && v$B_2752_out0;
assign v$G1_12395_out0 = v$A_7161_out0 && v$B_2756_out0;
assign v$G1_12400_out0 = v$A_7166_out0 && v$B_2761_out0;
assign v$SEL8_17658_out0 = v$OP1_3386_out0[23:1];
assign v$END_18274_out0 = v$A1A_11662_out1;
assign v$MUX2_2492_out0 = v$EN_1331_out0 ? v$MUX1_2349_out0 : v$IN_5018_out0;
assign v$MUX2_2494_out0 = v$EN_1333_out0 ? v$MUX1_2354_out0 : v$IN_5020_out0;
assign v$MUX2_2506_out0 = v$EN_1345_out0 ? v$MUX1_2397_out0 : v$IN_5032_out0;
assign v$MUX2_2508_out0 = v$EN_1347_out0 ? v$MUX1_2402_out0 : v$IN_5034_out0;
assign v$G2_5314_out0 = ((v$A_7154_out0 && !v$B_2749_out0) || (!v$A_7154_out0) && v$B_2749_out0);
assign v$G2_5315_out0 = ((v$A_7155_out0 && !v$B_2750_out0) || (!v$A_7155_out0) && v$B_2750_out0);
assign v$G2_5316_out0 = ((v$A_7156_out0 && !v$B_2751_out0) || (!v$A_7156_out0) && v$B_2751_out0);
assign v$G2_5318_out0 = ((v$A_7158_out0 && !v$B_2753_out0) || (!v$A_7158_out0) && v$B_2753_out0);
assign v$G2_5319_out0 = ((v$A_7159_out0 && !v$B_2754_out0) || (!v$A_7159_out0) && v$B_2754_out0);
assign v$G2_5320_out0 = ((v$A_7160_out0 && !v$B_2755_out0) || (!v$A_7160_out0) && v$B_2755_out0);
assign v$G2_5322_out0 = ((v$A_7162_out0 && !v$B_2757_out0) || (!v$A_7162_out0) && v$B_2757_out0);
assign v$G2_5323_out0 = ((v$A_7163_out0 && !v$B_2758_out0) || (!v$A_7163_out0) && v$B_2758_out0);
assign v$G2_5324_out0 = ((v$A_7164_out0 && !v$B_2759_out0) || (!v$A_7164_out0) && v$B_2759_out0);
assign v$G2_5325_out0 = ((v$A_7165_out0 && !v$B_2760_out0) || (!v$A_7165_out0) && v$B_2760_out0);
assign v$G2_5327_out0 = ((v$A_7167_out0 && !v$B_2762_out0) || (!v$A_7167_out0) && v$B_2762_out0);
assign v$G2_5328_out0 = ((v$A_7168_out0 && !v$B_2763_out0) || (!v$A_7168_out0) && v$B_2763_out0);
assign v$G2_5329_out0 = ((v$A_7169_out0 && !v$B_2764_out0) || (!v$A_7169_out0) && v$B_2764_out0);
assign v$G2_5330_out0 = ((v$A_7170_out0 && !v$B_2765_out0) || (!v$A_7170_out0) && v$B_2765_out0);
assign v$G2_5331_out0 = ((v$A_7171_out0 && !v$B_2766_out0) || (!v$A_7171_out0) && v$B_2766_out0);
assign v$G2_5332_out0 = ((v$A_7172_out0 && !v$B_2767_out0) || (!v$A_7172_out0) && v$B_2767_out0);
assign v$G_10103_out0 = v$G1_12383_out0;
assign v$G_10104_out0 = v$G1_12384_out0;
assign v$G_10105_out0 = v$G1_12385_out0;
assign v$G_10106_out0 = v$G1_12386_out0;
assign v$G_10107_out0 = v$G1_12387_out0;
assign v$G_10111_out0 = v$G1_12391_out0;
assign v$G_10115_out0 = v$G1_12395_out0;
assign v$G_10120_out0 = v$G1_12400_out0;
assign v$G1_12388_out0 = v$A_7154_out0 && v$B_2749_out0;
assign v$G1_12389_out0 = v$A_7155_out0 && v$B_2750_out0;
assign v$G1_12390_out0 = v$A_7156_out0 && v$B_2751_out0;
assign v$G1_12392_out0 = v$A_7158_out0 && v$B_2753_out0;
assign v$G1_12393_out0 = v$A_7159_out0 && v$B_2754_out0;
assign v$G1_12394_out0 = v$A_7160_out0 && v$B_2755_out0;
assign v$G1_12396_out0 = v$A_7162_out0 && v$B_2757_out0;
assign v$G1_12397_out0 = v$A_7163_out0 && v$B_2758_out0;
assign v$G1_12398_out0 = v$A_7164_out0 && v$B_2759_out0;
assign v$G1_12399_out0 = v$A_7165_out0 && v$B_2760_out0;
assign v$G1_12401_out0 = v$A_7167_out0 && v$B_2762_out0;
assign v$G1_12402_out0 = v$A_7168_out0 && v$B_2763_out0;
assign v$G1_12403_out0 = v$A_7169_out0 && v$B_2764_out0;
assign v$G1_12404_out0 = v$A_7170_out0 && v$B_2765_out0;
assign v$G1_12405_out0 = v$A_7171_out0 && v$B_2766_out0;
assign v$G1_12406_out0 = v$A_7172_out0 && v$B_2767_out0;
assign v$P_13916_out0 = v$G2_5309_out0;
assign v$P_13917_out0 = v$G2_5310_out0;
assign v$P_13918_out0 = v$G2_5311_out0;
assign v$P_13919_out0 = v$G2_5312_out0;
assign v$P_13920_out0 = v$G2_5313_out0;
assign v$P_13924_out0 = v$G2_5317_out0;
assign v$P_13928_out0 = v$G2_5321_out0;
assign v$P_13933_out0 = v$G2_5326_out0;
assign v$_18000_out0 = { v$SEL8_17658_out0,v$CIN_16819_out0 };
assign v$P12_237_out0 = v$P_13924_out0;
assign v$P21_4771_out0 = v$P_13918_out0;
assign v$P0_4812_out0 = v$P_13928_out0;
assign v$P15_6906_out0 = v$P_13920_out0;
assign v$G12_7044_out0 = v$G_10111_out0;
assign v$P6_8106_out0 = v$P_13916_out0;
assign v$G9_8927_out0 = v$G_10106_out0;
assign v$G_10108_out0 = v$G1_12388_out0;
assign v$G_10109_out0 = v$G1_12389_out0;
assign v$G_10110_out0 = v$G1_12390_out0;
assign v$G_10112_out0 = v$G1_12392_out0;
assign v$G_10113_out0 = v$G1_12393_out0;
assign v$G_10114_out0 = v$G1_12394_out0;
assign v$G_10116_out0 = v$G1_12396_out0;
assign v$G_10117_out0 = v$G1_12397_out0;
assign v$G_10118_out0 = v$G1_12398_out0;
assign v$G_10119_out0 = v$G1_12399_out0;
assign v$G_10121_out0 = v$G1_12401_out0;
assign v$G_10122_out0 = v$G1_12402_out0;
assign v$G_10123_out0 = v$G1_12403_out0;
assign v$G_10124_out0 = v$G1_12404_out0;
assign v$G_10125_out0 = v$G1_12405_out0;
assign v$G_10126_out0 = v$G1_12406_out0;
assign v$G15_11032_out0 = v$G_10107_out0;
assign v$G3_11106_out0 = v$G_10104_out0;
assign v$P18_11724_out0 = v$P_13933_out0;
assign v$G18_12940_out0 = v$G_10120_out0;
assign v$P_13921_out0 = v$G2_5314_out0;
assign v$P_13922_out0 = v$G2_5315_out0;
assign v$P_13923_out0 = v$G2_5316_out0;
assign v$P_13925_out0 = v$G2_5318_out0;
assign v$P_13926_out0 = v$G2_5319_out0;
assign v$P_13927_out0 = v$G2_5320_out0;
assign v$P_13929_out0 = v$G2_5322_out0;
assign v$P_13930_out0 = v$G2_5323_out0;
assign v$P_13931_out0 = v$G2_5324_out0;
assign v$P_13932_out0 = v$G2_5325_out0;
assign v$P_13934_out0 = v$G2_5327_out0;
assign v$P_13935_out0 = v$G2_5328_out0;
assign v$P_13936_out0 = v$G2_5329_out0;
assign v$P_13937_out0 = v$G2_5330_out0;
assign v$P_13938_out0 = v$G2_5331_out0;
assign v$P_13939_out0 = v$G2_5332_out0;
assign v$G21_14019_out0 = v$G_10105_out0;
assign v$OUT_14901_out0 = v$MUX2_2492_out0;
assign v$OUT_14906_out0 = v$MUX2_2494_out0;
assign v$OUT_14949_out0 = v$MUX2_2506_out0;
assign v$OUT_14954_out0 = v$MUX2_2508_out0;
assign {v$A1_15221_out1,v$A1_15221_out0 } = v$_18000_out0 + v$MUX1_8345_out0 + v$C6_11357_out0;
assign v$P3_15337_out0 = v$P_13917_out0;
assign v$G0_15944_out0 = v$G_10115_out0;
assign v$G6_16355_out0 = v$G_10103_out0;
assign v$P9_18447_out0 = v$P_13919_out0;
assign v$P5_223_out0 = v$P_13938_out0;
assign v$P10_346_out0 = v$P_13934_out0;
assign v$G$CD_1006_out0 = v$G6_16355_out0;
assign v$G$CD_1007_out0 = v$G3_11106_out0;
assign v$G$CD_1008_out0 = v$G12_7044_out0;
assign v$G$CD_1009_out0 = v$G9_8927_out0;
assign v$G$CD_1012_out0 = v$G18_12940_out0;
assign v$G$CD_1023_out0 = v$G15_11032_out0;
assign v$G$CD_1024_out0 = v$G21_14019_out0;
assign v$G7_1693_out0 = v$G_10108_out0;
assign v$P8_1705_out0 = v$P_13925_out0;
assign v$G10_1835_out0 = v$G_10121_out0;
assign v$G19_1883_out0 = v$G_10118_out0;
assign v$P$AB_2087_out0 = v$P0_4812_out0;
assign v$P$AB_2090_out0 = v$P18_11724_out0;
assign v$P$AB_2091_out0 = v$P21_4771_out0;
assign v$P$AB_2103_out0 = v$P12_237_out0;
assign v$P$AB_2105_out0 = v$P15_6906_out0;
assign v$P$AB_2108_out0 = v$P6_8106_out0;
assign v$P$AB_2114_out0 = v$P3_15337_out0;
assign v$P$AB_2119_out0 = v$P9_18447_out0;
assign v$P2_2221_out0 = v$P_13936_out0;
assign v$G8_2579_out0 = v$G_10112_out0;
assign v$G13_2830_out0 = v$G_10116_out0;
assign v$P1_2961_out0 = v$P_13922_out0;
assign v$P13_3034_out0 = v$P_13929_out0;
assign v$P14_3153_out0 = v$P_13923_out0;
assign v$P22_4736_out0 = v$P_13932_out0;
assign v$G1_5055_out0 = v$G_10109_out0;
assign v$G4_5737_out0 = v$G_10117_out0;
assign v$P23_6388_out0 = v$P_13927_out0;
assign v$P16_6964_out0 = v$P_13939_out0;
assign v$COUT_8118_out0 = v$A1_15221_out1;
assign v$G20_8227_out0 = v$G_10122_out0;
assign v$G$AB_9222_out0 = v$G0_15944_out0;
assign v$G$AB_9225_out0 = v$G18_12940_out0;
assign v$G$AB_9226_out0 = v$G21_14019_out0;
assign v$G$AB_9238_out0 = v$G12_7044_out0;
assign v$G$AB_9240_out0 = v$G15_11032_out0;
assign v$G$AB_9243_out0 = v$G6_16355_out0;
assign v$G$AB_9249_out0 = v$G3_11106_out0;
assign v$G$AB_9254_out0 = v$G9_8927_out0;
assign v$G17_9348_out0 = v$G_10113_out0;
assign v$P11_9613_out0 = v$P_13937_out0;
assign v$P$CD_10546_out0 = v$P6_8106_out0;
assign v$P$CD_10547_out0 = v$P3_15337_out0;
assign v$P$CD_10548_out0 = v$P12_237_out0;
assign v$P$CD_10549_out0 = v$P9_18447_out0;
assign v$P$CD_10552_out0 = v$P18_11724_out0;
assign v$P$CD_10563_out0 = v$P15_6906_out0;
assign v$P$CD_10564_out0 = v$P21_4771_out0;
assign v$P20_10661_out0 = v$P_13935_out0;
assign v$G5_10678_out0 = v$G_10125_out0;
assign v$G11_11065_out0 = v$G_10124_out0;
assign v$MUX1_11630_out0 = v$G2_17411_out0 ? v$C1_4454_out0 : v$OUT_14901_out0;
assign v$MUX1_11631_out0 = v$G2_17412_out0 ? v$C1_4455_out0 : v$OUT_14906_out0;
assign v$MUX1_11635_out0 = v$G2_17416_out0 ? v$C1_4459_out0 : v$OUT_14949_out0;
assign v$MUX1_11636_out0 = v$G2_17417_out0 ? v$C1_4460_out0 : v$OUT_14954_out0;
assign v$P17_11761_out0 = v$P_13926_out0;
assign v$P7_11771_out0 = v$P_13921_out0;
assign v$G22_12512_out0 = v$G_10119_out0;
assign v$P4_13638_out0 = v$P_13930_out0;
assign v$G23_14319_out0 = v$G_10114_out0;
assign v$SUM_15173_out0 = v$A1_15221_out0;
assign v$GATE2_15758_out0 = v$CIN_16108_out0 && v$P0_4812_out0;
assign v$G2_15962_out0 = v$G_10123_out0;
assign v$P19_16319_out0 = v$P_13931_out0;
assign v$G16_16450_out0 = v$G_10126_out0;
assign v$G14_17978_out0 = v$G_10110_out0;
assign v$GATE1_661_out0 = v$GATE2_15758_out0 || v$G0_15944_out0;
assign v$G$CD_997_out0 = v$G14_17978_out0;
assign v$G$CD_998_out0 = v$G8_2579_out0;
assign v$G$CD_1000_out0 = v$G1_5055_out0;
assign v$G$CD_1003_out0 = v$G19_1883_out0;
assign v$G$CD_1004_out0 = v$G22_12512_out0;
assign v$G$CD_1011_out0 = v$G23_14319_out0;
assign v$G$CD_1013_out0 = v$G2_15962_out0;
assign v$G$CD_1014_out0 = v$G5_10678_out0;
assign v$G$CD_1016_out0 = v$G13_2830_out0;
assign v$G$CD_1017_out0 = v$G17_9348_out0;
assign v$G$CD_1018_out0 = v$G16_16450_out0;
assign v$G$CD_1021_out0 = v$G7_1693_out0;
assign v$G$CD_1027_out0 = v$G4_5737_out0;
assign v$G$CD_1031_out0 = v$G20_8227_out0;
assign v$G$CD_1032_out0 = v$G10_1835_out0;
assign v$G$CD_1036_out0 = v$G11_11065_out0;
assign v$SUM_3473_out0 = v$SUM_15173_out0;
assign v$OUT_10011_out0 = v$MUX1_11630_out0;
assign v$OUT_10012_out0 = v$MUX1_11631_out0;
assign v$OUT_10016_out0 = v$MUX1_11635_out0;
assign v$OUT_10017_out0 = v$MUX1_11636_out0;
assign v$P$CD_10537_out0 = v$P14_3153_out0;
assign v$P$CD_10538_out0 = v$P8_1705_out0;
assign v$P$CD_10540_out0 = v$P1_2961_out0;
assign v$P$CD_10543_out0 = v$P19_16319_out0;
assign v$P$CD_10544_out0 = v$P22_4736_out0;
assign v$P$CD_10551_out0 = v$P23_6388_out0;
assign v$P$CD_10553_out0 = v$P2_2221_out0;
assign v$P$CD_10554_out0 = v$P5_223_out0;
assign v$P$CD_10556_out0 = v$P13_3034_out0;
assign v$P$CD_10557_out0 = v$P17_11761_out0;
assign v$P$CD_10558_out0 = v$P16_6964_out0;
assign v$P$CD_10561_out0 = v$P7_11771_out0;
assign v$P$CD_10567_out0 = v$P4_13638_out0;
assign v$P$CD_10571_out0 = v$P20_10661_out0;
assign v$P$CD_10572_out0 = v$P10_346_out0;
assign v$P$CD_10576_out0 = v$P11_9613_out0;
assign v$COUT_10735_out0 = v$COUT_8118_out0;
assign v$G8_11481_out0 = v$CINA_8550_out0 && v$P$AB_2087_out0;
assign v$G8_11484_out0 = v$CINA_8553_out0 && v$P$AB_2090_out0;
assign v$G8_11485_out0 = v$CINA_8554_out0 && v$P$AB_2091_out0;
assign v$G8_11497_out0 = v$CINA_8566_out0 && v$P$AB_2103_out0;
assign v$G8_11499_out0 = v$CINA_8568_out0 && v$P$AB_2105_out0;
assign v$G8_11502_out0 = v$CINA_8571_out0 && v$P$AB_2108_out0;
assign v$G8_11508_out0 = v$CINA_8577_out0 && v$P$AB_2114_out0;
assign v$G8_11513_out0 = v$CINA_8582_out0 && v$P$AB_2119_out0;
assign v$CIN_3895_out0 = v$COUT_10735_out0;
assign v$G5_4605_out0 = v$G$AB_9222_out0 && v$P$CD_10540_out0;
assign v$G5_4608_out0 = v$G$AB_9225_out0 && v$P$CD_10543_out0;
assign v$G5_4609_out0 = v$G$AB_9226_out0 && v$P$CD_10544_out0;
assign v$G5_4621_out0 = v$G$AB_9238_out0 && v$P$CD_10556_out0;
assign v$G5_4623_out0 = v$G$AB_9240_out0 && v$P$CD_10558_out0;
assign v$G5_4626_out0 = v$G$AB_9243_out0 && v$P$CD_10561_out0;
assign v$G5_4632_out0 = v$G$AB_9249_out0 && v$P$CD_10567_out0;
assign v$G5_4637_out0 = v$G$AB_9254_out0 && v$P$CD_10572_out0;
assign v$G1_5608_out0 = v$P$AB_2087_out0 && v$P$CD_10540_out0;
assign v$G1_5611_out0 = v$P$AB_2090_out0 && v$P$CD_10543_out0;
assign v$G1_5612_out0 = v$P$AB_2091_out0 && v$P$CD_10544_out0;
assign v$G1_5624_out0 = v$P$AB_2103_out0 && v$P$CD_10556_out0;
assign v$G1_5626_out0 = v$P$AB_2105_out0 && v$P$CD_10558_out0;
assign v$G1_5629_out0 = v$P$AB_2108_out0 && v$P$CD_10561_out0;
assign v$G1_5635_out0 = v$P$AB_2114_out0 && v$P$CD_10567_out0;
assign v$G1_5640_out0 = v$P$AB_2119_out0 && v$P$CD_10572_out0;
assign v$MUX4_5890_out0 = v$NEED$SHIFT$OP1_4821_out0 ? v$OUT_10012_out0 : v$OP1$MANTISA_11806_out0;
assign v$MUX4_5891_out0 = v$NEED$SHIFT$OP1_4822_out0 ? v$OUT_10017_out0 : v$OP1$MANTISA_11807_out0;
assign v$G7_9721_out0 = v$G8_11481_out0 && v$P$CD_10540_out0;
assign v$G7_9724_out0 = v$G8_11484_out0 && v$P$CD_10543_out0;
assign v$G7_9725_out0 = v$G8_11485_out0 && v$P$CD_10544_out0;
assign v$G7_9737_out0 = v$G8_11497_out0 && v$P$CD_10556_out0;
assign v$G7_9739_out0 = v$G8_11499_out0 && v$P$CD_10558_out0;
assign v$G7_9742_out0 = v$G8_11502_out0 && v$P$CD_10561_out0;
assign v$G7_9748_out0 = v$G8_11508_out0 && v$P$CD_10567_out0;
assign v$G7_9753_out0 = v$G8_11513_out0 && v$P$CD_10572_out0;
assign v$C0_10694_out0 = v$GATE1_661_out0;
assign v$MUX1_14183_out0 = v$NEED$SHIFT$OP1_4821_out0 ? v$OP2$MANTISA_3510_out0 : v$OUT_10011_out0;
assign v$MUX1_14184_out0 = v$NEED$SHIFT$OP1_4822_out0 ? v$OP2$MANTISA_3511_out0 : v$OUT_10016_out0;
assign v$OP1_14194_out0 = v$SUM_3473_out0;
assign v$SEL2_14411_out0 = v$SUM_3473_out0[0:0];
assign v$P$AD_773_out0 = v$G1_5608_out0;
assign v$P$AD_776_out0 = v$G1_5611_out0;
assign v$P$AD_777_out0 = v$G1_5612_out0;
assign v$P$AD_789_out0 = v$G1_5624_out0;
assign v$P$AD_791_out0 = v$G1_5626_out0;
assign v$P$AD_794_out0 = v$G1_5629_out0;
assign v$P$AD_800_out0 = v$G1_5635_out0;
assign v$P$AD_805_out0 = v$G1_5640_out0;
assign {v$A2A_1633_out1,v$A2A_1633_out0 } = v$A1_1712_out0 + v$B1_8125_out0 + v$C0_10694_out0;
assign v$OP1_3388_out0 = v$OP1_14194_out0;
assign v$XOR2_7849_out0 = v$MUX1_14183_out0 ^ v$MUX3_3771_out0;
assign v$XOR2_7850_out0 = v$MUX1_14184_out0 ^ v$MUX3_3772_out0;
assign v$SUM$2_9082_out0 = v$SEL2_14411_out0;
assign v$C0_9376_out0 = v$C0_10694_out0;
assign v$G4_11197_out0 = v$G5_4605_out0 || v$G$CD_1000_out0;
assign v$G4_11200_out0 = v$G5_4608_out0 || v$G$CD_1003_out0;
assign v$G4_11201_out0 = v$G5_4609_out0 || v$G$CD_1004_out0;
assign v$G4_11213_out0 = v$G5_4621_out0 || v$G$CD_1016_out0;
assign v$G4_11215_out0 = v$G5_4623_out0 || v$G$CD_1018_out0;
assign v$G4_11218_out0 = v$G5_4626_out0 || v$G$CD_1021_out0;
assign v$G4_11224_out0 = v$G5_4632_out0 || v$G$CD_1027_out0;
assign v$G4_11229_out0 = v$G5_4637_out0 || v$G$CD_1032_out0;
assign v$A1_13596_out0 = v$MUX4_5890_out0;
assign v$A1_13599_out0 = v$MUX4_5891_out0;
assign v$CIN_16821_out0 = v$CIN_3895_out0;
assign v$G6_519_out0 = v$G4_11197_out0 || v$G7_9721_out0;
assign v$G6_522_out0 = v$G4_11200_out0 || v$G7_9724_out0;
assign v$G6_523_out0 = v$G4_11201_out0 || v$G7_9725_out0;
assign v$G6_535_out0 = v$G4_11213_out0 || v$G7_9737_out0;
assign v$G6_537_out0 = v$G4_11215_out0 || v$G7_9739_out0;
assign v$G6_540_out0 = v$G4_11218_out0 || v$G7_9742_out0;
assign v$G6_546_out0 = v$G4_11224_out0 || v$G7_9748_out0;
assign v$G6_551_out0 = v$G4_11229_out0 || v$G7_9753_out0;
assign v$END1_1545_out0 = v$A2A_1633_out1;
assign v$P$AB_2084_out0 = v$P$AD_789_out0;
assign v$P$AB_2085_out0 = v$P$AD_794_out0;
assign v$P$AB_2098_out0 = v$P$AD_777_out0;
assign v$P$AB_2100_out0 = v$P$AD_773_out0;
assign v$P$AB_2101_out0 = v$P$AD_800_out0;
assign v$P$AB_2104_out0 = v$P$AD_791_out0;
assign v$P$AB_2118_out0 = v$P$AD_776_out0;
assign v$P$AB_2123_out0 = v$P$AD_805_out0;
assign v$_7540_out0 = v$A1_13596_out0[11:0];
assign v$_7540_out1 = v$A1_13596_out0[23:12];
assign v$_7543_out0 = v$A1_13599_out0[11:0];
assign v$_7543_out1 = v$A1_13599_out0[23:12];
assign v$B2_8416_out0 = v$XOR2_7849_out0;
assign v$B2_8419_out0 = v$XOR2_7850_out0;
assign v$P$CD_10541_out0 = v$P$AD_800_out0;
assign v$P$CD_10545_out0 = v$P$AD_777_out0;
assign v$P$CD_10566_out0 = v$P$AD_791_out0;
assign v$P$CD_10569_out0 = v$P$AD_789_out0;
assign v$P$CD_10570_out0 = v$P$AD_805_out0;
assign v$P$CD_10574_out0 = v$P$AD_776_out0;
assign v$P$CD_10575_out0 = v$P$AD_794_out0;
assign v$_13439_out0 = { v$A1A_11662_out0,v$A2A_1633_out0 };
assign v$G$AD_17172_out0 = v$G4_11197_out0;
assign v$G$AD_17175_out0 = v$G4_11200_out0;
assign v$G$AD_17176_out0 = v$G4_11201_out0;
assign v$G$AD_17188_out0 = v$G4_11213_out0;
assign v$G$AD_17190_out0 = v$G4_11215_out0;
assign v$G$AD_17193_out0 = v$G4_11218_out0;
assign v$G$AD_17199_out0 = v$G4_11224_out0;
assign v$G$AD_17204_out0 = v$G4_11229_out0;
assign v$SEL8_17660_out0 = v$OP1_3388_out0[23:1];
assign v$G$CD_1001_out0 = v$G$AD_17199_out0;
assign v$G$CD_1005_out0 = v$G$AD_17176_out0;
assign v$G$CD_1026_out0 = v$G$AD_17190_out0;
assign v$G$CD_1029_out0 = v$G$AD_17188_out0;
assign v$G$CD_1030_out0 = v$G$AD_17204_out0;
assign v$G$CD_1034_out0 = v$G$AD_17175_out0;
assign v$G$CD_1035_out0 = v$G$AD_17193_out0;
assign v$_3986_out0 = v$B2_8416_out0[11:0];
assign v$_3986_out1 = v$B2_8416_out0[23:12];
assign v$_3989_out0 = v$B2_8419_out0[11:0];
assign v$_3989_out1 = v$B2_8419_out0[23:12];
assign v$G1_5605_out0 = v$P$AB_2084_out0 && v$P$CD_10537_out0;
assign v$G1_5606_out0 = v$P$AB_2085_out0 && v$P$CD_10538_out0;
assign v$G1_5619_out0 = v$P$AB_2098_out0 && v$P$CD_10551_out0;
assign v$G1_5621_out0 = v$P$AB_2100_out0 && v$P$CD_10553_out0;
assign v$G1_5622_out0 = v$P$AB_2101_out0 && v$P$CD_10554_out0;
assign v$G1_5625_out0 = v$P$AB_2104_out0 && v$P$CD_10557_out0;
assign v$G1_5639_out0 = v$P$AB_2118_out0 && v$P$CD_10571_out0;
assign v$G1_5644_out0 = v$P$AB_2123_out0 && v$P$CD_10576_out0;
assign v$COUTD_6779_out0 = v$G6_519_out0;
assign v$COUTD_6782_out0 = v$G6_522_out0;
assign v$COUTD_6783_out0 = v$G6_523_out0;
assign v$COUTD_6795_out0 = v$G6_535_out0;
assign v$COUTD_6797_out0 = v$G6_537_out0;
assign v$COUTD_6800_out0 = v$G6_540_out0;
assign v$COUTD_6806_out0 = v$G6_546_out0;
assign v$COUTD_6811_out0 = v$G6_551_out0;
assign v$G$AB_9219_out0 = v$G$AD_17188_out0;
assign v$G$AB_9220_out0 = v$G$AD_17193_out0;
assign v$G$AB_9233_out0 = v$G$AD_17176_out0;
assign v$G$AB_9235_out0 = v$G$AD_17172_out0;
assign v$G$AB_9236_out0 = v$G$AD_17199_out0;
assign v$G$AB_9239_out0 = v$G$AD_17190_out0;
assign v$G$AB_9253_out0 = v$G$AD_17175_out0;
assign v$G$AB_9258_out0 = v$G$AD_17204_out0;
assign v$_16112_out0 = v$_7540_out0[5:0];
assign v$_16112_out1 = v$_7540_out0[11:6];
assign v$_16115_out0 = v$_7543_out0[5:0];
assign v$_16115_out1 = v$_7543_out0[11:6];
assign v$_17029_out0 = v$_7540_out1[5:0];
assign v$_17029_out1 = v$_7540_out1[11:6];
assign v$_17032_out0 = v$_7543_out1[5:0];
assign v$_17032_out1 = v$_7543_out1[11:6];
assign v$_18002_out0 = { v$SEL8_17660_out0,v$CIN_16821_out0 };
assign v$P$AD_770_out0 = v$G1_5605_out0;
assign v$P$AD_771_out0 = v$G1_5606_out0;
assign v$P$AD_784_out0 = v$G1_5619_out0;
assign v$P$AD_786_out0 = v$G1_5621_out0;
assign v$P$AD_787_out0 = v$G1_5622_out0;
assign v$P$AD_790_out0 = v$G1_5625_out0;
assign v$P$AD_804_out0 = v$G1_5639_out0;
assign v$P$AD_809_out0 = v$G1_5644_out0;
assign v$_1219_out0 = v$_3986_out1[5:0];
assign v$_1219_out1 = v$_3986_out1[11:6];
assign v$_1222_out0 = v$_3989_out1[5:0];
assign v$_1222_out1 = v$_3989_out1[11:6];
assign v$_1524_out0 = v$_3986_out0[5:0];
assign v$_1524_out1 = v$_3986_out0[11:6];
assign v$_1527_out0 = v$_3989_out0[5:0];
assign v$_1527_out1 = v$_3989_out0[11:6];
assign v$_1864_out0 = v$_17029_out1[2:0];
assign v$_1864_out1 = v$_17029_out1[5:3];
assign v$_1867_out0 = v$_17032_out1[2:0];
assign v$_1867_out1 = v$_17032_out1[5:3];
assign v$G5_4602_out0 = v$G$AB_9219_out0 && v$P$CD_10537_out0;
assign v$G5_4603_out0 = v$G$AB_9220_out0 && v$P$CD_10538_out0;
assign v$G5_4616_out0 = v$G$AB_9233_out0 && v$P$CD_10551_out0;
assign v$G5_4618_out0 = v$G$AB_9235_out0 && v$P$CD_10553_out0;
assign v$G5_4619_out0 = v$G$AB_9236_out0 && v$P$CD_10554_out0;
assign v$G5_4622_out0 = v$G$AB_9239_out0 && v$P$CD_10557_out0;
assign v$G5_4636_out0 = v$G$AB_9253_out0 && v$P$CD_10571_out0;
assign v$G5_4641_out0 = v$G$AB_9258_out0 && v$P$CD_10576_out0;
assign v$CINA_8547_out0 = v$COUTD_6795_out0;
assign v$CINA_8548_out0 = v$COUTD_6800_out0;
assign v$CINA_8561_out0 = v$COUTD_6783_out0;
assign v$CINA_8563_out0 = v$COUTD_6779_out0;
assign v$CINA_8564_out0 = v$COUTD_6806_out0;
assign v$CINA_8567_out0 = v$COUTD_6797_out0;
assign v$CINA_8581_out0 = v$COUTD_6782_out0;
assign v$CINA_8586_out0 = v$COUTD_6811_out0;
assign v$_10049_out0 = v$_17029_out0[2:0];
assign v$_10049_out1 = v$_17029_out0[5:3];
assign v$_10052_out0 = v$_17032_out0[2:0];
assign v$_10052_out1 = v$_17032_out0[5:3];
assign v$_13771_out0 = v$_16112_out0[2:0];
assign v$_13771_out1 = v$_16112_out0[5:3];
assign v$_13774_out0 = v$_16115_out0[2:0];
assign v$_13774_out1 = v$_16115_out0[5:3];
assign {v$A1_15223_out1,v$A1_15223_out0 } = v$_18002_out0 + v$MUX1_8347_out0 + v$C6_11359_out0;
assign v$C1_16783_out0 = v$COUTD_6779_out0;
assign v$_18421_out0 = v$_16112_out1[2:0];
assign v$_18421_out1 = v$_16112_out1[5:3];
assign v$_18424_out0 = v$_16115_out1[2:0];
assign v$_18424_out1 = v$_16115_out1[5:3];
assign v$_1303_out0 = v$_18421_out0[0:0];
assign v$_1303_out1 = v$_18421_out0[2:2];
assign v$_1306_out0 = v$_18424_out0[0:0];
assign v$_1306_out1 = v$_18424_out0[2:2];
assign v$_1354_out0 = v$_13771_out1[0:0];
assign v$_1354_out1 = v$_13771_out1[2:2];
assign v$_1357_out0 = v$_13774_out1[0:0];
assign v$_1357_out1 = v$_13774_out1[2:2];
assign v$_1855_out0 = v$_1864_out1[0:0];
assign v$_1855_out1 = v$_1864_out1[2:2];
assign v$_1858_out0 = v$_1867_out1[0:0];
assign v$_1858_out1 = v$_1867_out1[2:2];
assign v$P$AB_2083_out0 = v$P$AD_771_out0;
assign v$P$AB_2088_out0 = v$P$AD_786_out0;
assign v$P$AB_2094_out0 = v$P$AD_786_out0;
assign v$P$AB_2097_out0 = v$P$AD_804_out0;
assign v$P$AB_2102_out0 = v$P$AD_770_out0;
assign v$P$AB_2115_out0 = v$P$AD_786_out0;
assign v$_7068_out0 = v$_13771_out0[0:0];
assign v$_7068_out1 = v$_13771_out0[2:2];
assign v$_7071_out0 = v$_13774_out0[0:0];
assign v$_7071_out1 = v$_13774_out0[2:2];
assign v$COUT_8120_out0 = v$A1_15223_out1;
assign v$_9934_out0 = v$_1219_out1[2:0];
assign v$_9934_out1 = v$_1219_out1[5:3];
assign v$_9937_out0 = v$_1222_out1[2:0];
assign v$_9937_out1 = v$_1222_out1[5:3];
assign v$_10447_out0 = v$_10049_out0[0:0];
assign v$_10447_out1 = v$_10049_out0[2:2];
assign v$_10450_out0 = v$_10052_out0[0:0];
assign v$_10450_out1 = v$_10052_out0[2:2];
assign v$P$CD_10536_out0 = v$P$AD_809_out0;
assign v$P$CD_10542_out0 = v$P$AD_771_out0;
assign v$P$CD_10550_out0 = v$P$AD_784_out0;
assign v$P$CD_10555_out0 = v$P$AD_790_out0;
assign v$P$CD_10559_out0 = v$P$AD_804_out0;
assign v$P$CD_10560_out0 = v$P$AD_770_out0;
assign v$P$CD_10568_out0 = v$P$AD_787_out0;
assign v$_10911_out0 = v$_18421_out1[0:0];
assign v$_10911_out1 = v$_18421_out1[2:2];
assign v$_10914_out0 = v$_18424_out1[0:0];
assign v$_10914_out1 = v$_18424_out1[2:2];
assign v$_11100_out0 = v$_1864_out0[0:0];
assign v$_11100_out1 = v$_1864_out0[2:2];
assign v$_11103_out0 = v$_1867_out0[0:0];
assign v$_11103_out1 = v$_1867_out0[2:2];
assign v$G4_11194_out0 = v$G5_4602_out0 || v$G$CD_997_out0;
assign v$G4_11195_out0 = v$G5_4603_out0 || v$G$CD_998_out0;
assign v$G4_11208_out0 = v$G5_4616_out0 || v$G$CD_1011_out0;
assign v$G4_11210_out0 = v$G5_4618_out0 || v$G$CD_1013_out0;
assign v$G4_11211_out0 = v$G5_4619_out0 || v$G$CD_1014_out0;
assign v$G4_11214_out0 = v$G5_4622_out0 || v$G$CD_1017_out0;
assign v$G4_11228_out0 = v$G5_4636_out0 || v$G$CD_1031_out0;
assign v$G4_11233_out0 = v$G5_4641_out0 || v$G$CD_1036_out0;
assign v$G8_11478_out0 = v$CINA_8547_out0 && v$P$AB_2084_out0;
assign v$G8_11479_out0 = v$CINA_8548_out0 && v$P$AB_2085_out0;
assign v$G8_11492_out0 = v$CINA_8561_out0 && v$P$AB_2098_out0;
assign v$G8_11494_out0 = v$CINA_8563_out0 && v$P$AB_2100_out0;
assign v$G8_11495_out0 = v$CINA_8564_out0 && v$P$AB_2101_out0;
assign v$G8_11498_out0 = v$CINA_8567_out0 && v$P$AB_2104_out0;
assign v$G8_11512_out0 = v$CINA_8581_out0 && v$P$AB_2118_out0;
assign v$G8_11517_out0 = v$CINA_8586_out0 && v$P$AB_2123_out0;
assign v$C1_11851_out0 = v$C1_16783_out0;
assign {v$A3A_11953_out1,v$A3A_11953_out0 } = v$A2_18268_out0 + v$B2_3115_out0 + v$C1_16783_out0;
assign v$_12988_out0 = v$_1524_out1[2:0];
assign v$_12988_out1 = v$_1524_out1[5:3];
assign v$_12991_out0 = v$_1527_out1[2:0];
assign v$_12991_out1 = v$_1527_out1[5:3];
assign v$_13742_out0 = v$_1524_out0[2:0];
assign v$_13742_out1 = v$_1524_out0[5:3];
assign v$_13745_out0 = v$_1527_out0[2:0];
assign v$_13745_out1 = v$_1527_out0[5:3];
assign v$SUM_15175_out0 = v$A1_15223_out0;
assign v$_16131_out0 = v$_10049_out1[0:0];
assign v$_16131_out1 = v$_10049_out1[2:2];
assign v$_16134_out0 = v$_10052_out1[0:0];
assign v$_16134_out1 = v$_10052_out1[2:2];
assign v$_17733_out0 = v$_1219_out0[2:0];
assign v$_17733_out1 = v$_1219_out0[5:3];
assign v$_17736_out0 = v$_1222_out0[2:0];
assign v$_17736_out1 = v$_1222_out0[5:3];
assign v$A6_309_out0 = v$_1303_out0;
assign v$A6_312_out0 = v$_1306_out0;
assign v$A21_2599_out0 = v$_1855_out0;
assign v$A21_2602_out0 = v$_1858_out0;
assign v$_2923_out0 = v$_13742_out0[0:0];
assign v$_2923_out1 = v$_13742_out0[2:2];
assign v$_2926_out0 = v$_13745_out0[0:0];
assign v$_2926_out1 = v$_13745_out0[2:2];
assign v$A12_3139_out0 = v$_10447_out0;
assign v$A12_3142_out0 = v$_10450_out0;
assign v$A9_3436_out0 = v$_10911_out0;
assign v$A9_3439_out0 = v$_10914_out0;
assign v$SUM_3475_out0 = v$SUM_15175_out0;
assign v$A0_4309_out0 = v$_7068_out0;
assign v$A0_4312_out0 = v$_7071_out0;
assign v$END2_5236_out0 = v$A3A_11953_out1;
assign v$G1_5604_out0 = v$P$AB_2083_out0 && v$P$CD_10536_out0;
assign v$G1_5609_out0 = v$P$AB_2088_out0 && v$P$CD_10541_out0;
assign v$G1_5615_out0 = v$P$AB_2094_out0 && v$P$CD_10547_out0;
assign v$G1_5618_out0 = v$P$AB_2097_out0 && v$P$CD_10550_out0;
assign v$G1_5623_out0 = v$P$AB_2102_out0 && v$P$CD_10555_out0;
assign v$G1_5636_out0 = v$P$AB_2115_out0 && v$P$CD_10568_out0;
assign v$_5949_out0 = v$_16131_out1[0:0];
assign v$_5949_out1 = v$_16131_out1[1:1];
assign v$_5952_out0 = v$_16134_out1[0:0];
assign v$_5952_out1 = v$_16134_out1[1:1];
assign v$_7359_out0 = v$_1354_out1[0:0];
assign v$_7359_out1 = v$_1354_out1[1:1];
assign v$_7362_out0 = v$_1357_out1[0:0];
assign v$_7362_out1 = v$_1357_out1[1:1];
assign v$_7769_out0 = v$_17733_out0[0:0];
assign v$_7769_out1 = v$_17733_out0[2:2];
assign v$_7772_out0 = v$_17736_out0[0:0];
assign v$_7772_out1 = v$_17736_out0[2:2];
assign v$_8908_out0 = { v$C0_9376_out0,v$C1_11851_out0 };
assign v$_9063_out0 = v$_9934_out1[0:0];
assign v$_9063_out1 = v$_9934_out1[2:2];
assign v$_9066_out0 = v$_9937_out1[0:0];
assign v$_9066_out1 = v$_9937_out1[2:2];
assign v$G7_9718_out0 = v$G8_11478_out0 && v$P$CD_10537_out0;
assign v$G7_9719_out0 = v$G8_11479_out0 && v$P$CD_10538_out0;
assign v$G7_9732_out0 = v$G8_11492_out0 && v$P$CD_10551_out0;
assign v$G7_9734_out0 = v$G8_11494_out0 && v$P$CD_10553_out0;
assign v$G7_9735_out0 = v$G8_11495_out0 && v$P$CD_10554_out0;
assign v$G7_9738_out0 = v$G8_11498_out0 && v$P$CD_10557_out0;
assign v$G7_9752_out0 = v$G8_11512_out0 && v$P$CD_10571_out0;
assign v$G7_9757_out0 = v$G8_11517_out0 && v$P$CD_10576_out0;
assign v$_10285_out0 = v$_1855_out1[0:0];
assign v$_10285_out1 = v$_1855_out1[1:1];
assign v$_10288_out0 = v$_1858_out1[0:0];
assign v$_10288_out1 = v$_1858_out1[1:1];
assign v$COUT_10737_out0 = v$COUT_8120_out0;
assign v$_10773_out0 = v$_12988_out1[0:0];
assign v$_10773_out1 = v$_12988_out1[2:2];
assign v$_10776_out0 = v$_12991_out1[0:0];
assign v$_10776_out1 = v$_12991_out1[2:2];
assign v$_11619_out0 = v$_7068_out1[0:0];
assign v$_11619_out1 = v$_7068_out1[1:1];
assign v$_11622_out0 = v$_7071_out1[0:0];
assign v$_11622_out1 = v$_7071_out1[1:1];
assign v$A3_14608_out0 = v$_1354_out0;
assign v$A3_14611_out0 = v$_1357_out0;
assign v$_15149_out0 = v$_9934_out0[0:0];
assign v$_15149_out1 = v$_9934_out0[2:2];
assign v$_15152_out0 = v$_9937_out0[0:0];
assign v$_15152_out1 = v$_9937_out0[2:2];
assign v$_15742_out0 = v$_1303_out1[0:0];
assign v$_15742_out1 = v$_1303_out1[1:1];
assign v$_15745_out0 = v$_1306_out1[0:0];
assign v$_15745_out1 = v$_1306_out1[1:1];
assign v$_16183_out0 = v$_10447_out1[0:0];
assign v$_16183_out1 = v$_10447_out1[1:1];
assign v$_16186_out0 = v$_10450_out1[0:0];
assign v$_16186_out1 = v$_10450_out1[1:1];
assign v$_16266_out0 = v$_17733_out1[0:0];
assign v$_16266_out1 = v$_17733_out1[2:2];
assign v$_16269_out0 = v$_17736_out1[0:0];
assign v$_16269_out1 = v$_17736_out1[2:2];
assign v$_16705_out0 = v$_11100_out1[0:0];
assign v$_16705_out1 = v$_11100_out1[1:1];
assign v$_16708_out0 = v$_11103_out1[0:0];
assign v$_16708_out1 = v$_11103_out1[1:1];
assign v$_16741_out0 = v$_13742_out1[0:0];
assign v$_16741_out1 = v$_13742_out1[2:2];
assign v$_16744_out0 = v$_13745_out1[0:0];
assign v$_16744_out1 = v$_13745_out1[2:2];
assign v$G$AD_17169_out0 = v$G4_11194_out0;
assign v$G$AD_17170_out0 = v$G4_11195_out0;
assign v$G$AD_17183_out0 = v$G4_11208_out0;
assign v$G$AD_17185_out0 = v$G4_11210_out0;
assign v$G$AD_17186_out0 = v$G4_11211_out0;
assign v$G$AD_17189_out0 = v$G4_11214_out0;
assign v$G$AD_17203_out0 = v$G4_11228_out0;
assign v$G$AD_17208_out0 = v$G4_11233_out0;
assign v$A15_17319_out0 = v$_16131_out0;
assign v$A15_17322_out0 = v$_16134_out0;
assign v$A18_17696_out0 = v$_11100_out0;
assign v$A18_17699_out0 = v$_11103_out0;
assign v$_17756_out0 = v$_10911_out1[0:0];
assign v$_17756_out1 = v$_10911_out1[1:1];
assign v$_17759_out0 = v$_10914_out1[0:0];
assign v$_17759_out1 = v$_10914_out1[1:1];
assign v$_18189_out0 = v$_12988_out0[0:0];
assign v$_18189_out1 = v$_12988_out0[2:2];
assign v$_18192_out0 = v$_12991_out0[0:0];
assign v$_18192_out1 = v$_12991_out0[2:2];
assign v$G6_516_out0 = v$G4_11194_out0 || v$G7_9718_out0;
assign v$G6_517_out0 = v$G4_11195_out0 || v$G7_9719_out0;
assign v$G6_530_out0 = v$G4_11208_out0 || v$G7_9732_out0;
assign v$G6_532_out0 = v$G4_11210_out0 || v$G7_9734_out0;
assign v$G6_533_out0 = v$G4_11211_out0 || v$G7_9735_out0;
assign v$G6_536_out0 = v$G4_11214_out0 || v$G7_9738_out0;
assign v$G6_550_out0 = v$G4_11228_out0 || v$G7_9752_out0;
assign v$G6_555_out0 = v$G4_11233_out0 || v$G7_9757_out0;
assign v$A14_677_out0 = v$_16183_out1;
assign v$A14_680_out0 = v$_16186_out1;
assign v$P$AD_769_out0 = v$G1_5604_out0;
assign v$P$AD_774_out0 = v$G1_5609_out0;
assign v$P$AD_780_out0 = v$G1_5615_out0;
assign v$P$AD_783_out0 = v$G1_5618_out0;
assign v$P$AD_788_out0 = v$G1_5623_out0;
assign v$P$AD_801_out0 = v$G1_5636_out0;
assign v$G$CD_996_out0 = v$G$AD_17208_out0;
assign v$G$CD_1002_out0 = v$G$AD_17170_out0;
assign v$G$CD_1010_out0 = v$G$AD_17183_out0;
assign v$G$CD_1015_out0 = v$G$AD_17189_out0;
assign v$G$CD_1019_out0 = v$G$AD_17203_out0;
assign v$G$CD_1020_out0 = v$G$AD_17169_out0;
assign v$G$CD_1028_out0 = v$G$AD_17186_out0;
assign v$A19_1214_out0 = v$_16705_out0;
assign v$A19_1217_out0 = v$_16708_out0;
assign v$A10_1549_out0 = v$_17756_out0;
assign v$A10_1552_out0 = v$_17759_out0;
assign v$SEL3_1698_out0 = v$SUM_3475_out0[0:0];
assign v$A1_1711_out0 = v$_11619_out0;
assign v$A1_1714_out0 = v$_11622_out0;
assign v$B12_1951_out0 = v$_7769_out0;
assign v$B12_1954_out0 = v$_7772_out0;
assign v$B0_3201_out0 = v$_2923_out0;
assign v$B0_3204_out0 = v$_2926_out0;
assign v$CIN_3896_out0 = v$COUT_10737_out0;
assign v$B9_4066_out0 = v$_10773_out0;
assign v$B9_4069_out0 = v$_10776_out0;
assign v$A22_4425_out0 = v$_10285_out0;
assign v$A22_4428_out0 = v$_10288_out0;
assign v$A20_4437_out0 = v$_16705_out1;
assign v$A20_4440_out0 = v$_16708_out1;
assign v$A23_5064_out0 = v$_10285_out1;
assign v$A23_5067_out0 = v$_10288_out1;
assign v$A5_6666_out0 = v$_7359_out1;
assign v$A5_6669_out0 = v$_7362_out1;
assign v$_6899_out0 = v$_18189_out1[0:0];
assign v$_6899_out1 = v$_18189_out1[1:1];
assign v$_6902_out0 = v$_18192_out1[0:0];
assign v$_6902_out1 = v$_18192_out1[1:1];
assign v$_6978_out0 = v$_16741_out1[0:0];
assign v$_6978_out1 = v$_16741_out1[1:1];
assign v$_6981_out0 = v$_16744_out1[0:0];
assign v$_6981_out1 = v$_16744_out1[1:1];
assign v$A_7125_out0 = v$A6_309_out0;
assign v$A_7126_out0 = v$A3_14608_out0;
assign v$A_7127_out0 = v$A21_2599_out0;
assign v$A_7128_out0 = v$A9_3436_out0;
assign v$A_7129_out0 = v$A15_17319_out0;
assign v$A_7133_out0 = v$A12_3139_out0;
assign v$A_7137_out0 = v$A0_4309_out0;
assign v$A_7142_out0 = v$A18_17696_out0;
assign v$A_7197_out0 = v$A6_312_out0;
assign v$A_7198_out0 = v$A3_14611_out0;
assign v$A_7199_out0 = v$A21_2602_out0;
assign v$A_7200_out0 = v$A9_3439_out0;
assign v$A_7201_out0 = v$A15_17322_out0;
assign v$A_7205_out0 = v$A12_3142_out0;
assign v$A_7209_out0 = v$A0_4312_out0;
assign v$A_7214_out0 = v$A18_17699_out0;
assign v$G$AB_9218_out0 = v$G$AD_17170_out0;
assign v$G$AB_9223_out0 = v$G$AD_17185_out0;
assign v$G$AB_9229_out0 = v$G$AD_17185_out0;
assign v$G$AB_9232_out0 = v$G$AD_17203_out0;
assign v$G$AB_9237_out0 = v$G$AD_17169_out0;
assign v$G$AB_9250_out0 = v$G$AD_17185_out0;
assign v$_9382_out0 = v$_9063_out1[0:0];
assign v$_9382_out1 = v$_9063_out1[1:1];
assign v$_9385_out0 = v$_9066_out1[0:0];
assign v$_9385_out1 = v$_9066_out1[1:1];
assign v$B3_9472_out0 = v$_16741_out0;
assign v$B3_9475_out0 = v$_16744_out0;
assign v$_9498_out0 = v$_10773_out1[0:0];
assign v$_9498_out1 = v$_10773_out1[1:1];
assign v$_9501_out0 = v$_10776_out1[0:0];
assign v$_9501_out1 = v$_10776_out1[1:1];
assign v$A11_9963_out0 = v$_17756_out1;
assign v$A11_9966_out0 = v$_17759_out1;
assign v$B15_10022_out0 = v$_16266_out0;
assign v$B15_10025_out0 = v$_16269_out0;
assign v$B18_10868_out0 = v$_15149_out0;
assign v$B18_10871_out0 = v$_15152_out0;
assign v$_11023_out0 = v$_2923_out1[0:0];
assign v$_11023_out1 = v$_2923_out1[1:1];
assign v$_11026_out0 = v$_2926_out1[0:0];
assign v$_11026_out1 = v$_2926_out1[1:1];
assign v$_13181_out0 = v$_16266_out1[0:0];
assign v$_13181_out1 = v$_16266_out1[1:1];
assign v$_13184_out0 = v$_16269_out1[0:0];
assign v$_13184_out1 = v$_16269_out1[1:1];
assign v$B6_13299_out0 = v$_18189_out0;
assign v$B6_13302_out0 = v$_18192_out0;
assign v$A16_13615_out0 = v$_5949_out0;
assign v$A16_13618_out0 = v$_5952_out0;
assign v$A13_13863_out0 = v$_16183_out0;
assign v$A13_13866_out0 = v$_16186_out0;
assign v$OP1_14195_out0 = v$SUM_3475_out0;
assign v$A7_15308_out0 = v$_15742_out0;
assign v$A7_15311_out0 = v$_15745_out0;
assign v$_16590_out0 = v$_15149_out1[0:0];
assign v$_16590_out1 = v$_15149_out1[1:1];
assign v$_16593_out0 = v$_15152_out1[0:0];
assign v$_16593_out1 = v$_15152_out1[1:1];
assign v$A17_16723_out0 = v$_5949_out1;
assign v$A17_16726_out0 = v$_5952_out1;
assign v$_17326_out0 = v$_7769_out1[0:0];
assign v$_17326_out1 = v$_7769_out1[1:1];
assign v$_17329_out0 = v$_7772_out1[0:0];
assign v$_17329_out1 = v$_7772_out1[1:1];
assign v$A4_17499_out0 = v$_7359_out0;
assign v$A4_17502_out0 = v$_7362_out0;
assign v$B21_18083_out0 = v$_9063_out0;
assign v$B21_18086_out0 = v$_9066_out0;
assign v$A8_18091_out0 = v$_15742_out1;
assign v$A8_18094_out0 = v$_15745_out1;
assign v$A2_18267_out0 = v$_11619_out1;
assign v$A2_18270_out0 = v$_11622_out1;
assign v$B23_1284_out0 = v$_9382_out1;
assign v$B23_1287_out0 = v$_9385_out1;
assign v$P$AB_2089_out0 = v$P$AD_801_out0;
assign v$P$AB_2093_out0 = v$P$AD_801_out0;
assign v$P$AB_2112_out0 = v$P$AD_801_out0;
assign v$P$AB_2120_out0 = v$P$AD_788_out0;
assign v$P$AB_2122_out0 = v$P$AD_801_out0;
assign v$B_2720_out0 = v$B6_13299_out0;
assign v$B_2721_out0 = v$B3_9472_out0;
assign v$B_2722_out0 = v$B21_18083_out0;
assign v$B_2723_out0 = v$B9_4066_out0;
assign v$B_2724_out0 = v$B15_10022_out0;
assign v$B_2728_out0 = v$B12_1951_out0;
assign v$B_2732_out0 = v$B0_3201_out0;
assign v$B_2737_out0 = v$B18_10868_out0;
assign v$B_2792_out0 = v$B6_13302_out0;
assign v$B_2793_out0 = v$B3_9475_out0;
assign v$B_2794_out0 = v$B21_18086_out0;
assign v$B_2795_out0 = v$B9_4069_out0;
assign v$B_2796_out0 = v$B15_10025_out0;
assign v$B_2800_out0 = v$B12_1954_out0;
assign v$B_2804_out0 = v$B0_3204_out0;
assign v$B_2809_out0 = v$B18_10871_out0;
assign v$B2_3114_out0 = v$_11023_out1;
assign v$B2_3117_out0 = v$_11026_out1;
assign v$OP1_3389_out0 = v$OP1_14195_out0;
assign v$B20_3944_out0 = v$_16590_out1;
assign v$B20_3947_out0 = v$_16593_out1;
assign v$B14_4003_out0 = v$_17326_out1;
assign v$B14_4006_out0 = v$_17329_out1;
assign v$G5_4601_out0 = v$G$AB_9218_out0 && v$P$CD_10536_out0;
assign v$G5_4606_out0 = v$G$AB_9223_out0 && v$P$CD_10541_out0;
assign v$G5_4612_out0 = v$G$AB_9229_out0 && v$P$CD_10547_out0;
assign v$G5_4615_out0 = v$G$AB_9232_out0 && v$P$CD_10550_out0;
assign v$G5_4620_out0 = v$G$AB_9237_out0 && v$P$CD_10555_out0;
assign v$G5_4633_out0 = v$G$AB_9250_out0 && v$P$CD_10568_out0;
assign v$COUTD_6776_out0 = v$G6_516_out0;
assign v$COUTD_6777_out0 = v$G6_517_out0;
assign v$COUTD_6790_out0 = v$G6_530_out0;
assign v$COUTD_6792_out0 = v$G6_532_out0;
assign v$COUTD_6793_out0 = v$G6_533_out0;
assign v$COUTD_6796_out0 = v$G6_536_out0;
assign v$COUTD_6810_out0 = v$G6_550_out0;
assign v$COUTD_6815_out0 = v$G6_555_out0;
assign v$A_7130_out0 = v$A7_15308_out0;
assign v$A_7131_out0 = v$A1_1711_out0;
assign v$A_7132_out0 = v$A14_677_out0;
assign v$A_7134_out0 = v$A8_18091_out0;
assign v$A_7135_out0 = v$A17_16723_out0;
assign v$A_7136_out0 = v$A23_5064_out0;
assign v$A_7138_out0 = v$A13_13863_out0;
assign v$A_7139_out0 = v$A4_17499_out0;
assign v$A_7140_out0 = v$A19_1214_out0;
assign v$A_7141_out0 = v$A22_4425_out0;
assign v$A_7143_out0 = v$A10_1549_out0;
assign v$A_7144_out0 = v$A20_4437_out0;
assign v$A_7145_out0 = v$A2_18267_out0;
assign v$A_7146_out0 = v$A11_9963_out0;
assign v$A_7147_out0 = v$A5_6666_out0;
assign v$A_7148_out0 = v$A16_13615_out0;
assign v$A_7202_out0 = v$A7_15311_out0;
assign v$A_7203_out0 = v$A1_1714_out0;
assign v$A_7204_out0 = v$A14_680_out0;
assign v$A_7206_out0 = v$A8_18094_out0;
assign v$A_7207_out0 = v$A17_16726_out0;
assign v$A_7208_out0 = v$A23_5067_out0;
assign v$A_7210_out0 = v$A13_13866_out0;
assign v$A_7211_out0 = v$A4_17502_out0;
assign v$A_7212_out0 = v$A19_1217_out0;
assign v$A_7213_out0 = v$A22_4428_out0;
assign v$A_7215_out0 = v$A10_1552_out0;
assign v$A_7216_out0 = v$A20_4440_out0;
assign v$A_7217_out0 = v$A2_18270_out0;
assign v$A_7218_out0 = v$A11_9966_out0;
assign v$A_7219_out0 = v$A5_6669_out0;
assign v$A_7220_out0 = v$A16_13618_out0;
assign v$SUM$3_7904_out0 = v$SEL3_1698_out0;
assign v$B1_8124_out0 = v$_11023_out0;
assign v$B1_8127_out0 = v$_11026_out0;
assign v$B13_8676_out0 = v$_17326_out0;
assign v$B13_8679_out0 = v$_17329_out0;
assign v$B11_9117_out0 = v$_9498_out1;
assign v$B11_9120_out0 = v$_9501_out1;
assign v$B10_9878_out0 = v$_9498_out0;
assign v$B10_9881_out0 = v$_9501_out0;
assign v$P$CD_10539_out0 = v$P$AD_788_out0;
assign v$P$CD_10565_out0 = v$P$AD_769_out0;
assign v$P$CD_10573_out0 = v$P$AD_783_out0;
assign v$B22_10806_out0 = v$_9382_out0;
assign v$B22_10809_out0 = v$_9385_out0;
assign {v$A1A_11661_out1,v$A1A_11661_out0 } = v$A0_4309_out0 + v$B0_3201_out0 + v$C1_4465_out0;
assign {v$A1A_11664_out1,v$A1A_11664_out0 } = v$A0_4312_out0 + v$B0_3204_out0 + v$C1_4468_out0;
assign v$END11_12092_out0 = v$P$AD_780_out0;
assign v$B8_13139_out0 = v$_6899_out1;
assign v$B8_13142_out0 = v$_6902_out1;
assign v$B4_14664_out0 = v$_6978_out0;
assign v$B4_14667_out0 = v$_6981_out0;
assign v$B17_15536_out0 = v$_13181_out1;
assign v$B17_15539_out0 = v$_13184_out1;
assign v$B16_16415_out0 = v$_13181_out0;
assign v$B16_16418_out0 = v$_13184_out0;
assign v$B19_16790_out0 = v$_16590_out0;
assign v$B19_16793_out0 = v$_16593_out0;
assign v$CIN_16822_out0 = v$CIN_3896_out0;
assign v$B7_17041_out0 = v$_6899_out0;
assign v$B7_17044_out0 = v$_6902_out0;
assign v$END13_18069_out0 = v$P$AD_774_out0;
assign v$B5_18375_out0 = v$_6978_out1;
assign v$B5_18378_out0 = v$_6981_out1;
assign v$END1_1293_out0 = v$COUTD_6815_out0;
assign v$C2_2688_out0 = v$COUTD_6792_out0;
assign v$B_2725_out0 = v$B7_17041_out0;
assign v$B_2726_out0 = v$B1_8124_out0;
assign v$B_2727_out0 = v$B14_4003_out0;
assign v$B_2729_out0 = v$B8_13139_out0;
assign v$B_2730_out0 = v$B17_15536_out0;
assign v$B_2731_out0 = v$B23_1284_out0;
assign v$B_2733_out0 = v$B13_8676_out0;
assign v$B_2734_out0 = v$B4_14664_out0;
assign v$B_2735_out0 = v$B19_16790_out0;
assign v$B_2736_out0 = v$B22_10806_out0;
assign v$B_2738_out0 = v$B10_9878_out0;
assign v$B_2739_out0 = v$B20_3944_out0;
assign v$B_2740_out0 = v$B2_3114_out0;
assign v$B_2741_out0 = v$B11_9117_out0;
assign v$B_2742_out0 = v$B5_18375_out0;
assign v$B_2743_out0 = v$B16_16415_out0;
assign v$B_2797_out0 = v$B7_17044_out0;
assign v$B_2798_out0 = v$B1_8127_out0;
assign v$B_2799_out0 = v$B14_4006_out0;
assign v$B_2801_out0 = v$B8_13142_out0;
assign v$B_2802_out0 = v$B17_15539_out0;
assign v$B_2803_out0 = v$B23_1287_out0;
assign v$B_2805_out0 = v$B13_8679_out0;
assign v$B_2806_out0 = v$B4_14667_out0;
assign v$B_2807_out0 = v$B19_16793_out0;
assign v$B_2808_out0 = v$B22_10809_out0;
assign v$B_2810_out0 = v$B10_9881_out0;
assign v$B_2811_out0 = v$B20_3947_out0;
assign v$B_2812_out0 = v$B2_3117_out0;
assign v$B_2813_out0 = v$B11_9120_out0;
assign v$B_2814_out0 = v$B5_18378_out0;
assign v$B_2815_out0 = v$B16_16418_out0;
assign v$END_3321_out0 = v$COUTD_6793_out0;
assign v$END3_3447_out0 = v$COUTD_6790_out0;
assign v$G2_5285_out0 = ((v$A_7125_out0 && !v$B_2720_out0) || (!v$A_7125_out0) && v$B_2720_out0);
assign v$G2_5286_out0 = ((v$A_7126_out0 && !v$B_2721_out0) || (!v$A_7126_out0) && v$B_2721_out0);
assign v$G2_5287_out0 = ((v$A_7127_out0 && !v$B_2722_out0) || (!v$A_7127_out0) && v$B_2722_out0);
assign v$G2_5288_out0 = ((v$A_7128_out0 && !v$B_2723_out0) || (!v$A_7128_out0) && v$B_2723_out0);
assign v$G2_5289_out0 = ((v$A_7129_out0 && !v$B_2724_out0) || (!v$A_7129_out0) && v$B_2724_out0);
assign v$G2_5293_out0 = ((v$A_7133_out0 && !v$B_2728_out0) || (!v$A_7133_out0) && v$B_2728_out0);
assign v$G2_5297_out0 = ((v$A_7137_out0 && !v$B_2732_out0) || (!v$A_7137_out0) && v$B_2732_out0);
assign v$G2_5302_out0 = ((v$A_7142_out0 && !v$B_2737_out0) || (!v$A_7142_out0) && v$B_2737_out0);
assign v$G2_5357_out0 = ((v$A_7197_out0 && !v$B_2792_out0) || (!v$A_7197_out0) && v$B_2792_out0);
assign v$G2_5358_out0 = ((v$A_7198_out0 && !v$B_2793_out0) || (!v$A_7198_out0) && v$B_2793_out0);
assign v$G2_5359_out0 = ((v$A_7199_out0 && !v$B_2794_out0) || (!v$A_7199_out0) && v$B_2794_out0);
assign v$G2_5360_out0 = ((v$A_7200_out0 && !v$B_2795_out0) || (!v$A_7200_out0) && v$B_2795_out0);
assign v$G2_5361_out0 = ((v$A_7201_out0 && !v$B_2796_out0) || (!v$A_7201_out0) && v$B_2796_out0);
assign v$G2_5365_out0 = ((v$A_7205_out0 && !v$B_2800_out0) || (!v$A_7205_out0) && v$B_2800_out0);
assign v$G2_5369_out0 = ((v$A_7209_out0 && !v$B_2804_out0) || (!v$A_7209_out0) && v$B_2804_out0);
assign v$G2_5374_out0 = ((v$A_7214_out0 && !v$B_2809_out0) || (!v$A_7214_out0) && v$B_2809_out0);
assign v$G1_5610_out0 = v$P$AB_2089_out0 && v$P$CD_10542_out0;
assign v$G1_5614_out0 = v$P$AB_2093_out0 && v$P$CD_10546_out0;
assign v$G1_5633_out0 = v$P$AB_2112_out0 && v$P$CD_10565_out0;
assign v$G1_5641_out0 = v$P$AB_2120_out0 && v$P$CD_10573_out0;
assign v$G1_5643_out0 = v$P$AB_2122_out0 && v$P$CD_10575_out0;
assign v$END2_7753_out0 = v$COUTD_6796_out0;
assign v$CINA_8546_out0 = v$COUTD_6777_out0;
assign v$CINA_8551_out0 = v$COUTD_6792_out0;
assign v$CINA_8557_out0 = v$COUTD_6792_out0;
assign v$CINA_8560_out0 = v$COUTD_6810_out0;
assign v$CINA_8565_out0 = v$COUTD_6776_out0;
assign v$CINA_8578_out0 = v$COUTD_6792_out0;
assign v$END45_9059_out0 = v$COUTD_6810_out0;
assign v$G4_11193_out0 = v$G5_4601_out0 || v$G$CD_996_out0;
assign v$G4_11198_out0 = v$G5_4606_out0 || v$G$CD_1001_out0;
assign v$G4_11204_out0 = v$G5_4612_out0 || v$G$CD_1007_out0;
assign v$G4_11207_out0 = v$G5_4615_out0 || v$G$CD_1010_out0;
assign v$G4_11212_out0 = v$G5_4620_out0 || v$G$CD_1015_out0;
assign v$G4_11225_out0 = v$G5_4633_out0 || v$G$CD_1028_out0;
assign v$G1_12359_out0 = v$A_7125_out0 && v$B_2720_out0;
assign v$G1_12360_out0 = v$A_7126_out0 && v$B_2721_out0;
assign v$G1_12361_out0 = v$A_7127_out0 && v$B_2722_out0;
assign v$G1_12362_out0 = v$A_7128_out0 && v$B_2723_out0;
assign v$G1_12363_out0 = v$A_7129_out0 && v$B_2724_out0;
assign v$G1_12367_out0 = v$A_7133_out0 && v$B_2728_out0;
assign v$G1_12371_out0 = v$A_7137_out0 && v$B_2732_out0;
assign v$G1_12376_out0 = v$A_7142_out0 && v$B_2737_out0;
assign v$G1_12431_out0 = v$A_7197_out0 && v$B_2792_out0;
assign v$G1_12432_out0 = v$A_7198_out0 && v$B_2793_out0;
assign v$G1_12433_out0 = v$A_7199_out0 && v$B_2794_out0;
assign v$G1_12434_out0 = v$A_7200_out0 && v$B_2795_out0;
assign v$G1_12435_out0 = v$A_7201_out0 && v$B_2796_out0;
assign v$G1_12439_out0 = v$A_7205_out0 && v$B_2800_out0;
assign v$G1_12443_out0 = v$A_7209_out0 && v$B_2804_out0;
assign v$G1_12448_out0 = v$A_7214_out0 && v$B_2809_out0;
assign v$SEL8_17661_out0 = v$OP1_3389_out0[23:1];
assign v$END_18273_out0 = v$A1A_11661_out1;
assign v$END_18276_out0 = v$A1A_11664_out1;
assign v$P$AD_775_out0 = v$G1_5610_out0;
assign v$P$AD_779_out0 = v$G1_5614_out0;
assign v$P$AD_798_out0 = v$G1_5633_out0;
assign v$P$AD_806_out0 = v$G1_5641_out0;
assign v$P$AD_808_out0 = v$G1_5643_out0;
assign v$G2_5290_out0 = ((v$A_7130_out0 && !v$B_2725_out0) || (!v$A_7130_out0) && v$B_2725_out0);
assign v$G2_5291_out0 = ((v$A_7131_out0 && !v$B_2726_out0) || (!v$A_7131_out0) && v$B_2726_out0);
assign v$G2_5292_out0 = ((v$A_7132_out0 && !v$B_2727_out0) || (!v$A_7132_out0) && v$B_2727_out0);
assign v$G2_5294_out0 = ((v$A_7134_out0 && !v$B_2729_out0) || (!v$A_7134_out0) && v$B_2729_out0);
assign v$G2_5295_out0 = ((v$A_7135_out0 && !v$B_2730_out0) || (!v$A_7135_out0) && v$B_2730_out0);
assign v$G2_5296_out0 = ((v$A_7136_out0 && !v$B_2731_out0) || (!v$A_7136_out0) && v$B_2731_out0);
assign v$G2_5298_out0 = ((v$A_7138_out0 && !v$B_2733_out0) || (!v$A_7138_out0) && v$B_2733_out0);
assign v$G2_5299_out0 = ((v$A_7139_out0 && !v$B_2734_out0) || (!v$A_7139_out0) && v$B_2734_out0);
assign v$G2_5300_out0 = ((v$A_7140_out0 && !v$B_2735_out0) || (!v$A_7140_out0) && v$B_2735_out0);
assign v$G2_5301_out0 = ((v$A_7141_out0 && !v$B_2736_out0) || (!v$A_7141_out0) && v$B_2736_out0);
assign v$G2_5303_out0 = ((v$A_7143_out0 && !v$B_2738_out0) || (!v$A_7143_out0) && v$B_2738_out0);
assign v$G2_5304_out0 = ((v$A_7144_out0 && !v$B_2739_out0) || (!v$A_7144_out0) && v$B_2739_out0);
assign v$G2_5305_out0 = ((v$A_7145_out0 && !v$B_2740_out0) || (!v$A_7145_out0) && v$B_2740_out0);
assign v$G2_5306_out0 = ((v$A_7146_out0 && !v$B_2741_out0) || (!v$A_7146_out0) && v$B_2741_out0);
assign v$G2_5307_out0 = ((v$A_7147_out0 && !v$B_2742_out0) || (!v$A_7147_out0) && v$B_2742_out0);
assign v$G2_5308_out0 = ((v$A_7148_out0 && !v$B_2743_out0) || (!v$A_7148_out0) && v$B_2743_out0);
assign v$G2_5362_out0 = ((v$A_7202_out0 && !v$B_2797_out0) || (!v$A_7202_out0) && v$B_2797_out0);
assign v$G2_5363_out0 = ((v$A_7203_out0 && !v$B_2798_out0) || (!v$A_7203_out0) && v$B_2798_out0);
assign v$G2_5364_out0 = ((v$A_7204_out0 && !v$B_2799_out0) || (!v$A_7204_out0) && v$B_2799_out0);
assign v$G2_5366_out0 = ((v$A_7206_out0 && !v$B_2801_out0) || (!v$A_7206_out0) && v$B_2801_out0);
assign v$G2_5367_out0 = ((v$A_7207_out0 && !v$B_2802_out0) || (!v$A_7207_out0) && v$B_2802_out0);
assign v$G2_5368_out0 = ((v$A_7208_out0 && !v$B_2803_out0) || (!v$A_7208_out0) && v$B_2803_out0);
assign v$G2_5370_out0 = ((v$A_7210_out0 && !v$B_2805_out0) || (!v$A_7210_out0) && v$B_2805_out0);
assign v$G2_5371_out0 = ((v$A_7211_out0 && !v$B_2806_out0) || (!v$A_7211_out0) && v$B_2806_out0);
assign v$G2_5372_out0 = ((v$A_7212_out0 && !v$B_2807_out0) || (!v$A_7212_out0) && v$B_2807_out0);
assign v$G2_5373_out0 = ((v$A_7213_out0 && !v$B_2808_out0) || (!v$A_7213_out0) && v$B_2808_out0);
assign v$G2_5375_out0 = ((v$A_7215_out0 && !v$B_2810_out0) || (!v$A_7215_out0) && v$B_2810_out0);
assign v$G2_5376_out0 = ((v$A_7216_out0 && !v$B_2811_out0) || (!v$A_7216_out0) && v$B_2811_out0);
assign v$G2_5377_out0 = ((v$A_7217_out0 && !v$B_2812_out0) || (!v$A_7217_out0) && v$B_2812_out0);
assign v$G2_5378_out0 = ((v$A_7218_out0 && !v$B_2813_out0) || (!v$A_7218_out0) && v$B_2813_out0);
assign v$G2_5379_out0 = ((v$A_7219_out0 && !v$B_2814_out0) || (!v$A_7219_out0) && v$B_2814_out0);
assign v$G2_5380_out0 = ((v$A_7220_out0 && !v$B_2815_out0) || (!v$A_7220_out0) && v$B_2815_out0);
assign v$G_10079_out0 = v$G1_12359_out0;
assign v$G_10080_out0 = v$G1_12360_out0;
assign v$G_10081_out0 = v$G1_12361_out0;
assign v$G_10082_out0 = v$G1_12362_out0;
assign v$G_10083_out0 = v$G1_12363_out0;
assign v$G_10087_out0 = v$G1_12367_out0;
assign v$G_10091_out0 = v$G1_12371_out0;
assign v$G_10096_out0 = v$G1_12376_out0;
assign v$G_10151_out0 = v$G1_12431_out0;
assign v$G_10152_out0 = v$G1_12432_out0;
assign v$G_10153_out0 = v$G1_12433_out0;
assign v$G_10154_out0 = v$G1_12434_out0;
assign v$G_10155_out0 = v$G1_12435_out0;
assign v$G_10159_out0 = v$G1_12439_out0;
assign v$G_10163_out0 = v$G1_12443_out0;
assign v$G_10168_out0 = v$G1_12448_out0;
assign v$G8_11477_out0 = v$CINA_8546_out0 && v$P$AB_2083_out0;
assign v$G8_11482_out0 = v$CINA_8551_out0 && v$P$AB_2088_out0;
assign v$G8_11488_out0 = v$CINA_8557_out0 && v$P$AB_2094_out0;
assign v$G8_11491_out0 = v$CINA_8560_out0 && v$P$AB_2097_out0;
assign v$G8_11496_out0 = v$CINA_8565_out0 && v$P$AB_2102_out0;
assign v$G8_11509_out0 = v$CINA_8578_out0 && v$P$AB_2115_out0;
assign v$G1_12364_out0 = v$A_7130_out0 && v$B_2725_out0;
assign v$G1_12365_out0 = v$A_7131_out0 && v$B_2726_out0;
assign v$G1_12366_out0 = v$A_7132_out0 && v$B_2727_out0;
assign v$G1_12368_out0 = v$A_7134_out0 && v$B_2729_out0;
assign v$G1_12369_out0 = v$A_7135_out0 && v$B_2730_out0;
assign v$G1_12370_out0 = v$A_7136_out0 && v$B_2731_out0;
assign v$G1_12372_out0 = v$A_7138_out0 && v$B_2733_out0;
assign v$G1_12373_out0 = v$A_7139_out0 && v$B_2734_out0;
assign v$G1_12374_out0 = v$A_7140_out0 && v$B_2735_out0;
assign v$G1_12375_out0 = v$A_7141_out0 && v$B_2736_out0;
assign v$G1_12377_out0 = v$A_7143_out0 && v$B_2738_out0;
assign v$G1_12378_out0 = v$A_7144_out0 && v$B_2739_out0;
assign v$G1_12379_out0 = v$A_7145_out0 && v$B_2740_out0;
assign v$G1_12380_out0 = v$A_7146_out0 && v$B_2741_out0;
assign v$G1_12381_out0 = v$A_7147_out0 && v$B_2742_out0;
assign v$G1_12382_out0 = v$A_7148_out0 && v$B_2743_out0;
assign v$G1_12436_out0 = v$A_7202_out0 && v$B_2797_out0;
assign v$G1_12437_out0 = v$A_7203_out0 && v$B_2798_out0;
assign v$G1_12438_out0 = v$A_7204_out0 && v$B_2799_out0;
assign v$G1_12440_out0 = v$A_7206_out0 && v$B_2801_out0;
assign v$G1_12441_out0 = v$A_7207_out0 && v$B_2802_out0;
assign v$G1_12442_out0 = v$A_7208_out0 && v$B_2803_out0;
assign v$G1_12444_out0 = v$A_7210_out0 && v$B_2805_out0;
assign v$G1_12445_out0 = v$A_7211_out0 && v$B_2806_out0;
assign v$G1_12446_out0 = v$A_7212_out0 && v$B_2807_out0;
assign v$G1_12447_out0 = v$A_7213_out0 && v$B_2808_out0;
assign v$G1_12449_out0 = v$A_7215_out0 && v$B_2810_out0;
assign v$G1_12450_out0 = v$A_7216_out0 && v$B_2811_out0;
assign v$G1_12451_out0 = v$A_7217_out0 && v$B_2812_out0;
assign v$G1_12452_out0 = v$A_7218_out0 && v$B_2813_out0;
assign v$G1_12453_out0 = v$A_7219_out0 && v$B_2814_out0;
assign v$G1_12454_out0 = v$A_7220_out0 && v$B_2815_out0;
assign {v$A4A_13156_out1,v$A4A_13156_out0 } = v$A3_14609_out0 + v$B3_9473_out0 + v$C2_2688_out0;
assign v$P_13892_out0 = v$G2_5285_out0;
assign v$P_13893_out0 = v$G2_5286_out0;
assign v$P_13894_out0 = v$G2_5287_out0;
assign v$P_13895_out0 = v$G2_5288_out0;
assign v$P_13896_out0 = v$G2_5289_out0;
assign v$P_13900_out0 = v$G2_5293_out0;
assign v$P_13904_out0 = v$G2_5297_out0;
assign v$P_13909_out0 = v$G2_5302_out0;
assign v$P_13964_out0 = v$G2_5357_out0;
assign v$P_13965_out0 = v$G2_5358_out0;
assign v$P_13966_out0 = v$G2_5359_out0;
assign v$P_13967_out0 = v$G2_5360_out0;
assign v$P_13968_out0 = v$G2_5361_out0;
assign v$P_13972_out0 = v$G2_5365_out0;
assign v$P_13976_out0 = v$G2_5369_out0;
assign v$P_13981_out0 = v$G2_5374_out0;
assign v$G$AD_17168_out0 = v$G4_11193_out0;
assign v$G$AD_17173_out0 = v$G4_11198_out0;
assign v$G$AD_17179_out0 = v$G4_11204_out0;
assign v$G$AD_17182_out0 = v$G4_11207_out0;
assign v$G$AD_17187_out0 = v$G4_11212_out0;
assign v$G$AD_17200_out0 = v$G4_11225_out0;
assign v$_18003_out0 = { v$SEL8_17661_out0,v$CIN_16822_out0 };
assign v$C2_18181_out0 = v$C2_2688_out0;
assign v$P12_236_out0 = v$P_13900_out0;
assign v$P12_239_out0 = v$P_13972_out0;
assign v$G$CD_999_out0 = v$G$AD_17187_out0;
assign v$G$CD_1025_out0 = v$G$AD_17168_out0;
assign v$G$CD_1033_out0 = v$G$AD_17182_out0;
assign v$END10_1153_out0 = v$G$AD_17179_out0;
assign v$P$AB_2086_out0 = v$P$AD_798_out0;
assign v$P$AB_2095_out0 = v$P$AD_798_out0;
assign v$P$AB_2096_out0 = v$P$AD_775_out0;
assign v$P$AB_2107_out0 = v$P$AD_798_out0;
assign v$P$AB_2109_out0 = v$P$AD_798_out0;
assign v$P$AB_2116_out0 = v$P$AD_798_out0;
assign v$P$AB_2117_out0 = v$P$AD_775_out0;
assign v$P21_4770_out0 = v$P_13894_out0;
assign v$P21_4773_out0 = v$P_13966_out0;
assign v$P0_4811_out0 = v$P_13904_out0;
assign v$P0_4814_out0 = v$P_13976_out0;
assign v$P15_6905_out0 = v$P_13896_out0;
assign v$P15_6908_out0 = v$P_13968_out0;
assign v$G12_7043_out0 = v$G_10087_out0;
assign v$G12_7046_out0 = v$G_10159_out0;
assign v$END15_7384_out0 = v$P$AD_779_out0;
assign v$END17_7639_out0 = v$P$AD_808_out0;
assign v$END3_7934_out0 = v$A4A_13156_out1;
assign v$P6_8105_out0 = v$P_13892_out0;
assign v$P6_8108_out0 = v$P_13964_out0;
assign v$G9_8926_out0 = v$G_10082_out0;
assign v$G9_8929_out0 = v$G_10154_out0;
assign v$G$AB_9224_out0 = v$G$AD_17200_out0;
assign v$G$AB_9228_out0 = v$G$AD_17200_out0;
assign v$G$AB_9247_out0 = v$G$AD_17200_out0;
assign v$G$AB_9255_out0 = v$G$AD_17187_out0;
assign v$G$AB_9257_out0 = v$G$AD_17200_out0;
assign v$G7_9717_out0 = v$G8_11477_out0 && v$P$CD_10536_out0;
assign v$G7_9722_out0 = v$G8_11482_out0 && v$P$CD_10541_out0;
assign v$G7_9728_out0 = v$G8_11488_out0 && v$P$CD_10547_out0;
assign v$G7_9731_out0 = v$G8_11491_out0 && v$P$CD_10550_out0;
assign v$G7_9736_out0 = v$G8_11496_out0 && v$P$CD_10555_out0;
assign v$G7_9749_out0 = v$G8_11509_out0 && v$P$CD_10568_out0;
assign v$G_10084_out0 = v$G1_12364_out0;
assign v$G_10085_out0 = v$G1_12365_out0;
assign v$G_10086_out0 = v$G1_12366_out0;
assign v$G_10088_out0 = v$G1_12368_out0;
assign v$G_10089_out0 = v$G1_12369_out0;
assign v$G_10090_out0 = v$G1_12370_out0;
assign v$G_10092_out0 = v$G1_12372_out0;
assign v$G_10093_out0 = v$G1_12373_out0;
assign v$G_10094_out0 = v$G1_12374_out0;
assign v$G_10095_out0 = v$G1_12375_out0;
assign v$G_10097_out0 = v$G1_12377_out0;
assign v$G_10098_out0 = v$G1_12378_out0;
assign v$G_10099_out0 = v$G1_12379_out0;
assign v$G_10100_out0 = v$G1_12380_out0;
assign v$G_10101_out0 = v$G1_12381_out0;
assign v$G_10102_out0 = v$G1_12382_out0;
assign v$G_10156_out0 = v$G1_12436_out0;
assign v$G_10157_out0 = v$G1_12437_out0;
assign v$G_10158_out0 = v$G1_12438_out0;
assign v$G_10160_out0 = v$G1_12440_out0;
assign v$G_10161_out0 = v$G1_12441_out0;
assign v$G_10162_out0 = v$G1_12442_out0;
assign v$G_10164_out0 = v$G1_12444_out0;
assign v$G_10165_out0 = v$G1_12445_out0;
assign v$G_10166_out0 = v$G1_12446_out0;
assign v$G_10167_out0 = v$G1_12447_out0;
assign v$G_10169_out0 = v$G1_12449_out0;
assign v$G_10170_out0 = v$G1_12450_out0;
assign v$G_10171_out0 = v$G1_12451_out0;
assign v$G_10172_out0 = v$G1_12452_out0;
assign v$G_10173_out0 = v$G1_12453_out0;
assign v$G_10174_out0 = v$G1_12454_out0;
assign v$P$CD_10562_out0 = v$P$AD_806_out0;
assign v$END12_10782_out0 = v$G$AD_17173_out0;
assign v$G15_11031_out0 = v$G_10083_out0;
assign v$G15_11034_out0 = v$G_10155_out0;
assign v$G3_11105_out0 = v$G_10080_out0;
assign v$G3_11108_out0 = v$G_10152_out0;
assign v$END19_11657_out0 = v$P$AD_775_out0;
assign v$P18_11723_out0 = v$P_13909_out0;
assign v$P18_11726_out0 = v$P_13981_out0;
assign v$G18_12939_out0 = v$G_10096_out0;
assign v$G18_12942_out0 = v$G_10168_out0;
assign v$P_13897_out0 = v$G2_5290_out0;
assign v$P_13898_out0 = v$G2_5291_out0;
assign v$P_13899_out0 = v$G2_5292_out0;
assign v$P_13901_out0 = v$G2_5294_out0;
assign v$P_13902_out0 = v$G2_5295_out0;
assign v$P_13903_out0 = v$G2_5296_out0;
assign v$P_13905_out0 = v$G2_5298_out0;
assign v$P_13906_out0 = v$G2_5299_out0;
assign v$P_13907_out0 = v$G2_5300_out0;
assign v$P_13908_out0 = v$G2_5301_out0;
assign v$P_13910_out0 = v$G2_5303_out0;
assign v$P_13911_out0 = v$G2_5304_out0;
assign v$P_13912_out0 = v$G2_5305_out0;
assign v$P_13913_out0 = v$G2_5306_out0;
assign v$P_13914_out0 = v$G2_5307_out0;
assign v$P_13915_out0 = v$G2_5308_out0;
assign v$P_13969_out0 = v$G2_5362_out0;
assign v$P_13970_out0 = v$G2_5363_out0;
assign v$P_13971_out0 = v$G2_5364_out0;
assign v$P_13973_out0 = v$G2_5366_out0;
assign v$P_13974_out0 = v$G2_5367_out0;
assign v$P_13975_out0 = v$G2_5368_out0;
assign v$P_13977_out0 = v$G2_5370_out0;
assign v$P_13978_out0 = v$G2_5371_out0;
assign v$P_13979_out0 = v$G2_5372_out0;
assign v$P_13980_out0 = v$G2_5373_out0;
assign v$P_13982_out0 = v$G2_5375_out0;
assign v$P_13983_out0 = v$G2_5376_out0;
assign v$P_13984_out0 = v$G2_5377_out0;
assign v$P_13985_out0 = v$G2_5378_out0;
assign v$P_13986_out0 = v$G2_5379_out0;
assign v$P_13987_out0 = v$G2_5380_out0;
assign v$G21_14018_out0 = v$G_10081_out0;
assign v$G21_14021_out0 = v$G_10153_out0;
assign {v$A1_15224_out1,v$A1_15224_out0 } = v$_18003_out0 + v$MUX1_8348_out0 + v$C6_11360_out0;
assign v$P3_15336_out0 = v$P_13893_out0;
assign v$P3_15339_out0 = v$P_13965_out0;
assign v$G0_15943_out0 = v$G_10091_out0;
assign v$G0_15946_out0 = v$G_10163_out0;
assign v$G6_16354_out0 = v$G_10079_out0;
assign v$G6_16357_out0 = v$G_10151_out0;
assign v$P9_18446_out0 = v$P_13895_out0;
assign v$P9_18449_out0 = v$P_13967_out0;
assign v$_18666_out0 = { v$A3A_11953_out0,v$A4A_13156_out0 };
assign v$P5_222_out0 = v$P_13914_out0;
assign v$P5_225_out0 = v$P_13986_out0;
assign v$P10_345_out0 = v$P_13910_out0;
assign v$P10_348_out0 = v$P_13982_out0;
assign v$G6_515_out0 = v$G4_11193_out0 || v$G7_9717_out0;
assign v$G6_520_out0 = v$G4_11198_out0 || v$G7_9722_out0;
assign v$G6_526_out0 = v$G4_11204_out0 || v$G7_9728_out0;
assign v$G6_529_out0 = v$G4_11207_out0 || v$G7_9731_out0;
assign v$G6_534_out0 = v$G4_11212_out0 || v$G7_9736_out0;
assign v$G6_547_out0 = v$G4_11225_out0 || v$G7_9749_out0;
assign v$G$CD_965_out0 = v$G6_16354_out0;
assign v$G$CD_966_out0 = v$G3_11105_out0;
assign v$G$CD_967_out0 = v$G12_7043_out0;
assign v$G$CD_968_out0 = v$G9_8926_out0;
assign v$G$CD_971_out0 = v$G18_12939_out0;
assign v$G$CD_982_out0 = v$G15_11031_out0;
assign v$G$CD_983_out0 = v$G21_14018_out0;
assign v$G$CD_1088_out0 = v$G6_16357_out0;
assign v$G$CD_1089_out0 = v$G3_11108_out0;
assign v$G$CD_1090_out0 = v$G12_7046_out0;
assign v$G$CD_1091_out0 = v$G9_8929_out0;
assign v$G$CD_1094_out0 = v$G18_12942_out0;
assign v$G$CD_1105_out0 = v$G15_11034_out0;
assign v$G$CD_1106_out0 = v$G21_14021_out0;
assign v$G7_1692_out0 = v$G_10084_out0;
assign v$G7_1695_out0 = v$G_10156_out0;
assign v$P8_1704_out0 = v$P_13901_out0;
assign v$P8_1707_out0 = v$P_13973_out0;
assign v$G10_1834_out0 = v$G_10097_out0;
assign v$G10_1837_out0 = v$G_10169_out0;
assign v$G19_1882_out0 = v$G_10094_out0;
assign v$G19_1885_out0 = v$G_10166_out0;
assign v$P$AB_2046_out0 = v$P0_4811_out0;
assign v$P$AB_2049_out0 = v$P18_11723_out0;
assign v$P$AB_2050_out0 = v$P21_4770_out0;
assign v$P$AB_2062_out0 = v$P12_236_out0;
assign v$P$AB_2064_out0 = v$P15_6905_out0;
assign v$P$AB_2067_out0 = v$P6_8105_out0;
assign v$P$AB_2073_out0 = v$P3_15336_out0;
assign v$P$AB_2078_out0 = v$P9_18446_out0;
assign v$P$AB_2169_out0 = v$P0_4814_out0;
assign v$P$AB_2172_out0 = v$P18_11726_out0;
assign v$P$AB_2173_out0 = v$P21_4773_out0;
assign v$P$AB_2185_out0 = v$P12_239_out0;
assign v$P$AB_2187_out0 = v$P15_6908_out0;
assign v$P$AB_2190_out0 = v$P6_8108_out0;
assign v$P$AB_2196_out0 = v$P3_15339_out0;
assign v$P$AB_2201_out0 = v$P9_18449_out0;
assign v$P2_2220_out0 = v$P_13912_out0;
assign v$P2_2223_out0 = v$P_13984_out0;
assign v$G8_2578_out0 = v$G_10088_out0;
assign v$G8_2581_out0 = v$G_10160_out0;
assign v$G13_2829_out0 = v$G_10092_out0;
assign v$G13_2832_out0 = v$G_10164_out0;
assign v$P1_2960_out0 = v$P_13898_out0;
assign v$P1_2963_out0 = v$P_13970_out0;
assign v$P13_3033_out0 = v$P_13905_out0;
assign v$P13_3036_out0 = v$P_13977_out0;
assign v$P14_3152_out0 = v$P_13899_out0;
assign v$P14_3155_out0 = v$P_13971_out0;
assign v$G5_4607_out0 = v$G$AB_9224_out0 && v$P$CD_10542_out0;
assign v$G5_4611_out0 = v$G$AB_9228_out0 && v$P$CD_10546_out0;
assign v$G5_4630_out0 = v$G$AB_9247_out0 && v$P$CD_10565_out0;
assign v$G5_4638_out0 = v$G$AB_9255_out0 && v$P$CD_10573_out0;
assign v$G5_4640_out0 = v$G$AB_9257_out0 && v$P$CD_10575_out0;
assign v$P22_4735_out0 = v$P_13908_out0;
assign v$P22_4738_out0 = v$P_13980_out0;
assign v$G1_5054_out0 = v$G_10085_out0;
assign v$G1_5057_out0 = v$G_10157_out0;
assign v$G1_5607_out0 = v$P$AB_2086_out0 && v$P$CD_10539_out0;
assign v$G1_5616_out0 = v$P$AB_2095_out0 && v$P$CD_10548_out0;
assign v$G1_5617_out0 = v$P$AB_2096_out0 && v$P$CD_10549_out0;
assign v$G1_5628_out0 = v$P$AB_2107_out0 && v$P$CD_10560_out0;
assign v$G1_5630_out0 = v$P$AB_2109_out0 && v$P$CD_10562_out0;
assign v$G1_5637_out0 = v$P$AB_2116_out0 && v$P$CD_10569_out0;
assign v$G1_5638_out0 = v$P$AB_2117_out0 && v$P$CD_10570_out0;
assign v$G4_5736_out0 = v$G_10093_out0;
assign v$G4_5739_out0 = v$G_10165_out0;
assign v$P23_6387_out0 = v$P_13903_out0;
assign v$P23_6390_out0 = v$P_13975_out0;
assign v$P16_6963_out0 = v$P_13915_out0;
assign v$P16_6966_out0 = v$P_13987_out0;
assign v$COUT_8121_out0 = v$A1_15224_out1;
assign v$G20_8226_out0 = v$G_10098_out0;
assign v$G20_8229_out0 = v$G_10170_out0;
assign v$G$AB_9181_out0 = v$G0_15943_out0;
assign v$G$AB_9184_out0 = v$G18_12939_out0;
assign v$G$AB_9185_out0 = v$G21_14018_out0;
assign v$G$AB_9197_out0 = v$G12_7043_out0;
assign v$G$AB_9199_out0 = v$G15_11031_out0;
assign v$G$AB_9202_out0 = v$G6_16354_out0;
assign v$G$AB_9208_out0 = v$G3_11105_out0;
assign v$G$AB_9213_out0 = v$G9_8926_out0;
assign v$G$AB_9304_out0 = v$G0_15946_out0;
assign v$G$AB_9307_out0 = v$G18_12942_out0;
assign v$G$AB_9308_out0 = v$G21_14021_out0;
assign v$G$AB_9320_out0 = v$G12_7046_out0;
assign v$G$AB_9322_out0 = v$G15_11034_out0;
assign v$G$AB_9325_out0 = v$G6_16357_out0;
assign v$G$AB_9331_out0 = v$G3_11108_out0;
assign v$G$AB_9336_out0 = v$G9_8929_out0;
assign v$G17_9347_out0 = v$G_10089_out0;
assign v$G17_9350_out0 = v$G_10161_out0;
assign v$P11_9612_out0 = v$P_13913_out0;
assign v$P11_9615_out0 = v$P_13985_out0;
assign v$_10357_out0 = { v$_13439_out0,v$_18666_out0 };
assign v$P$CD_10505_out0 = v$P6_8105_out0;
assign v$P$CD_10506_out0 = v$P3_15336_out0;
assign v$P$CD_10507_out0 = v$P12_236_out0;
assign v$P$CD_10508_out0 = v$P9_18446_out0;
assign v$P$CD_10511_out0 = v$P18_11723_out0;
assign v$P$CD_10522_out0 = v$P15_6905_out0;
assign v$P$CD_10523_out0 = v$P21_4770_out0;
assign v$P$CD_10628_out0 = v$P6_8108_out0;
assign v$P$CD_10629_out0 = v$P3_15339_out0;
assign v$P$CD_10630_out0 = v$P12_239_out0;
assign v$P$CD_10631_out0 = v$P9_18449_out0;
assign v$P$CD_10634_out0 = v$P18_11726_out0;
assign v$P$CD_10645_out0 = v$P15_6908_out0;
assign v$P$CD_10646_out0 = v$P21_4773_out0;
assign v$P20_10660_out0 = v$P_13911_out0;
assign v$P20_10663_out0 = v$P_13983_out0;
assign v$G5_10677_out0 = v$G_10101_out0;
assign v$G5_10680_out0 = v$G_10173_out0;
assign v$G11_11064_out0 = v$G_10100_out0;
assign v$G11_11067_out0 = v$G_10172_out0;
assign v$P17_11760_out0 = v$P_13902_out0;
assign v$P17_11763_out0 = v$P_13974_out0;
assign v$P7_11770_out0 = v$P_13897_out0;
assign v$P7_11773_out0 = v$P_13969_out0;
assign v$G22_12511_out0 = v$G_10095_out0;
assign v$G22_12514_out0 = v$G_10167_out0;
assign v$P4_13637_out0 = v$P_13906_out0;
assign v$P4_13640_out0 = v$P_13978_out0;
assign v$G23_14318_out0 = v$G_10090_out0;
assign v$G23_14321_out0 = v$G_10162_out0;
assign v$SUM_15176_out0 = v$A1_15224_out0;
assign v$GATE2_15757_out0 = v$CIN_16107_out0 && v$P0_4811_out0;
assign v$GATE2_15760_out0 = v$CIN_16110_out0 && v$P0_4814_out0;
assign v$G2_15961_out0 = v$G_10099_out0;
assign v$G2_15964_out0 = v$G_10171_out0;
assign v$P19_16318_out0 = v$P_13907_out0;
assign v$P19_16321_out0 = v$P_13979_out0;
assign v$G16_16449_out0 = v$G_10102_out0;
assign v$G16_16452_out0 = v$G_10174_out0;
assign v$G14_17977_out0 = v$G_10086_out0;
assign v$G14_17980_out0 = v$G_10158_out0;
assign v$GATE1_660_out0 = v$GATE2_15757_out0 || v$G0_15943_out0;
assign v$GATE1_663_out0 = v$GATE2_15760_out0 || v$G0_15946_out0;
assign v$P$AD_772_out0 = v$G1_5607_out0;
assign v$P$AD_781_out0 = v$G1_5616_out0;
assign v$P$AD_782_out0 = v$G1_5617_out0;
assign v$P$AD_793_out0 = v$G1_5628_out0;
assign v$P$AD_795_out0 = v$G1_5630_out0;
assign v$P$AD_802_out0 = v$G1_5637_out0;
assign v$P$AD_803_out0 = v$G1_5638_out0;
assign v$G$CD_956_out0 = v$G14_17977_out0;
assign v$G$CD_957_out0 = v$G8_2578_out0;
assign v$G$CD_959_out0 = v$G1_5054_out0;
assign v$G$CD_962_out0 = v$G19_1882_out0;
assign v$G$CD_963_out0 = v$G22_12511_out0;
assign v$G$CD_970_out0 = v$G23_14318_out0;
assign v$G$CD_972_out0 = v$G2_15961_out0;
assign v$G$CD_973_out0 = v$G5_10677_out0;
assign v$G$CD_975_out0 = v$G13_2829_out0;
assign v$G$CD_976_out0 = v$G17_9347_out0;
assign v$G$CD_977_out0 = v$G16_16449_out0;
assign v$G$CD_980_out0 = v$G7_1692_out0;
assign v$G$CD_986_out0 = v$G4_5736_out0;
assign v$G$CD_990_out0 = v$G20_8226_out0;
assign v$G$CD_991_out0 = v$G10_1834_out0;
assign v$G$CD_995_out0 = v$G11_11064_out0;
assign v$G$CD_1079_out0 = v$G14_17980_out0;
assign v$G$CD_1080_out0 = v$G8_2581_out0;
assign v$G$CD_1082_out0 = v$G1_5057_out0;
assign v$G$CD_1085_out0 = v$G19_1885_out0;
assign v$G$CD_1086_out0 = v$G22_12514_out0;
assign v$G$CD_1093_out0 = v$G23_14321_out0;
assign v$G$CD_1095_out0 = v$G2_15964_out0;
assign v$G$CD_1096_out0 = v$G5_10680_out0;
assign v$G$CD_1098_out0 = v$G13_2832_out0;
assign v$G$CD_1099_out0 = v$G17_9350_out0;
assign v$G$CD_1100_out0 = v$G16_16452_out0;
assign v$G$CD_1103_out0 = v$G7_1695_out0;
assign v$G$CD_1109_out0 = v$G4_5739_out0;
assign v$G$CD_1113_out0 = v$G20_8229_out0;
assign v$G$CD_1114_out0 = v$G10_1837_out0;
assign v$G$CD_1118_out0 = v$G11_11067_out0;
assign v$SUM_3476_out0 = v$SUM_15176_out0;
assign v$COUTD_6775_out0 = v$G6_515_out0;
assign v$COUTD_6780_out0 = v$G6_520_out0;
assign v$COUTD_6786_out0 = v$G6_526_out0;
assign v$COUTD_6789_out0 = v$G6_529_out0;
assign v$COUTD_6794_out0 = v$G6_534_out0;
assign v$COUTD_6807_out0 = v$G6_547_out0;
assign v$P$CD_10496_out0 = v$P14_3152_out0;
assign v$P$CD_10497_out0 = v$P8_1704_out0;
assign v$P$CD_10499_out0 = v$P1_2960_out0;
assign v$P$CD_10502_out0 = v$P19_16318_out0;
assign v$P$CD_10503_out0 = v$P22_4735_out0;
assign v$P$CD_10510_out0 = v$P23_6387_out0;
assign v$P$CD_10512_out0 = v$P2_2220_out0;
assign v$P$CD_10513_out0 = v$P5_222_out0;
assign v$P$CD_10515_out0 = v$P13_3033_out0;
assign v$P$CD_10516_out0 = v$P17_11760_out0;
assign v$P$CD_10517_out0 = v$P16_6963_out0;
assign v$P$CD_10520_out0 = v$P7_11770_out0;
assign v$P$CD_10526_out0 = v$P4_13637_out0;
assign v$P$CD_10530_out0 = v$P20_10660_out0;
assign v$P$CD_10531_out0 = v$P10_345_out0;
assign v$P$CD_10535_out0 = v$P11_9612_out0;
assign v$P$CD_10619_out0 = v$P14_3155_out0;
assign v$P$CD_10620_out0 = v$P8_1707_out0;
assign v$P$CD_10622_out0 = v$P1_2963_out0;
assign v$P$CD_10625_out0 = v$P19_16321_out0;
assign v$P$CD_10626_out0 = v$P22_4738_out0;
assign v$P$CD_10633_out0 = v$P23_6390_out0;
assign v$P$CD_10635_out0 = v$P2_2223_out0;
assign v$P$CD_10636_out0 = v$P5_225_out0;
assign v$P$CD_10638_out0 = v$P13_3036_out0;
assign v$P$CD_10639_out0 = v$P17_11763_out0;
assign v$P$CD_10640_out0 = v$P16_6966_out0;
assign v$P$CD_10643_out0 = v$P7_11773_out0;
assign v$P$CD_10649_out0 = v$P4_13640_out0;
assign v$P$CD_10653_out0 = v$P20_10663_out0;
assign v$P$CD_10654_out0 = v$P10_348_out0;
assign v$P$CD_10658_out0 = v$P11_9615_out0;
assign v$COUT_10738_out0 = v$COUT_8121_out0;
assign v$G4_11199_out0 = v$G5_4607_out0 || v$G$CD_1002_out0;
assign v$G4_11203_out0 = v$G5_4611_out0 || v$G$CD_1006_out0;
assign v$G4_11222_out0 = v$G5_4630_out0 || v$G$CD_1025_out0;
assign v$G4_11230_out0 = v$G5_4638_out0 || v$G$CD_1033_out0;
assign v$G4_11232_out0 = v$G5_4640_out0 || v$G$CD_1035_out0;
assign v$G8_11440_out0 = v$CINA_8509_out0 && v$P$AB_2046_out0;
assign v$G8_11443_out0 = v$CINA_8512_out0 && v$P$AB_2049_out0;
assign v$G8_11444_out0 = v$CINA_8513_out0 && v$P$AB_2050_out0;
assign v$G8_11456_out0 = v$CINA_8525_out0 && v$P$AB_2062_out0;
assign v$G8_11458_out0 = v$CINA_8527_out0 && v$P$AB_2064_out0;
assign v$G8_11461_out0 = v$CINA_8530_out0 && v$P$AB_2067_out0;
assign v$G8_11467_out0 = v$CINA_8536_out0 && v$P$AB_2073_out0;
assign v$G8_11472_out0 = v$CINA_8541_out0 && v$P$AB_2078_out0;
assign v$G8_11563_out0 = v$CINA_8632_out0 && v$P$AB_2169_out0;
assign v$G8_11566_out0 = v$CINA_8635_out0 && v$P$AB_2172_out0;
assign v$G8_11567_out0 = v$CINA_8636_out0 && v$P$AB_2173_out0;
assign v$G8_11579_out0 = v$CINA_8648_out0 && v$P$AB_2185_out0;
assign v$G8_11581_out0 = v$CINA_8650_out0 && v$P$AB_2187_out0;
assign v$G8_11584_out0 = v$CINA_8653_out0 && v$P$AB_2190_out0;
assign v$G8_11590_out0 = v$CINA_8659_out0 && v$P$AB_2196_out0;
assign v$G8_11595_out0 = v$CINA_8664_out0 && v$P$AB_2201_out0;
assign v$SEL4_1186_out0 = v$SUM_3476_out0[0:0];
assign v$C4_1261_out0 = v$COUTD_6780_out0;
assign v$P$AB_2099_out0 = v$P$AD_772_out0;
assign v$P$AB_2106_out0 = v$P$AD_772_out0;
assign v$P$AB_2110_out0 = v$P$AD_793_out0;
assign v$P$AB_2113_out0 = v$P$AD_793_out0;
assign v$P$AB_2121_out0 = v$P$AD_772_out0;
assign v$END27_2212_out0 = v$P$AD_802_out0;
assign v$CIN_3897_out0 = v$COUT_10738_out0;
assign v$END21_4342_out0 = v$P$AD_782_out0;
assign v$G5_4564_out0 = v$G$AB_9181_out0 && v$P$CD_10499_out0;
assign v$G5_4567_out0 = v$G$AB_9184_out0 && v$P$CD_10502_out0;
assign v$G5_4568_out0 = v$G$AB_9185_out0 && v$P$CD_10503_out0;
assign v$G5_4580_out0 = v$G$AB_9197_out0 && v$P$CD_10515_out0;
assign v$G5_4582_out0 = v$G$AB_9199_out0 && v$P$CD_10517_out0;
assign v$G5_4585_out0 = v$G$AB_9202_out0 && v$P$CD_10520_out0;
assign v$G5_4591_out0 = v$G$AB_9208_out0 && v$P$CD_10526_out0;
assign v$G5_4596_out0 = v$G$AB_9213_out0 && v$P$CD_10531_out0;
assign v$G5_4687_out0 = v$G$AB_9304_out0 && v$P$CD_10622_out0;
assign v$G5_4690_out0 = v$G$AB_9307_out0 && v$P$CD_10625_out0;
assign v$G5_4691_out0 = v$G$AB_9308_out0 && v$P$CD_10626_out0;
assign v$G5_4703_out0 = v$G$AB_9320_out0 && v$P$CD_10638_out0;
assign v$G5_4705_out0 = v$G$AB_9322_out0 && v$P$CD_10640_out0;
assign v$G5_4708_out0 = v$G$AB_9325_out0 && v$P$CD_10643_out0;
assign v$G5_4714_out0 = v$G$AB_9331_out0 && v$P$CD_10649_out0;
assign v$G5_4719_out0 = v$G$AB_9336_out0 && v$P$CD_10654_out0;
assign v$G1_5567_out0 = v$P$AB_2046_out0 && v$P$CD_10499_out0;
assign v$G1_5570_out0 = v$P$AB_2049_out0 && v$P$CD_10502_out0;
assign v$G1_5571_out0 = v$P$AB_2050_out0 && v$P$CD_10503_out0;
assign v$G1_5583_out0 = v$P$AB_2062_out0 && v$P$CD_10515_out0;
assign v$G1_5585_out0 = v$P$AB_2064_out0 && v$P$CD_10517_out0;
assign v$G1_5588_out0 = v$P$AB_2067_out0 && v$P$CD_10520_out0;
assign v$G1_5594_out0 = v$P$AB_2073_out0 && v$P$CD_10526_out0;
assign v$G1_5599_out0 = v$P$AB_2078_out0 && v$P$CD_10531_out0;
assign v$G1_5690_out0 = v$P$AB_2169_out0 && v$P$CD_10622_out0;
assign v$G1_5693_out0 = v$P$AB_2172_out0 && v$P$CD_10625_out0;
assign v$G1_5694_out0 = v$P$AB_2173_out0 && v$P$CD_10626_out0;
assign v$G1_5706_out0 = v$P$AB_2185_out0 && v$P$CD_10638_out0;
assign v$G1_5708_out0 = v$P$AB_2187_out0 && v$P$CD_10640_out0;
assign v$G1_5711_out0 = v$P$AB_2190_out0 && v$P$CD_10643_out0;
assign v$G1_5717_out0 = v$P$AB_2196_out0 && v$P$CD_10649_out0;
assign v$G1_5722_out0 = v$P$AB_2201_out0 && v$P$CD_10654_out0;
assign v$END40_5777_out0 = v$COUTD_6794_out0;
assign v$END29_5887_out0 = v$P$AD_793_out0;
assign v$CINA_8552_out0 = v$COUTD_6807_out0;
assign v$CINA_8556_out0 = v$COUTD_6807_out0;
assign v$CINA_8575_out0 = v$COUTD_6807_out0;
assign v$CINA_8583_out0 = v$COUTD_6794_out0;
assign v$CINA_8585_out0 = v$COUTD_6807_out0;
assign v$END4_9369_out0 = v$COUTD_6775_out0;
assign v$G7_9680_out0 = v$G8_11440_out0 && v$P$CD_10499_out0;
assign v$G7_9683_out0 = v$G8_11443_out0 && v$P$CD_10502_out0;
assign v$G7_9684_out0 = v$G8_11444_out0 && v$P$CD_10503_out0;
assign v$G7_9696_out0 = v$G8_11456_out0 && v$P$CD_10515_out0;
assign v$G7_9698_out0 = v$G8_11458_out0 && v$P$CD_10517_out0;
assign v$G7_9701_out0 = v$G8_11461_out0 && v$P$CD_10520_out0;
assign v$G7_9707_out0 = v$G8_11467_out0 && v$P$CD_10526_out0;
assign v$G7_9712_out0 = v$G8_11472_out0 && v$P$CD_10531_out0;
assign v$G7_9803_out0 = v$G8_11563_out0 && v$P$CD_10622_out0;
assign v$G7_9806_out0 = v$G8_11566_out0 && v$P$CD_10625_out0;
assign v$G7_9807_out0 = v$G8_11567_out0 && v$P$CD_10626_out0;
assign v$G7_9819_out0 = v$G8_11579_out0 && v$P$CD_10638_out0;
assign v$G7_9821_out0 = v$G8_11581_out0 && v$P$CD_10640_out0;
assign v$G7_9824_out0 = v$G8_11584_out0 && v$P$CD_10643_out0;
assign v$G7_9830_out0 = v$G8_11590_out0 && v$P$CD_10649_out0;
assign v$G7_9835_out0 = v$G8_11595_out0 && v$P$CD_10654_out0;
assign v$C0_10693_out0 = v$GATE1_660_out0;
assign v$C0_10696_out0 = v$GATE1_663_out0;
assign v$END52_11975_out0 = v$P$AD_795_out0;
assign v$OP1_14196_out0 = v$SUM_3476_out0;
assign v$END60_15134_out0 = v$COUTD_6789_out0;
assign v$C3_15728_out0 = v$COUTD_6786_out0;
assign v$C5_15917_out0 = v$COUTD_6807_out0;
assign v$END23_16719_out0 = v$P$AD_803_out0;
assign v$END25_17072_out0 = v$P$AD_781_out0;
assign v$G$AD_17174_out0 = v$G4_11199_out0;
assign v$G$AD_17178_out0 = v$G4_11203_out0;
assign v$G$AD_17197_out0 = v$G4_11222_out0;
assign v$G$AD_17205_out0 = v$G4_11230_out0;
assign v$G$AD_17207_out0 = v$G4_11232_out0;
assign v$END16_218_out0 = v$G$AD_17207_out0;
assign v$END14_276_out0 = v$G$AD_17178_out0;
assign v$P$AD_732_out0 = v$G1_5567_out0;
assign v$P$AD_735_out0 = v$G1_5570_out0;
assign v$P$AD_736_out0 = v$G1_5571_out0;
assign v$P$AD_748_out0 = v$G1_5583_out0;
assign v$P$AD_750_out0 = v$G1_5585_out0;
assign v$P$AD_753_out0 = v$G1_5588_out0;
assign v$P$AD_759_out0 = v$G1_5594_out0;
assign v$P$AD_764_out0 = v$G1_5599_out0;
assign v$P$AD_855_out0 = v$G1_5690_out0;
assign v$P$AD_858_out0 = v$G1_5693_out0;
assign v$P$AD_859_out0 = v$G1_5694_out0;
assign v$P$AD_871_out0 = v$G1_5706_out0;
assign v$P$AD_873_out0 = v$G1_5708_out0;
assign v$P$AD_876_out0 = v$G1_5711_out0;
assign v$P$AD_882_out0 = v$G1_5717_out0;
assign v$P$AD_887_out0 = v$G1_5722_out0;
assign v$G$CD_1022_out0 = v$G$AD_17205_out0;
assign {v$A2A_1632_out1,v$A2A_1632_out0 } = v$A1_1711_out0 + v$B1_8124_out0 + v$C0_10693_out0;
assign {v$A2A_1635_out1,v$A2A_1635_out0 } = v$A1_1714_out0 + v$B1_8127_out0 + v$C0_10696_out0;
assign {v$A7A_1659_out1,v$A7A_1659_out0 } = v$A5_6667_out0 + v$B5_18376_out0 + v$C4_1261_out0;
assign v$C4_1878_out0 = v$C4_1261_out0;
assign {v$A6A_3123_out1,v$A6A_3123_out0 } = v$A6_310_out0 + v$B6_13300_out0 + v$C5_15917_out0;
assign v$OP1_3390_out0 = v$OP1_14196_out0;
assign v$G1_5620_out0 = v$P$AB_2099_out0 && v$P$CD_10552_out0;
assign v$G1_5627_out0 = v$P$AB_2106_out0 && v$P$CD_10559_out0;
assign v$G1_5631_out0 = v$P$AB_2110_out0 && v$P$CD_10563_out0;
assign v$G1_5634_out0 = v$P$AB_2113_out0 && v$P$CD_10566_out0;
assign v$G1_5642_out0 = v$P$AB_2121_out0 && v$P$CD_10574_out0;
assign v$G$AB_9221_out0 = v$G$AD_17197_out0;
assign v$G$AB_9230_out0 = v$G$AD_17197_out0;
assign v$G$AB_9231_out0 = v$G$AD_17174_out0;
assign v$G$AB_9242_out0 = v$G$AD_17197_out0;
assign v$G$AB_9244_out0 = v$G$AD_17197_out0;
assign v$G$AB_9251_out0 = v$G$AD_17197_out0;
assign v$G$AB_9252_out0 = v$G$AD_17174_out0;
assign v$C0_9375_out0 = v$C0_10693_out0;
assign v$C0_9378_out0 = v$C0_10696_out0;
assign v$G4_11156_out0 = v$G5_4564_out0 || v$G$CD_959_out0;
assign v$G4_11159_out0 = v$G5_4567_out0 || v$G$CD_962_out0;
assign v$G4_11160_out0 = v$G5_4568_out0 || v$G$CD_963_out0;
assign v$G4_11172_out0 = v$G5_4580_out0 || v$G$CD_975_out0;
assign v$G4_11174_out0 = v$G5_4582_out0 || v$G$CD_977_out0;
assign v$G4_11177_out0 = v$G5_4585_out0 || v$G$CD_980_out0;
assign v$G4_11183_out0 = v$G5_4591_out0 || v$G$CD_986_out0;
assign v$G4_11188_out0 = v$G5_4596_out0 || v$G$CD_991_out0;
assign v$G4_11279_out0 = v$G5_4687_out0 || v$G$CD_1082_out0;
assign v$G4_11282_out0 = v$G5_4690_out0 || v$G$CD_1085_out0;
assign v$G4_11283_out0 = v$G5_4691_out0 || v$G$CD_1086_out0;
assign v$G4_11295_out0 = v$G5_4703_out0 || v$G$CD_1098_out0;
assign v$G4_11297_out0 = v$G5_4705_out0 || v$G$CD_1100_out0;
assign v$G4_11300_out0 = v$G5_4708_out0 || v$G$CD_1103_out0;
assign v$G4_11306_out0 = v$G5_4714_out0 || v$G$CD_1109_out0;
assign v$G4_11311_out0 = v$G5_4719_out0 || v$G$CD_1114_out0;
assign v$G8_11483_out0 = v$CINA_8552_out0 && v$P$AB_2089_out0;
assign v$G8_11487_out0 = v$CINA_8556_out0 && v$P$AB_2093_out0;
assign v$G8_11506_out0 = v$CINA_8575_out0 && v$P$AB_2112_out0;
assign v$G8_11514_out0 = v$CINA_8583_out0 && v$P$AB_2120_out0;
assign v$G8_11516_out0 = v$CINA_8585_out0 && v$P$AB_2122_out0;
assign v$C5_11688_out0 = v$C5_15917_out0;
assign v$END18_11948_out0 = v$G$AD_17174_out0;
assign v$SUM$4_15246_out0 = v$SEL4_1186_out0;
assign v$C3_15819_out0 = v$C3_15728_out0;
assign {v$A5A_16101_out1,v$A5A_16101_out0 } = v$A4_17500_out0 + v$B4_14665_out0 + v$C3_15728_out0;
assign v$CIN_16823_out0 = v$CIN_3897_out0;
assign v$_84_out0 = { v$A5A_16101_out0,v$A7A_1659_out0 };
assign v$G6_478_out0 = v$G4_11156_out0 || v$G7_9680_out0;
assign v$G6_481_out0 = v$G4_11159_out0 || v$G7_9683_out0;
assign v$G6_482_out0 = v$G4_11160_out0 || v$G7_9684_out0;
assign v$G6_494_out0 = v$G4_11172_out0 || v$G7_9696_out0;
assign v$G6_496_out0 = v$G4_11174_out0 || v$G7_9698_out0;
assign v$G6_499_out0 = v$G4_11177_out0 || v$G7_9701_out0;
assign v$G6_505_out0 = v$G4_11183_out0 || v$G7_9707_out0;
assign v$G6_510_out0 = v$G4_11188_out0 || v$G7_9712_out0;
assign v$G6_601_out0 = v$G4_11279_out0 || v$G7_9803_out0;
assign v$G6_604_out0 = v$G4_11282_out0 || v$G7_9806_out0;
assign v$G6_605_out0 = v$G4_11283_out0 || v$G7_9807_out0;
assign v$G6_617_out0 = v$G4_11295_out0 || v$G7_9819_out0;
assign v$G6_619_out0 = v$G4_11297_out0 || v$G7_9821_out0;
assign v$G6_622_out0 = v$G4_11300_out0 || v$G7_9824_out0;
assign v$G6_628_out0 = v$G4_11306_out0 || v$G7_9830_out0;
assign v$G6_633_out0 = v$G4_11311_out0 || v$G7_9835_out0;
assign v$P$AD_785_out0 = v$G1_5620_out0;
assign v$P$AD_792_out0 = v$G1_5627_out0;
assign v$P$AD_796_out0 = v$G1_5631_out0;
assign v$P$AD_799_out0 = v$G1_5634_out0;
assign v$P$AD_807_out0 = v$G1_5642_out0;
assign v$END1_1544_out0 = v$A2A_1632_out1;
assign v$END1_1547_out0 = v$A2A_1635_out1;
assign v$P$AB_2043_out0 = v$P$AD_748_out0;
assign v$P$AB_2044_out0 = v$P$AD_753_out0;
assign v$P$AB_2057_out0 = v$P$AD_736_out0;
assign v$P$AB_2059_out0 = v$P$AD_732_out0;
assign v$P$AB_2060_out0 = v$P$AD_759_out0;
assign v$P$AB_2063_out0 = v$P$AD_750_out0;
assign v$P$AB_2077_out0 = v$P$AD_735_out0;
assign v$P$AB_2082_out0 = v$P$AD_764_out0;
assign v$P$AB_2166_out0 = v$P$AD_871_out0;
assign v$P$AB_2167_out0 = v$P$AD_876_out0;
assign v$P$AB_2180_out0 = v$P$AD_859_out0;
assign v$P$AB_2182_out0 = v$P$AD_855_out0;
assign v$P$AB_2183_out0 = v$P$AD_882_out0;
assign v$P$AB_2186_out0 = v$P$AD_873_out0;
assign v$P$AB_2200_out0 = v$P$AD_858_out0;
assign v$P$AB_2205_out0 = v$P$AD_887_out0;
assign v$_2455_out0 = { v$C4_1878_out0,v$C5_11688_out0 };
assign v$END5_4145_out0 = v$A7A_1659_out1;
assign v$G5_4604_out0 = v$G$AB_9221_out0 && v$P$CD_10539_out0;
assign v$G5_4613_out0 = v$G$AB_9230_out0 && v$P$CD_10548_out0;
assign v$G5_4614_out0 = v$G$AB_9231_out0 && v$P$CD_10549_out0;
assign v$G5_4625_out0 = v$G$AB_9242_out0 && v$P$CD_10560_out0;
assign v$G5_4627_out0 = v$G$AB_9244_out0 && v$P$CD_10562_out0;
assign v$G5_4634_out0 = v$G$AB_9251_out0 && v$P$CD_10569_out0;
assign v$G5_4635_out0 = v$G$AB_9252_out0 && v$P$CD_10570_out0;
assign v$END4_5248_out0 = v$A5A_16101_out1;
assign v$G7_9723_out0 = v$G8_11483_out0 && v$P$CD_10542_out0;
assign v$G7_9727_out0 = v$G8_11487_out0 && v$P$CD_10546_out0;
assign v$G7_9746_out0 = v$G8_11506_out0 && v$P$CD_10565_out0;
assign v$G7_9754_out0 = v$G8_11514_out0 && v$P$CD_10573_out0;
assign v$G7_9756_out0 = v$G8_11516_out0 && v$P$CD_10575_out0;
assign v$P$CD_10500_out0 = v$P$AD_759_out0;
assign v$P$CD_10504_out0 = v$P$AD_736_out0;
assign v$P$CD_10525_out0 = v$P$AD_750_out0;
assign v$P$CD_10528_out0 = v$P$AD_748_out0;
assign v$P$CD_10529_out0 = v$P$AD_764_out0;
assign v$P$CD_10533_out0 = v$P$AD_735_out0;
assign v$P$CD_10534_out0 = v$P$AD_753_out0;
assign v$P$CD_10623_out0 = v$P$AD_882_out0;
assign v$P$CD_10627_out0 = v$P$AD_859_out0;
assign v$P$CD_10648_out0 = v$P$AD_873_out0;
assign v$P$CD_10651_out0 = v$P$AD_871_out0;
assign v$P$CD_10652_out0 = v$P$AD_887_out0;
assign v$P$CD_10656_out0 = v$P$AD_858_out0;
assign v$P$CD_10657_out0 = v$P$AD_876_out0;
assign v$_13438_out0 = { v$A1A_11661_out0,v$A2A_1632_out0 };
assign v$_13441_out0 = { v$A1A_11664_out0,v$A2A_1635_out0 };
assign v$_15000_out0 = { v$C2_18181_out0,v$C3_15819_out0 };
assign v$END6_15251_out0 = v$A6A_3123_out1;
assign v$G$AD_17131_out0 = v$G4_11156_out0;
assign v$G$AD_17134_out0 = v$G4_11159_out0;
assign v$G$AD_17135_out0 = v$G4_11160_out0;
assign v$G$AD_17147_out0 = v$G4_11172_out0;
assign v$G$AD_17149_out0 = v$G4_11174_out0;
assign v$G$AD_17152_out0 = v$G4_11177_out0;
assign v$G$AD_17158_out0 = v$G4_11183_out0;
assign v$G$AD_17163_out0 = v$G4_11188_out0;
assign v$G$AD_17254_out0 = v$G4_11279_out0;
assign v$G$AD_17257_out0 = v$G4_11282_out0;
assign v$G$AD_17258_out0 = v$G4_11283_out0;
assign v$G$AD_17270_out0 = v$G4_11295_out0;
assign v$G$AD_17272_out0 = v$G4_11297_out0;
assign v$G$AD_17275_out0 = v$G4_11300_out0;
assign v$G$AD_17281_out0 = v$G4_11306_out0;
assign v$G$AD_17286_out0 = v$G4_11311_out0;
assign v$SEL8_17662_out0 = v$OP1_3390_out0[23:1];
assign v$END33_266_out0 = v$P$AD_799_out0;
assign v$G6_521_out0 = v$G4_11199_out0 || v$G7_9723_out0;
assign v$G6_525_out0 = v$G4_11203_out0 || v$G7_9727_out0;
assign v$G6_544_out0 = v$G4_11222_out0 || v$G7_9746_out0;
assign v$G6_552_out0 = v$G4_11230_out0 || v$G7_9754_out0;
assign v$G6_554_out0 = v$G4_11232_out0 || v$G7_9756_out0;
assign v$G$CD_960_out0 = v$G$AD_17158_out0;
assign v$G$CD_964_out0 = v$G$AD_17135_out0;
assign v$G$CD_985_out0 = v$G$AD_17149_out0;
assign v$G$CD_988_out0 = v$G$AD_17147_out0;
assign v$G$CD_989_out0 = v$G$AD_17163_out0;
assign v$G$CD_993_out0 = v$G$AD_17134_out0;
assign v$G$CD_994_out0 = v$G$AD_17152_out0;
assign v$G$CD_1083_out0 = v$G$AD_17281_out0;
assign v$G$CD_1087_out0 = v$G$AD_17258_out0;
assign v$G$CD_1108_out0 = v$G$AD_17272_out0;
assign v$G$CD_1111_out0 = v$G$AD_17270_out0;
assign v$G$CD_1112_out0 = v$G$AD_17286_out0;
assign v$G$CD_1116_out0 = v$G$AD_17257_out0;
assign v$G$CD_1117_out0 = v$G$AD_17275_out0;
assign v$P$AB_2092_out0 = v$P$AD_792_out0;
assign v$P$AB_2111_out0 = v$P$AD_792_out0;
assign v$END47_2681_out0 = v$P$AD_792_out0;
assign v$G1_5564_out0 = v$P$AB_2043_out0 && v$P$CD_10496_out0;
assign v$G1_5565_out0 = v$P$AB_2044_out0 && v$P$CD_10497_out0;
assign v$G1_5578_out0 = v$P$AB_2057_out0 && v$P$CD_10510_out0;
assign v$G1_5580_out0 = v$P$AB_2059_out0 && v$P$CD_10512_out0;
assign v$G1_5581_out0 = v$P$AB_2060_out0 && v$P$CD_10513_out0;
assign v$G1_5584_out0 = v$P$AB_2063_out0 && v$P$CD_10516_out0;
assign v$G1_5598_out0 = v$P$AB_2077_out0 && v$P$CD_10530_out0;
assign v$G1_5603_out0 = v$P$AB_2082_out0 && v$P$CD_10535_out0;
assign v$G1_5687_out0 = v$P$AB_2166_out0 && v$P$CD_10619_out0;
assign v$G1_5688_out0 = v$P$AB_2167_out0 && v$P$CD_10620_out0;
assign v$G1_5701_out0 = v$P$AB_2180_out0 && v$P$CD_10633_out0;
assign v$G1_5703_out0 = v$P$AB_2182_out0 && v$P$CD_10635_out0;
assign v$G1_5704_out0 = v$P$AB_2183_out0 && v$P$CD_10636_out0;
assign v$G1_5707_out0 = v$P$AB_2186_out0 && v$P$CD_10639_out0;
assign v$G1_5721_out0 = v$P$AB_2200_out0 && v$P$CD_10653_out0;
assign v$G1_5726_out0 = v$P$AB_2205_out0 && v$P$CD_10658_out0;
assign v$COUTD_6738_out0 = v$G6_478_out0;
assign v$COUTD_6741_out0 = v$G6_481_out0;
assign v$COUTD_6742_out0 = v$G6_482_out0;
assign v$COUTD_6754_out0 = v$G6_494_out0;
assign v$COUTD_6756_out0 = v$G6_496_out0;
assign v$COUTD_6759_out0 = v$G6_499_out0;
assign v$COUTD_6765_out0 = v$G6_505_out0;
assign v$COUTD_6770_out0 = v$G6_510_out0;
assign v$COUTD_6861_out0 = v$G6_601_out0;
assign v$COUTD_6864_out0 = v$G6_604_out0;
assign v$COUTD_6865_out0 = v$G6_605_out0;
assign v$COUTD_6877_out0 = v$G6_617_out0;
assign v$COUTD_6879_out0 = v$G6_619_out0;
assign v$COUTD_6882_out0 = v$G6_622_out0;
assign v$COUTD_6888_out0 = v$G6_628_out0;
assign v$COUTD_6893_out0 = v$G6_633_out0;
assign v$_7255_out0 = { v$_8908_out0,v$_15000_out0 };
assign v$G$AB_9178_out0 = v$G$AD_17147_out0;
assign v$G$AB_9179_out0 = v$G$AD_17152_out0;
assign v$G$AB_9192_out0 = v$G$AD_17135_out0;
assign v$G$AB_9194_out0 = v$G$AD_17131_out0;
assign v$G$AB_9195_out0 = v$G$AD_17158_out0;
assign v$G$AB_9198_out0 = v$G$AD_17149_out0;
assign v$G$AB_9212_out0 = v$G$AD_17134_out0;
assign v$G$AB_9217_out0 = v$G$AD_17163_out0;
assign v$G$AB_9301_out0 = v$G$AD_17270_out0;
assign v$G$AB_9302_out0 = v$G$AD_17275_out0;
assign v$G$AB_9315_out0 = v$G$AD_17258_out0;
assign v$G$AB_9317_out0 = v$G$AD_17254_out0;
assign v$G$AB_9318_out0 = v$G$AD_17281_out0;
assign v$G$AB_9321_out0 = v$G$AD_17272_out0;
assign v$G$AB_9335_out0 = v$G$AD_17257_out0;
assign v$G$AB_9340_out0 = v$G$AD_17286_out0;
assign v$G4_11196_out0 = v$G5_4604_out0 || v$G$CD_999_out0;
assign v$G4_11205_out0 = v$G5_4613_out0 || v$G$CD_1008_out0;
assign v$G4_11206_out0 = v$G5_4614_out0 || v$G$CD_1009_out0;
assign v$G4_11217_out0 = v$G5_4625_out0 || v$G$CD_1020_out0;
assign v$G4_11219_out0 = v$G5_4627_out0 || v$G$CD_1022_out0;
assign v$G4_11226_out0 = v$G5_4634_out0 || v$G$CD_1029_out0;
assign v$G4_11227_out0 = v$G5_4635_out0 || v$G$CD_1030_out0;
assign v$END44_15667_out0 = v$P$AD_807_out0;
assign v$_18004_out0 = { v$SEL8_17662_out0,v$CIN_16823_out0 };
assign v$END42_18313_out0 = v$P$AD_785_out0;
assign v$END31_18522_out0 = v$P$AD_796_out0;
assign v$P$AD_729_out0 = v$G1_5564_out0;
assign v$P$AD_730_out0 = v$G1_5565_out0;
assign v$P$AD_743_out0 = v$G1_5578_out0;
assign v$P$AD_745_out0 = v$G1_5580_out0;
assign v$P$AD_746_out0 = v$G1_5581_out0;
assign v$P$AD_749_out0 = v$G1_5584_out0;
assign v$P$AD_763_out0 = v$G1_5598_out0;
assign v$P$AD_768_out0 = v$G1_5603_out0;
assign v$P$AD_852_out0 = v$G1_5687_out0;
assign v$P$AD_853_out0 = v$G1_5688_out0;
assign v$P$AD_866_out0 = v$G1_5701_out0;
assign v$P$AD_868_out0 = v$G1_5703_out0;
assign v$P$AD_869_out0 = v$G1_5704_out0;
assign v$P$AD_872_out0 = v$G1_5707_out0;
assign v$P$AD_886_out0 = v$G1_5721_out0;
assign v$P$AD_891_out0 = v$G1_5726_out0;
assign v$G5_4561_out0 = v$G$AB_9178_out0 && v$P$CD_10496_out0;
assign v$G5_4562_out0 = v$G$AB_9179_out0 && v$P$CD_10497_out0;
assign v$G5_4575_out0 = v$G$AB_9192_out0 && v$P$CD_10510_out0;
assign v$G5_4577_out0 = v$G$AB_9194_out0 && v$P$CD_10512_out0;
assign v$G5_4578_out0 = v$G$AB_9195_out0 && v$P$CD_10513_out0;
assign v$G5_4581_out0 = v$G$AB_9198_out0 && v$P$CD_10516_out0;
assign v$G5_4595_out0 = v$G$AB_9212_out0 && v$P$CD_10530_out0;
assign v$G5_4600_out0 = v$G$AB_9217_out0 && v$P$CD_10535_out0;
assign v$G5_4684_out0 = v$G$AB_9301_out0 && v$P$CD_10619_out0;
assign v$G5_4685_out0 = v$G$AB_9302_out0 && v$P$CD_10620_out0;
assign v$G5_4698_out0 = v$G$AB_9315_out0 && v$P$CD_10633_out0;
assign v$G5_4700_out0 = v$G$AB_9317_out0 && v$P$CD_10635_out0;
assign v$G5_4701_out0 = v$G$AB_9318_out0 && v$P$CD_10636_out0;
assign v$G5_4704_out0 = v$G$AB_9321_out0 && v$P$CD_10639_out0;
assign v$G5_4718_out0 = v$G$AB_9335_out0 && v$P$CD_10653_out0;
assign v$G5_4723_out0 = v$G$AB_9340_out0 && v$P$CD_10658_out0;
assign v$G1_5613_out0 = v$P$AB_2092_out0 && v$P$CD_10545_out0;
assign v$G1_5632_out0 = v$P$AB_2111_out0 && v$P$CD_10564_out0;
assign v$COUTD_6781_out0 = v$G6_521_out0;
assign v$COUTD_6785_out0 = v$G6_525_out0;
assign v$COUTD_6804_out0 = v$G6_544_out0;
assign v$COUTD_6812_out0 = v$G6_552_out0;
assign v$COUTD_6814_out0 = v$G6_554_out0;
assign v$CINA_8506_out0 = v$COUTD_6754_out0;
assign v$CINA_8507_out0 = v$COUTD_6759_out0;
assign v$CINA_8520_out0 = v$COUTD_6742_out0;
assign v$CINA_8522_out0 = v$COUTD_6738_out0;
assign v$CINA_8523_out0 = v$COUTD_6765_out0;
assign v$CINA_8526_out0 = v$COUTD_6756_out0;
assign v$CINA_8540_out0 = v$COUTD_6741_out0;
assign v$CINA_8545_out0 = v$COUTD_6770_out0;
assign v$CINA_8629_out0 = v$COUTD_6877_out0;
assign v$CINA_8630_out0 = v$COUTD_6882_out0;
assign v$CINA_8643_out0 = v$COUTD_6865_out0;
assign v$CINA_8645_out0 = v$COUTD_6861_out0;
assign v$CINA_8646_out0 = v$COUTD_6888_out0;
assign v$CINA_8649_out0 = v$COUTD_6879_out0;
assign v$CINA_8663_out0 = v$COUTD_6864_out0;
assign v$CINA_8668_out0 = v$COUTD_6893_out0;
assign {v$A1_15225_out1,v$A1_15225_out0 } = v$_18004_out0 + v$MUX1_8349_out0 + v$C6_11361_out0;
assign v$C1_16782_out0 = v$COUTD_6738_out0;
assign v$C1_16785_out0 = v$COUTD_6861_out0;
assign v$G$AD_17171_out0 = v$G4_11196_out0;
assign v$G$AD_17180_out0 = v$G4_11205_out0;
assign v$G$AD_17181_out0 = v$G4_11206_out0;
assign v$G$AD_17192_out0 = v$G4_11217_out0;
assign v$G$AD_17194_out0 = v$G4_11219_out0;
assign v$G$AD_17201_out0 = v$G4_11226_out0;
assign v$G$AD_17202_out0 = v$G4_11227_out0;
assign v$END53_319_out0 = v$G$AD_17194_out0;
assign v$P$AD_778_out0 = v$G1_5613_out0;
assign v$P$AD_797_out0 = v$G1_5632_out0;
assign v$P$AB_2042_out0 = v$P$AD_730_out0;
assign v$P$AB_2047_out0 = v$P$AD_745_out0;
assign v$P$AB_2053_out0 = v$P$AD_745_out0;
assign v$P$AB_2056_out0 = v$P$AD_763_out0;
assign v$P$AB_2061_out0 = v$P$AD_729_out0;
assign v$P$AB_2074_out0 = v$P$AD_745_out0;
assign v$P$AB_2165_out0 = v$P$AD_853_out0;
assign v$P$AB_2170_out0 = v$P$AD_868_out0;
assign v$P$AB_2176_out0 = v$P$AD_868_out0;
assign v$P$AB_2179_out0 = v$P$AD_886_out0;
assign v$P$AB_2184_out0 = v$P$AD_852_out0;
assign v$P$AB_2197_out0 = v$P$AD_868_out0;
assign v$END26_6437_out0 = v$G$AD_17201_out0;
assign v$C8_7432_out0 = v$COUTD_6781_out0;
assign v$COUT_8122_out0 = v$A1_15225_out1;
assign v$CINA_8549_out0 = v$COUTD_6804_out0;
assign v$CINA_8558_out0 = v$COUTD_6804_out0;
assign v$CINA_8559_out0 = v$COUTD_6781_out0;
assign v$CINA_8570_out0 = v$COUTD_6804_out0;
assign v$CINA_8572_out0 = v$COUTD_6804_out0;
assign v$CINA_8579_out0 = v$COUTD_6804_out0;
assign v$CINA_8580_out0 = v$COUTD_6781_out0;
assign v$G$AB_9234_out0 = v$G$AD_17171_out0;
assign v$G$AB_9241_out0 = v$G$AD_17171_out0;
assign v$G$AB_9245_out0 = v$G$AD_17192_out0;
assign v$G$AB_9248_out0 = v$G$AD_17192_out0;
assign v$G$AB_9256_out0 = v$G$AD_17171_out0;
assign v$C6_9588_out0 = v$COUTD_6785_out0;
assign v$P$CD_10495_out0 = v$P$AD_768_out0;
assign v$P$CD_10501_out0 = v$P$AD_730_out0;
assign v$P$CD_10509_out0 = v$P$AD_743_out0;
assign v$P$CD_10514_out0 = v$P$AD_749_out0;
assign v$P$CD_10518_out0 = v$P$AD_763_out0;
assign v$P$CD_10519_out0 = v$P$AD_729_out0;
assign v$P$CD_10527_out0 = v$P$AD_746_out0;
assign v$P$CD_10618_out0 = v$P$AD_891_out0;
assign v$P$CD_10624_out0 = v$P$AD_853_out0;
assign v$P$CD_10632_out0 = v$P$AD_866_out0;
assign v$P$CD_10637_out0 = v$P$AD_872_out0;
assign v$P$CD_10641_out0 = v$P$AD_886_out0;
assign v$P$CD_10642_out0 = v$P$AD_852_out0;
assign v$P$CD_10650_out0 = v$P$AD_869_out0;
assign v$C7_10971_out0 = v$COUTD_6814_out0;
assign v$G4_11153_out0 = v$G5_4561_out0 || v$G$CD_956_out0;
assign v$G4_11154_out0 = v$G5_4562_out0 || v$G$CD_957_out0;
assign v$G4_11167_out0 = v$G5_4575_out0 || v$G$CD_970_out0;
assign v$G4_11169_out0 = v$G5_4577_out0 || v$G$CD_972_out0;
assign v$G4_11170_out0 = v$G5_4578_out0 || v$G$CD_973_out0;
assign v$G4_11173_out0 = v$G5_4581_out0 || v$G$CD_976_out0;
assign v$G4_11187_out0 = v$G5_4595_out0 || v$G$CD_990_out0;
assign v$G4_11192_out0 = v$G5_4600_out0 || v$G$CD_995_out0;
assign v$G4_11276_out0 = v$G5_4684_out0 || v$G$CD_1079_out0;
assign v$G4_11277_out0 = v$G5_4685_out0 || v$G$CD_1080_out0;
assign v$G4_11290_out0 = v$G5_4698_out0 || v$G$CD_1093_out0;
assign v$G4_11292_out0 = v$G5_4700_out0 || v$G$CD_1095_out0;
assign v$G4_11293_out0 = v$G5_4701_out0 || v$G$CD_1096_out0;
assign v$G4_11296_out0 = v$G5_4704_out0 || v$G$CD_1099_out0;
assign v$G4_11310_out0 = v$G5_4718_out0 || v$G$CD_1113_out0;
assign v$G4_11315_out0 = v$G5_4723_out0 || v$G$CD_1118_out0;
assign v$G8_11437_out0 = v$CINA_8506_out0 && v$P$AB_2043_out0;
assign v$G8_11438_out0 = v$CINA_8507_out0 && v$P$AB_2044_out0;
assign v$G8_11451_out0 = v$CINA_8520_out0 && v$P$AB_2057_out0;
assign v$G8_11453_out0 = v$CINA_8522_out0 && v$P$AB_2059_out0;
assign v$G8_11454_out0 = v$CINA_8523_out0 && v$P$AB_2060_out0;
assign v$G8_11457_out0 = v$CINA_8526_out0 && v$P$AB_2063_out0;
assign v$G8_11471_out0 = v$CINA_8540_out0 && v$P$AB_2077_out0;
assign v$G8_11476_out0 = v$CINA_8545_out0 && v$P$AB_2082_out0;
assign v$G8_11560_out0 = v$CINA_8629_out0 && v$P$AB_2166_out0;
assign v$G8_11561_out0 = v$CINA_8630_out0 && v$P$AB_2167_out0;
assign v$G8_11574_out0 = v$CINA_8643_out0 && v$P$AB_2180_out0;
assign v$G8_11576_out0 = v$CINA_8645_out0 && v$P$AB_2182_out0;
assign v$G8_11577_out0 = v$CINA_8646_out0 && v$P$AB_2183_out0;
assign v$G8_11580_out0 = v$CINA_8649_out0 && v$P$AB_2186_out0;
assign v$G8_11594_out0 = v$CINA_8663_out0 && v$P$AB_2200_out0;
assign v$G8_11599_out0 = v$CINA_8668_out0 && v$P$AB_2205_out0;
assign v$C1_11850_out0 = v$C1_16782_out0;
assign v$C1_11853_out0 = v$C1_16785_out0;
assign {v$A3A_11952_out1,v$A3A_11952_out0 } = v$A2_18267_out0 + v$B2_3114_out0 + v$C1_16782_out0;
assign {v$A3A_11955_out1,v$A3A_11955_out0 } = v$A2_18270_out0 + v$B2_3117_out0 + v$C1_16785_out0;
assign v$END20_13266_out0 = v$G$AD_17181_out0;
assign v$END28_13671_out0 = v$G$AD_17192_out0;
assign v$C11_14798_out0 = v$COUTD_6804_out0;
assign v$SUM_15177_out0 = v$A1_15225_out0;
assign v$END22_15486_out0 = v$G$AD_17202_out0;
assign v$END24_16405_out0 = v$G$AD_17180_out0;
assign v$END61_17958_out0 = v$COUTD_6812_out0;
assign {v$A8A_1507_out1,v$A8A_1507_out0 } = v$A7_15309_out0 + v$B7_17042_out0 + v$C6_9588_out0;
assign {v$A17A_2489_out1,v$A17A_2489_out0 } = v$A12_3140_out0 + v$B12_1952_out0 + v$C11_14798_out0;
assign v$SUM_3477_out0 = v$SUM_15177_out0;
assign v$G5_4617_out0 = v$G$AB_9234_out0 && v$P$CD_10552_out0;
assign v$G5_4624_out0 = v$G$AB_9241_out0 && v$P$CD_10559_out0;
assign v$G5_4628_out0 = v$G$AB_9245_out0 && v$P$CD_10563_out0;
assign v$G5_4631_out0 = v$G$AB_9248_out0 && v$P$CD_10566_out0;
assign v$G5_4639_out0 = v$G$AB_9256_out0 && v$P$CD_10574_out0;
assign v$END2_5235_out0 = v$A3A_11952_out1;
assign v$END2_5238_out0 = v$A3A_11955_out1;
assign v$G1_5563_out0 = v$P$AB_2042_out0 && v$P$CD_10495_out0;
assign v$G1_5568_out0 = v$P$AB_2047_out0 && v$P$CD_10500_out0;
assign v$G1_5574_out0 = v$P$AB_2053_out0 && v$P$CD_10506_out0;
assign v$G1_5577_out0 = v$P$AB_2056_out0 && v$P$CD_10509_out0;
assign v$G1_5582_out0 = v$P$AB_2061_out0 && v$P$CD_10514_out0;
assign v$G1_5595_out0 = v$P$AB_2074_out0 && v$P$CD_10527_out0;
assign v$G1_5686_out0 = v$P$AB_2165_out0 && v$P$CD_10618_out0;
assign v$G1_5691_out0 = v$P$AB_2170_out0 && v$P$CD_10623_out0;
assign v$G1_5697_out0 = v$P$AB_2176_out0 && v$P$CD_10629_out0;
assign v$G1_5700_out0 = v$P$AB_2179_out0 && v$P$CD_10632_out0;
assign v$G1_5705_out0 = v$P$AB_2184_out0 && v$P$CD_10637_out0;
assign v$G1_5718_out0 = v$P$AB_2197_out0 && v$P$CD_10650_out0;
assign v$C6_7057_out0 = v$C6_9588_out0;
assign v$_8907_out0 = { v$C0_9375_out0,v$C1_11850_out0 };
assign v$_8910_out0 = { v$C0_9378_out0,v$C1_11853_out0 };
assign v$C11_9512_out0 = v$C11_14798_out0;
assign v$G7_9677_out0 = v$G8_11437_out0 && v$P$CD_10496_out0;
assign v$G7_9678_out0 = v$G8_11438_out0 && v$P$CD_10497_out0;
assign v$G7_9691_out0 = v$G8_11451_out0 && v$P$CD_10510_out0;
assign v$G7_9693_out0 = v$G8_11453_out0 && v$P$CD_10512_out0;
assign v$G7_9694_out0 = v$G8_11454_out0 && v$P$CD_10513_out0;
assign v$G7_9697_out0 = v$G8_11457_out0 && v$P$CD_10516_out0;
assign v$G7_9711_out0 = v$G8_11471_out0 && v$P$CD_10530_out0;
assign v$G7_9716_out0 = v$G8_11476_out0 && v$P$CD_10535_out0;
assign v$G7_9800_out0 = v$G8_11560_out0 && v$P$CD_10619_out0;
assign v$G7_9801_out0 = v$G8_11561_out0 && v$P$CD_10620_out0;
assign v$G7_9814_out0 = v$G8_11574_out0 && v$P$CD_10633_out0;
assign v$G7_9816_out0 = v$G8_11576_out0 && v$P$CD_10635_out0;
assign v$G7_9817_out0 = v$G8_11577_out0 && v$P$CD_10636_out0;
assign v$G7_9820_out0 = v$G8_11580_out0 && v$P$CD_10639_out0;
assign v$G7_9834_out0 = v$G8_11594_out0 && v$P$CD_10653_out0;
assign v$G7_9839_out0 = v$G8_11599_out0 && v$P$CD_10658_out0;
assign {v$A9A_10413_out1,v$A9A_10413_out0 } = v$A8_18092_out0 + v$B8_13140_out0 + v$C7_10971_out0;
assign v$COUT_10739_out0 = v$COUT_8122_out0;
assign v$G8_11480_out0 = v$CINA_8549_out0 && v$P$AB_2086_out0;
assign v$G8_11489_out0 = v$CINA_8558_out0 && v$P$AB_2095_out0;
assign v$G8_11490_out0 = v$CINA_8559_out0 && v$P$AB_2096_out0;
assign v$G8_11501_out0 = v$CINA_8570_out0 && v$P$AB_2107_out0;
assign v$G8_11503_out0 = v$CINA_8572_out0 && v$P$AB_2109_out0;
assign v$G8_11510_out0 = v$CINA_8579_out0 && v$P$AB_2116_out0;
assign v$G8_11511_out0 = v$CINA_8580_out0 && v$P$AB_2117_out0;
assign v$END51_11678_out0 = v$P$AD_778_out0;
assign {v$A10A_16004_out1,v$A10A_16004_out0 } = v$A9_3437_out0 + v$B9_4067_out0 + v$C8_7432_out0;
assign v$C7_16432_out0 = v$C7_10971_out0;
assign v$G$AD_17128_out0 = v$G4_11153_out0;
assign v$G$AD_17129_out0 = v$G4_11154_out0;
assign v$G$AD_17142_out0 = v$G4_11167_out0;
assign v$G$AD_17144_out0 = v$G4_11169_out0;
assign v$G$AD_17145_out0 = v$G4_11170_out0;
assign v$G$AD_17148_out0 = v$G4_11173_out0;
assign v$G$AD_17162_out0 = v$G4_11187_out0;
assign v$G$AD_17167_out0 = v$G4_11192_out0;
assign v$G$AD_17251_out0 = v$G4_11276_out0;
assign v$G$AD_17252_out0 = v$G4_11277_out0;
assign v$G$AD_17265_out0 = v$G4_11290_out0;
assign v$G$AD_17267_out0 = v$G4_11292_out0;
assign v$G$AD_17268_out0 = v$G4_11293_out0;
assign v$G$AD_17271_out0 = v$G4_11296_out0;
assign v$G$AD_17285_out0 = v$G4_11310_out0;
assign v$G$AD_17290_out0 = v$G4_11315_out0;
assign v$END49_18452_out0 = v$P$AD_797_out0;
assign v$C8_18499_out0 = v$C8_7432_out0;
assign v$G6_475_out0 = v$G4_11153_out0 || v$G7_9677_out0;
assign v$G6_476_out0 = v$G4_11154_out0 || v$G7_9678_out0;
assign v$G6_489_out0 = v$G4_11167_out0 || v$G7_9691_out0;
assign v$G6_491_out0 = v$G4_11169_out0 || v$G7_9693_out0;
assign v$G6_492_out0 = v$G4_11170_out0 || v$G7_9694_out0;
assign v$G6_495_out0 = v$G4_11173_out0 || v$G7_9697_out0;
assign v$G6_509_out0 = v$G4_11187_out0 || v$G7_9711_out0;
assign v$G6_514_out0 = v$G4_11192_out0 || v$G7_9716_out0;
assign v$G6_598_out0 = v$G4_11276_out0 || v$G7_9800_out0;
assign v$G6_599_out0 = v$G4_11277_out0 || v$G7_9801_out0;
assign v$G6_612_out0 = v$G4_11290_out0 || v$G7_9814_out0;
assign v$G6_614_out0 = v$G4_11292_out0 || v$G7_9816_out0;
assign v$G6_615_out0 = v$G4_11293_out0 || v$G7_9817_out0;
assign v$G6_618_out0 = v$G4_11296_out0 || v$G7_9820_out0;
assign v$G6_632_out0 = v$G4_11310_out0 || v$G7_9834_out0;
assign v$G6_637_out0 = v$G4_11315_out0 || v$G7_9839_out0;
assign v$P$AD_728_out0 = v$G1_5563_out0;
assign v$P$AD_733_out0 = v$G1_5568_out0;
assign v$P$AD_739_out0 = v$G1_5574_out0;
assign v$P$AD_742_out0 = v$G1_5577_out0;
assign v$P$AD_747_out0 = v$G1_5582_out0;
assign v$P$AD_760_out0 = v$G1_5595_out0;
assign v$P$AD_851_out0 = v$G1_5686_out0;
assign v$P$AD_856_out0 = v$G1_5691_out0;
assign v$P$AD_862_out0 = v$G1_5697_out0;
assign v$P$AD_865_out0 = v$G1_5700_out0;
assign v$P$AD_870_out0 = v$G1_5705_out0;
assign v$P$AD_883_out0 = v$G1_5718_out0;
assign v$G$CD_955_out0 = v$G$AD_17167_out0;
assign v$G$CD_961_out0 = v$G$AD_17129_out0;
assign v$G$CD_969_out0 = v$G$AD_17142_out0;
assign v$G$CD_974_out0 = v$G$AD_17148_out0;
assign v$G$CD_978_out0 = v$G$AD_17162_out0;
assign v$G$CD_979_out0 = v$G$AD_17128_out0;
assign v$G$CD_987_out0 = v$G$AD_17145_out0;
assign v$G$CD_1078_out0 = v$G$AD_17290_out0;
assign v$G$CD_1084_out0 = v$G$AD_17252_out0;
assign v$G$CD_1092_out0 = v$G$AD_17265_out0;
assign v$G$CD_1097_out0 = v$G$AD_17271_out0;
assign v$G$CD_1101_out0 = v$G$AD_17285_out0;
assign v$G$CD_1102_out0 = v$G$AD_17251_out0;
assign v$G$CD_1110_out0 = v$G$AD_17268_out0;
assign v$END7_3361_out0 = v$A8A_1507_out1;
assign v$_3638_out0 = { v$A6A_3123_out0,v$A8A_1507_out0 };
assign v$CIN_3894_out0 = v$COUT_10739_out0;
assign v$END8_3903_out0 = v$A9A_10413_out1;
assign v$END9_4235_out0 = v$A10A_16004_out1;
assign v$SEL9_5394_out0 = v$SUM_3477_out0[0:0];
assign v$G$AB_9177_out0 = v$G$AD_17129_out0;
assign v$G$AB_9182_out0 = v$G$AD_17144_out0;
assign v$G$AB_9188_out0 = v$G$AD_17144_out0;
assign v$G$AB_9191_out0 = v$G$AD_17162_out0;
assign v$G$AB_9196_out0 = v$G$AD_17128_out0;
assign v$G$AB_9209_out0 = v$G$AD_17144_out0;
assign v$G$AB_9300_out0 = v$G$AD_17252_out0;
assign v$G$AB_9305_out0 = v$G$AD_17267_out0;
assign v$G$AB_9311_out0 = v$G$AD_17267_out0;
assign v$G$AB_9314_out0 = v$G$AD_17285_out0;
assign v$G$AB_9319_out0 = v$G$AD_17251_out0;
assign v$G$AB_9332_out0 = v$G$AD_17267_out0;
assign v$ENDw_9553_out0 = v$A17A_2489_out1;
assign v$G7_9720_out0 = v$G8_11480_out0 && v$P$CD_10539_out0;
assign v$G7_9729_out0 = v$G8_11489_out0 && v$P$CD_10548_out0;
assign v$G7_9730_out0 = v$G8_11490_out0 && v$P$CD_10549_out0;
assign v$G7_9741_out0 = v$G8_11501_out0 && v$P$CD_10560_out0;
assign v$G7_9743_out0 = v$G8_11503_out0 && v$P$CD_10562_out0;
assign v$G7_9750_out0 = v$G8_11510_out0 && v$P$CD_10569_out0;
assign v$G7_9751_out0 = v$G8_11511_out0 && v$P$CD_10570_out0;
assign v$G4_11209_out0 = v$G5_4617_out0 || v$G$CD_1012_out0;
assign v$G4_11216_out0 = v$G5_4624_out0 || v$G$CD_1019_out0;
assign v$G4_11220_out0 = v$G5_4628_out0 || v$G$CD_1023_out0;
assign v$G4_11223_out0 = v$G5_4631_out0 || v$G$CD_1026_out0;
assign v$G4_11231_out0 = v$G5_4639_out0 || v$G$CD_1034_out0;
assign v$OP1_14193_out0 = v$SUM_3477_out0;
assign v$_15015_out0 = { v$A9A_10413_out0,v$A10A_16004_out0 };
assign v$_16312_out0 = { v$C6_7057_out0,v$C7_16432_out0 };
assign v$G6_518_out0 = v$G4_11196_out0 || v$G7_9720_out0;
assign v$G6_527_out0 = v$G4_11205_out0 || v$G7_9729_out0;
assign v$G6_528_out0 = v$G4_11206_out0 || v$G7_9730_out0;
assign v$G6_539_out0 = v$G4_11217_out0 || v$G7_9741_out0;
assign v$G6_541_out0 = v$G4_11219_out0 || v$G7_9743_out0;
assign v$G6_548_out0 = v$G4_11226_out0 || v$G7_9750_out0;
assign v$G6_549_out0 = v$G4_11227_out0 || v$G7_9751_out0;
assign v$P$AB_2048_out0 = v$P$AD_760_out0;
assign v$P$AB_2052_out0 = v$P$AD_760_out0;
assign v$P$AB_2071_out0 = v$P$AD_760_out0;
assign v$P$AB_2079_out0 = v$P$AD_747_out0;
assign v$P$AB_2081_out0 = v$P$AD_760_out0;
assign v$P$AB_2171_out0 = v$P$AD_883_out0;
assign v$P$AB_2175_out0 = v$P$AD_883_out0;
assign v$P$AB_2194_out0 = v$P$AD_883_out0;
assign v$P$AB_2202_out0 = v$P$AD_870_out0;
assign v$P$AB_2204_out0 = v$P$AD_883_out0;
assign v$OP1_3387_out0 = v$OP1_14193_out0;
assign v$G5_4560_out0 = v$G$AB_9177_out0 && v$P$CD_10495_out0;
assign v$G5_4565_out0 = v$G$AB_9182_out0 && v$P$CD_10500_out0;
assign v$G5_4571_out0 = v$G$AB_9188_out0 && v$P$CD_10506_out0;
assign v$G5_4574_out0 = v$G$AB_9191_out0 && v$P$CD_10509_out0;
assign v$G5_4579_out0 = v$G$AB_9196_out0 && v$P$CD_10514_out0;
assign v$G5_4592_out0 = v$G$AB_9209_out0 && v$P$CD_10527_out0;
assign v$G5_4683_out0 = v$G$AB_9300_out0 && v$P$CD_10618_out0;
assign v$G5_4688_out0 = v$G$AB_9305_out0 && v$P$CD_10623_out0;
assign v$G5_4694_out0 = v$G$AB_9311_out0 && v$P$CD_10629_out0;
assign v$G5_4697_out0 = v$G$AB_9314_out0 && v$P$CD_10632_out0;
assign v$G5_4702_out0 = v$G$AB_9319_out0 && v$P$CD_10637_out0;
assign v$G5_4715_out0 = v$G$AB_9332_out0 && v$P$CD_10650_out0;
assign v$COUTD_6735_out0 = v$G6_475_out0;
assign v$COUTD_6736_out0 = v$G6_476_out0;
assign v$COUTD_6749_out0 = v$G6_489_out0;
assign v$COUTD_6751_out0 = v$G6_491_out0;
assign v$COUTD_6752_out0 = v$G6_492_out0;
assign v$COUTD_6755_out0 = v$G6_495_out0;
assign v$COUTD_6769_out0 = v$G6_509_out0;
assign v$COUTD_6774_out0 = v$G6_514_out0;
assign v$COUTD_6858_out0 = v$G6_598_out0;
assign v$COUTD_6859_out0 = v$G6_599_out0;
assign v$COUTD_6872_out0 = v$G6_612_out0;
assign v$COUTD_6874_out0 = v$G6_614_out0;
assign v$COUTD_6875_out0 = v$G6_615_out0;
assign v$COUTD_6878_out0 = v$G6_618_out0;
assign v$COUTD_6892_out0 = v$G6_632_out0;
assign v$COUTD_6897_out0 = v$G6_637_out0;
assign v$_7406_out0 = { v$_2455_out0,v$_16312_out0 };
assign v$SUM$5_7817_out0 = v$SEL9_5394_out0;
assign v$P$CD_10498_out0 = v$P$AD_747_out0;
assign v$P$CD_10524_out0 = v$P$AD_728_out0;
assign v$P$CD_10532_out0 = v$P$AD_742_out0;
assign v$P$CD_10621_out0 = v$P$AD_870_out0;
assign v$P$CD_10647_out0 = v$P$AD_851_out0;
assign v$P$CD_10655_out0 = v$P$AD_865_out0;
assign v$END11_12091_out0 = v$P$AD_739_out0;
assign v$END11_12094_out0 = v$P$AD_862_out0;
assign v$CIN_16820_out0 = v$CIN_3894_out0;
assign v$G$AD_17184_out0 = v$G4_11209_out0;
assign v$G$AD_17191_out0 = v$G4_11216_out0;
assign v$G$AD_17195_out0 = v$G4_11220_out0;
assign v$G$AD_17198_out0 = v$G4_11223_out0;
assign v$G$AD_17206_out0 = v$G4_11231_out0;
assign v$_17966_out0 = { v$_84_out0,v$_3638_out0 };
assign v$END13_18068_out0 = v$P$AD_733_out0;
assign v$END13_18071_out0 = v$P$AD_856_out0;
assign v$END1_1292_out0 = v$COUTD_6774_out0;
assign v$END1_1295_out0 = v$COUTD_6897_out0;
assign v$END32_2472_out0 = v$G$AD_17198_out0;
assign v$C2_2687_out0 = v$COUTD_6751_out0;
assign v$C2_2690_out0 = v$COUTD_6874_out0;
assign v$END_3320_out0 = v$COUTD_6752_out0;
assign v$END_3323_out0 = v$COUTD_6875_out0;
assign v$END3_3446_out0 = v$COUTD_6749_out0;
assign v$END3_3449_out0 = v$COUTD_6872_out0;
assign v$G1_5569_out0 = v$P$AB_2048_out0 && v$P$CD_10501_out0;
assign v$G1_5573_out0 = v$P$AB_2052_out0 && v$P$CD_10505_out0;
assign v$G1_5592_out0 = v$P$AB_2071_out0 && v$P$CD_10524_out0;
assign v$G1_5600_out0 = v$P$AB_2079_out0 && v$P$CD_10532_out0;
assign v$G1_5602_out0 = v$P$AB_2081_out0 && v$P$CD_10534_out0;
assign v$G1_5692_out0 = v$P$AB_2171_out0 && v$P$CD_10624_out0;
assign v$G1_5696_out0 = v$P$AB_2175_out0 && v$P$CD_10628_out0;
assign v$G1_5715_out0 = v$P$AB_2194_out0 && v$P$CD_10647_out0;
assign v$G1_5723_out0 = v$P$AB_2202_out0 && v$P$CD_10655_out0;
assign v$G1_5725_out0 = v$P$AB_2204_out0 && v$P$CD_10657_out0;
assign v$COUTD_6778_out0 = v$G6_518_out0;
assign v$COUTD_6787_out0 = v$G6_527_out0;
assign v$COUTD_6788_out0 = v$G6_528_out0;
assign v$COUTD_6799_out0 = v$G6_539_out0;
assign v$COUTD_6801_out0 = v$G6_541_out0;
assign v$COUTD_6808_out0 = v$G6_548_out0;
assign v$COUTD_6809_out0 = v$G6_549_out0;
assign v$END2_7752_out0 = v$COUTD_6755_out0;
assign v$END2_7755_out0 = v$COUTD_6878_out0;
assign v$_7792_out0 = { v$_7255_out0,v$_7406_out0 };
assign v$CINA_8505_out0 = v$COUTD_6736_out0;
assign v$CINA_8510_out0 = v$COUTD_6751_out0;
assign v$CINA_8516_out0 = v$COUTD_6751_out0;
assign v$CINA_8519_out0 = v$COUTD_6769_out0;
assign v$CINA_8524_out0 = v$COUTD_6735_out0;
assign v$CINA_8537_out0 = v$COUTD_6751_out0;
assign v$CINA_8628_out0 = v$COUTD_6859_out0;
assign v$CINA_8633_out0 = v$COUTD_6874_out0;
assign v$CINA_8639_out0 = v$COUTD_6874_out0;
assign v$CINA_8642_out0 = v$COUTD_6892_out0;
assign v$CINA_8647_out0 = v$COUTD_6858_out0;
assign v$CINA_8660_out0 = v$COUTD_6874_out0;
assign v$END45_9058_out0 = v$COUTD_6769_out0;
assign v$END45_9061_out0 = v$COUTD_6892_out0;
assign v$G$AB_9227_out0 = v$G$AD_17191_out0;
assign v$G$AB_9246_out0 = v$G$AD_17191_out0;
assign v$G4_11152_out0 = v$G5_4560_out0 || v$G$CD_955_out0;
assign v$G4_11157_out0 = v$G5_4565_out0 || v$G$CD_960_out0;
assign v$G4_11163_out0 = v$G5_4571_out0 || v$G$CD_966_out0;
assign v$G4_11166_out0 = v$G5_4574_out0 || v$G$CD_969_out0;
assign v$G4_11171_out0 = v$G5_4579_out0 || v$G$CD_974_out0;
assign v$G4_11184_out0 = v$G5_4592_out0 || v$G$CD_987_out0;
assign v$G4_11275_out0 = v$G5_4683_out0 || v$G$CD_1078_out0;
assign v$G4_11280_out0 = v$G5_4688_out0 || v$G$CD_1083_out0;
assign v$G4_11286_out0 = v$G5_4694_out0 || v$G$CD_1089_out0;
assign v$G4_11289_out0 = v$G5_4697_out0 || v$G$CD_1092_out0;
assign v$G4_11294_out0 = v$G5_4702_out0 || v$G$CD_1097_out0;
assign v$G4_11307_out0 = v$G5_4715_out0 || v$G$CD_1110_out0;
assign v$END43_13194_out0 = v$G$AD_17206_out0;
assign v$END46_15047_out0 = v$G$AD_17191_out0;
assign v$END30_15715_out0 = v$G$AD_17195_out0;
assign v$END41_16667_out0 = v$G$AD_17184_out0;
assign v$SEL8_17659_out0 = v$OP1_3387_out0[23:1];
assign v$_17750_out0 = { v$_10357_out0,v$_17966_out0 };
assign v$C14_281_out0 = v$COUTD_6799_out0;
assign v$P$AD_734_out0 = v$G1_5569_out0;
assign v$P$AD_738_out0 = v$G1_5573_out0;
assign v$P$AD_757_out0 = v$G1_5592_out0;
assign v$P$AD_765_out0 = v$G1_5600_out0;
assign v$P$AD_767_out0 = v$G1_5602_out0;
assign v$P$AD_857_out0 = v$G1_5692_out0;
assign v$P$AD_861_out0 = v$G1_5696_out0;
assign v$P$AD_880_out0 = v$G1_5715_out0;
assign v$P$AD_888_out0 = v$G1_5723_out0;
assign v$P$AD_890_out0 = v$G1_5725_out0;
assign v$C17_2522_out0 = v$COUTD_6778_out0;
assign v$G5_4610_out0 = v$G$AB_9227_out0 && v$P$CD_10545_out0;
assign v$G5_4629_out0 = v$G$AB_9246_out0 && v$P$CD_10564_out0;
assign v$C23_4845_out0 = v$COUTD_6801_out0;
assign v$C9_5939_out0 = v$COUTD_6788_out0;
assign v$CINA_8562_out0 = v$COUTD_6778_out0;
assign v$CINA_8569_out0 = v$COUTD_6778_out0;
assign v$CINA_8573_out0 = v$COUTD_6799_out0;
assign v$CINA_8576_out0 = v$COUTD_6799_out0;
assign v$CINA_8584_out0 = v$COUTD_6778_out0;
assign v$G8_11436_out0 = v$CINA_8505_out0 && v$P$AB_2042_out0;
assign v$G8_11441_out0 = v$CINA_8510_out0 && v$P$AB_2047_out0;
assign v$G8_11447_out0 = v$CINA_8516_out0 && v$P$AB_2053_out0;
assign v$G8_11450_out0 = v$CINA_8519_out0 && v$P$AB_2056_out0;
assign v$G8_11455_out0 = v$CINA_8524_out0 && v$P$AB_2061_out0;
assign v$G8_11468_out0 = v$CINA_8537_out0 && v$P$AB_2074_out0;
assign v$G8_11559_out0 = v$CINA_8628_out0 && v$P$AB_2165_out0;
assign v$G8_11564_out0 = v$CINA_8633_out0 && v$P$AB_2170_out0;
assign v$G8_11570_out0 = v$CINA_8639_out0 && v$P$AB_2176_out0;
assign v$G8_11573_out0 = v$CINA_8642_out0 && v$P$AB_2179_out0;
assign v$G8_11578_out0 = v$CINA_8647_out0 && v$P$AB_2184_out0;
assign v$G8_11591_out0 = v$CINA_8660_out0 && v$P$AB_2197_out0;
assign v$C13_11778_out0 = v$COUTD_6808_out0;
assign v$C10_12734_out0 = v$COUTD_6809_out0;
assign {v$A4A_13155_out1,v$A4A_13155_out0 } = v$A3_14608_out0 + v$B3_9472_out0 + v$C2_2687_out0;
assign {v$A4A_13158_out1,v$A4A_13158_out0 } = v$A3_14611_out0 + v$B3_9475_out0 + v$C2_2690_out0;
assign v$C12_13522_out0 = v$COUTD_6787_out0;
assign v$G$AD_17127_out0 = v$G4_11152_out0;
assign v$G$AD_17132_out0 = v$G4_11157_out0;
assign v$G$AD_17138_out0 = v$G4_11163_out0;
assign v$G$AD_17141_out0 = v$G4_11166_out0;
assign v$G$AD_17146_out0 = v$G4_11171_out0;
assign v$G$AD_17159_out0 = v$G4_11184_out0;
assign v$G$AD_17250_out0 = v$G4_11275_out0;
assign v$G$AD_17255_out0 = v$G4_11280_out0;
assign v$G$AD_17261_out0 = v$G4_11286_out0;
assign v$G$AD_17264_out0 = v$G4_11289_out0;
assign v$G$AD_17269_out0 = v$G4_11294_out0;
assign v$G$AD_17282_out0 = v$G4_11307_out0;
assign v$_18001_out0 = { v$SEL8_17659_out0,v$CIN_16820_out0 };
assign v$C2_18180_out0 = v$C2_2687_out0;
assign v$C2_18183_out0 = v$C2_2690_out0;
assign v$C14_327_out0 = v$C14_281_out0;
assign v$G$CD_958_out0 = v$G$AD_17146_out0;
assign v$G$CD_984_out0 = v$G$AD_17127_out0;
assign v$G$CD_992_out0 = v$G$AD_17141_out0;
assign v$G$CD_1081_out0 = v$G$AD_17269_out0;
assign v$G$CD_1107_out0 = v$G$AD_17250_out0;
assign v$G$CD_1115_out0 = v$G$AD_17264_out0;
assign v$END10_1152_out0 = v$G$AD_17138_out0;
assign v$END10_1155_out0 = v$G$AD_17261_out0;
assign v$C10_1942_out0 = v$C10_12734_out0;
assign v$P$AB_2045_out0 = v$P$AD_757_out0;
assign v$P$AB_2054_out0 = v$P$AD_757_out0;
assign v$P$AB_2055_out0 = v$P$AD_734_out0;
assign v$P$AB_2066_out0 = v$P$AD_757_out0;
assign v$P$AB_2068_out0 = v$P$AD_757_out0;
assign v$P$AB_2075_out0 = v$P$AD_757_out0;
assign v$P$AB_2076_out0 = v$P$AD_734_out0;
assign v$P$AB_2168_out0 = v$P$AD_880_out0;
assign v$P$AB_2177_out0 = v$P$AD_880_out0;
assign v$P$AB_2178_out0 = v$P$AD_857_out0;
assign v$P$AB_2189_out0 = v$P$AD_880_out0;
assign v$P$AB_2191_out0 = v$P$AD_880_out0;
assign v$P$AB_2198_out0 = v$P$AD_880_out0;
assign v$P$AB_2199_out0 = v$P$AD_857_out0;
assign {v$A12A_4447_out1,v$A12A_4447_out0 } = v$A11_9964_out0 + v$B11_9118_out0 + v$C10_12734_out0;
assign v$C17_6068_out0 = v$C17_2522_out0;
assign {v$A13_7242_out1,v$A13_7242_out0 } = v$A15_17320_out0 + v$B15_10023_out0 + v$C14_281_out0;
assign v$END15_7383_out0 = v$P$AD_738_out0;
assign v$END15_7386_out0 = v$P$AD_861_out0;
assign v$END17_7638_out0 = v$P$AD_767_out0;
assign v$END17_7641_out0 = v$P$AD_890_out0;
assign v$END3_7933_out0 = v$A4A_13155_out1;
assign v$END3_7936_out0 = v$A4A_13158_out1;
assign v$G$AB_9183_out0 = v$G$AD_17159_out0;
assign v$G$AB_9187_out0 = v$G$AD_17159_out0;
assign v$G$AB_9206_out0 = v$G$AD_17159_out0;
assign v$G$AB_9214_out0 = v$G$AD_17146_out0;
assign v$G$AB_9216_out0 = v$G$AD_17159_out0;
assign v$G$AB_9306_out0 = v$G$AD_17282_out0;
assign v$G$AB_9310_out0 = v$G$AD_17282_out0;
assign v$G$AB_9329_out0 = v$G$AD_17282_out0;
assign v$G$AB_9337_out0 = v$G$AD_17269_out0;
assign v$G$AB_9339_out0 = v$G$AD_17282_out0;
assign v$C12_9396_out0 = v$C12_13522_out0;
assign v$G7_9676_out0 = v$G8_11436_out0 && v$P$CD_10495_out0;
assign v$G7_9681_out0 = v$G8_11441_out0 && v$P$CD_10500_out0;
assign v$G7_9687_out0 = v$G8_11447_out0 && v$P$CD_10506_out0;
assign v$G7_9690_out0 = v$G8_11450_out0 && v$P$CD_10509_out0;
assign v$G7_9695_out0 = v$G8_11455_out0 && v$P$CD_10514_out0;
assign v$G7_9708_out0 = v$G8_11468_out0 && v$P$CD_10527_out0;
assign v$G7_9799_out0 = v$G8_11559_out0 && v$P$CD_10618_out0;
assign v$G7_9804_out0 = v$G8_11564_out0 && v$P$CD_10623_out0;
assign v$G7_9810_out0 = v$G8_11570_out0 && v$P$CD_10629_out0;
assign v$G7_9813_out0 = v$G8_11573_out0 && v$P$CD_10632_out0;
assign v$G7_9818_out0 = v$G8_11578_out0 && v$P$CD_10637_out0;
assign v$G7_9831_out0 = v$G8_11591_out0 && v$P$CD_10650_out0;
assign {v$A18_10034_out1,v$A18_10034_out0 } = v$A13_13864_out0 + v$B13_8677_out0 + v$C12_13522_out0;
assign v$P$CD_10521_out0 = v$P$AD_765_out0;
assign v$P$CD_10644_out0 = v$P$AD_888_out0;
assign v$END12_10781_out0 = v$G$AD_17132_out0;
assign v$END12_10784_out0 = v$G$AD_17255_out0;
assign v$G4_11202_out0 = v$G5_4610_out0 || v$G$CD_1005_out0;
assign v$G4_11221_out0 = v$G5_4629_out0 || v$G$CD_1024_out0;
assign v$G8_11493_out0 = v$CINA_8562_out0 && v$P$AB_2099_out0;
assign v$G8_11500_out0 = v$CINA_8569_out0 && v$P$AB_2106_out0;
assign v$G8_11504_out0 = v$CINA_8573_out0 && v$P$AB_2110_out0;
assign v$G8_11507_out0 = v$CINA_8576_out0 && v$P$AB_2113_out0;
assign v$G8_11515_out0 = v$CINA_8584_out0 && v$P$AB_2121_out0;
assign v$END19_11656_out0 = v$P$AD_734_out0;
assign v$END19_11659_out0 = v$P$AD_857_out0;
assign v$C9_12157_out0 = v$C9_5939_out0;
assign {v$A15_13218_out1,v$A15_13218_out0 } = v$A18_17697_out0 + v$B18_10869_out0 + v$C17_2522_out0;
assign {v$A16A_14561_out1,v$A16A_14561_out0 } = v$A10_1550_out0 + v$B10_9879_out0 + v$C9_5939_out0;
assign {v$A1_15222_out1,v$A1_15222_out0 } = v$_18001_out0 + v$MUX1_8346_out0 + v$C6_11358_out0;
assign v$C23_16151_out0 = v$C23_4845_out0;
assign {v$A20_16376_out1,v$A20_16376_out0 } = v$A14_678_out0 + v$B14_4004_out0 + v$C13_11778_out0;
assign v$C13_18591_out0 = v$C13_11778_out0;
assign v$_18665_out0 = { v$A3A_11952_out0,v$A4A_13155_out0 };
assign v$_18668_out0 = { v$A3A_11955_out0,v$A4A_13158_out0 };
assign v$G6_474_out0 = v$G4_11152_out0 || v$G7_9676_out0;
assign v$G6_479_out0 = v$G4_11157_out0 || v$G7_9681_out0;
assign v$G6_485_out0 = v$G4_11163_out0 || v$G7_9687_out0;
assign v$G6_488_out0 = v$G4_11166_out0 || v$G7_9690_out0;
assign v$G6_493_out0 = v$G4_11171_out0 || v$G7_9695_out0;
assign v$G6_506_out0 = v$G4_11184_out0 || v$G7_9708_out0;
assign v$G6_597_out0 = v$G4_11275_out0 || v$G7_9799_out0;
assign v$G6_602_out0 = v$G4_11280_out0 || v$G7_9804_out0;
assign v$G6_608_out0 = v$G4_11286_out0 || v$G7_9810_out0;
assign v$G6_611_out0 = v$G4_11289_out0 || v$G7_9813_out0;
assign v$G6_616_out0 = v$G4_11294_out0 || v$G7_9818_out0;
assign v$G6_629_out0 = v$G4_11307_out0 || v$G7_9831_out0;
assign v$ENDq_1460_out0 = v$A12A_4447_out1;
assign v$G5_4566_out0 = v$G$AB_9183_out0 && v$P$CD_10501_out0;
assign v$G5_4570_out0 = v$G$AB_9187_out0 && v$P$CD_10505_out0;
assign v$G5_4589_out0 = v$G$AB_9206_out0 && v$P$CD_10524_out0;
assign v$G5_4597_out0 = v$G$AB_9214_out0 && v$P$CD_10532_out0;
assign v$G5_4599_out0 = v$G$AB_9216_out0 && v$P$CD_10534_out0;
assign v$G5_4689_out0 = v$G$AB_9306_out0 && v$P$CD_10624_out0;
assign v$G5_4693_out0 = v$G$AB_9310_out0 && v$P$CD_10628_out0;
assign v$G5_4712_out0 = v$G$AB_9329_out0 && v$P$CD_10647_out0;
assign v$G5_4720_out0 = v$G$AB_9337_out0 && v$P$CD_10655_out0;
assign v$G5_4722_out0 = v$G$AB_9339_out0 && v$P$CD_10657_out0;
assign v$G1_5566_out0 = v$P$AB_2045_out0 && v$P$CD_10498_out0;
assign v$G1_5575_out0 = v$P$AB_2054_out0 && v$P$CD_10507_out0;
assign v$G1_5576_out0 = v$P$AB_2055_out0 && v$P$CD_10508_out0;
assign v$G1_5587_out0 = v$P$AB_2066_out0 && v$P$CD_10519_out0;
assign v$G1_5589_out0 = v$P$AB_2068_out0 && v$P$CD_10521_out0;
assign v$G1_5596_out0 = v$P$AB_2075_out0 && v$P$CD_10528_out0;
assign v$G1_5597_out0 = v$P$AB_2076_out0 && v$P$CD_10529_out0;
assign v$G1_5689_out0 = v$P$AB_2168_out0 && v$P$CD_10621_out0;
assign v$G1_5698_out0 = v$P$AB_2177_out0 && v$P$CD_10630_out0;
assign v$G1_5699_out0 = v$P$AB_2178_out0 && v$P$CD_10631_out0;
assign v$G1_5710_out0 = v$P$AB_2189_out0 && v$P$CD_10642_out0;
assign v$G1_5712_out0 = v$P$AB_2191_out0 && v$P$CD_10644_out0;
assign v$G1_5719_out0 = v$P$AB_2198_out0 && v$P$CD_10651_out0;
assign v$G1_5720_out0 = v$P$AB_2199_out0 && v$P$CD_10652_out0;
assign v$_5898_out0 = { v$A17A_2489_out0,v$A18_10034_out0 };
assign v$CARRY_6334_out0 = v$C23_16151_out0;
assign v$ENDr_7524_out0 = v$A20_16376_out1;
assign v$_7554_out0 = { v$C8_18499_out0,v$C9_12157_out0 };
assign v$COUT_8119_out0 = v$A1_15222_out1;
assign v$ENDi_8684_out0 = v$A15_13218_out1;
assign v$END0_9354_out0 = v$A16A_14561_out1;
assign v$G7_9733_out0 = v$G8_11493_out0 && v$P$CD_10552_out0;
assign v$G7_9740_out0 = v$G8_11500_out0 && v$P$CD_10559_out0;
assign v$G7_9744_out0 = v$G8_11504_out0 && v$P$CD_10563_out0;
assign v$G7_9747_out0 = v$G8_11507_out0 && v$P$CD_10566_out0;
assign v$G7_9755_out0 = v$G8_11515_out0 && v$P$CD_10574_out0;
assign v$_10239_out0 = { v$C12_9396_out0,v$C13_18591_out0 };
assign v$ENDt_10260_out0 = v$A13_7242_out1;
assign v$_10356_out0 = { v$_13438_out0,v$_18665_out0 };
assign v$_10359_out0 = { v$_13441_out0,v$_18668_out0 };
assign v$_10960_out0 = { v$A16A_14561_out0,v$A12A_4447_out0 };
assign v$_14838_out0 = { v$C10_1942_out0,v$C11_9512_out0 };
assign v$SUM_15174_out0 = v$A1_15222_out0;
assign v$G$AD_17177_out0 = v$G4_11202_out0;
assign v$G$AD_17196_out0 = v$G4_11221_out0;
assign v$_17458_out0 = { v$A20_16376_out0,v$A13_7242_out0 };
assign v$ENDe_17894_out0 = v$A18_10034_out1;
assign v$G6_531_out0 = v$G4_11209_out0 || v$G7_9733_out0;
assign v$G6_538_out0 = v$G4_11216_out0 || v$G7_9740_out0;
assign v$G6_542_out0 = v$G4_11220_out0 || v$G7_9744_out0;
assign v$G6_545_out0 = v$G4_11223_out0 || v$G7_9747_out0;
assign v$G6_553_out0 = v$G4_11231_out0 || v$G7_9755_out0;
assign v$P$AD_731_out0 = v$G1_5566_out0;
assign v$P$AD_740_out0 = v$G1_5575_out0;
assign v$P$AD_741_out0 = v$G1_5576_out0;
assign v$P$AD_752_out0 = v$G1_5587_out0;
assign v$P$AD_754_out0 = v$G1_5589_out0;
assign v$P$AD_761_out0 = v$G1_5596_out0;
assign v$P$AD_762_out0 = v$G1_5597_out0;
assign v$P$AD_854_out0 = v$G1_5689_out0;
assign v$P$AD_863_out0 = v$G1_5698_out0;
assign v$P$AD_864_out0 = v$G1_5699_out0;
assign v$P$AD_875_out0 = v$G1_5710_out0;
assign v$P$AD_877_out0 = v$G1_5712_out0;
assign v$P$AD_884_out0 = v$G1_5719_out0;
assign v$P$AD_885_out0 = v$G1_5720_out0;
assign v$_1559_out0 = { v$_15015_out0,v$_10960_out0 };
assign v$SUM_3474_out0 = v$SUM_15174_out0;
assign v$COUTD_6734_out0 = v$G6_474_out0;
assign v$COUTD_6739_out0 = v$G6_479_out0;
assign v$COUTD_6745_out0 = v$G6_485_out0;
assign v$COUTD_6748_out0 = v$G6_488_out0;
assign v$COUTD_6753_out0 = v$G6_493_out0;
assign v$COUTD_6766_out0 = v$G6_506_out0;
assign v$COUTD_6857_out0 = v$G6_597_out0;
assign v$COUTD_6862_out0 = v$G6_602_out0;
assign v$COUTD_6868_out0 = v$G6_608_out0;
assign v$COUTD_6871_out0 = v$G6_611_out0;
assign v$COUTD_6876_out0 = v$G6_616_out0;
assign v$COUTD_6889_out0 = v$G6_629_out0;
assign v$END50_7415_out0 = v$G$AD_17177_out0;
assign v$END48_10367_out0 = v$G$AD_17196_out0;
assign v$COUT_10736_out0 = v$COUT_8119_out0;
assign v$G4_11158_out0 = v$G5_4566_out0 || v$G$CD_961_out0;
assign v$G4_11162_out0 = v$G5_4570_out0 || v$G$CD_965_out0;
assign v$G4_11181_out0 = v$G5_4589_out0 || v$G$CD_984_out0;
assign v$G4_11189_out0 = v$G5_4597_out0 || v$G$CD_992_out0;
assign v$G4_11191_out0 = v$G5_4599_out0 || v$G$CD_994_out0;
assign v$G4_11281_out0 = v$G5_4689_out0 || v$G$CD_1084_out0;
assign v$G4_11285_out0 = v$G5_4693_out0 || v$G$CD_1088_out0;
assign v$G4_11304_out0 = v$G5_4712_out0 || v$G$CD_1107_out0;
assign v$G4_11312_out0 = v$G5_4720_out0 || v$G$CD_1115_out0;
assign v$G4_11314_out0 = v$G5_4722_out0 || v$G$CD_1117_out0;
assign v$_14295_out0 = { v$_5898_out0,v$_17458_out0 };
assign v$_18305_out0 = { v$_7554_out0,v$_14838_out0 };
assign v$_1175_out0 = { v$_1559_out0,v$_14295_out0 };
assign v$C4_1260_out0 = v$COUTD_6739_out0;
assign v$C4_1263_out0 = v$COUTD_6862_out0;
assign v$SEL10_1815_out0 = v$SUM_3474_out0[0:0];
assign v$P$AB_2058_out0 = v$P$AD_731_out0;
assign v$P$AB_2065_out0 = v$P$AD_731_out0;
assign v$P$AB_2069_out0 = v$P$AD_752_out0;
assign v$P$AB_2072_out0 = v$P$AD_752_out0;
assign v$P$AB_2080_out0 = v$P$AD_731_out0;
assign v$P$AB_2181_out0 = v$P$AD_854_out0;
assign v$P$AB_2188_out0 = v$P$AD_854_out0;
assign v$P$AB_2192_out0 = v$P$AD_875_out0;
assign v$P$AB_2195_out0 = v$P$AD_875_out0;
assign v$P$AB_2203_out0 = v$P$AD_854_out0;
assign v$END27_2211_out0 = v$P$AD_761_out0;
assign v$END27_2214_out0 = v$P$AD_884_out0;
assign v$CIN_3892_out0 = v$COUT_10736_out0;
assign v$END21_4341_out0 = v$P$AD_741_out0;
assign v$END21_4344_out0 = v$P$AD_864_out0;
assign v$END40_5776_out0 = v$COUTD_6753_out0;
assign v$END40_5779_out0 = v$COUTD_6876_out0;
assign v$END29_5886_out0 = v$P$AD_752_out0;
assign v$END29_5889_out0 = v$P$AD_875_out0;
assign v$COUTD_6791_out0 = v$G6_531_out0;
assign v$COUTD_6798_out0 = v$G6_538_out0;
assign v$COUTD_6802_out0 = v$G6_542_out0;
assign v$COUTD_6805_out0 = v$G6_545_out0;
assign v$COUTD_6813_out0 = v$G6_553_out0;
assign v$CINA_8511_out0 = v$COUTD_6766_out0;
assign v$CINA_8515_out0 = v$COUTD_6766_out0;
assign v$CINA_8534_out0 = v$COUTD_6766_out0;
assign v$CINA_8542_out0 = v$COUTD_6753_out0;
assign v$CINA_8544_out0 = v$COUTD_6766_out0;
assign v$CINA_8634_out0 = v$COUTD_6889_out0;
assign v$CINA_8638_out0 = v$COUTD_6889_out0;
assign v$CINA_8657_out0 = v$COUTD_6889_out0;
assign v$CINA_8665_out0 = v$COUTD_6876_out0;
assign v$CINA_8667_out0 = v$COUTD_6889_out0;
assign v$END4_9368_out0 = v$COUTD_6734_out0;
assign v$END4_9371_out0 = v$COUTD_6857_out0;
assign v$END52_11974_out0 = v$P$AD_754_out0;
assign v$END52_11977_out0 = v$P$AD_877_out0;
assign v$OP1_14191_out0 = v$SUM_3474_out0;
assign v$END60_15133_out0 = v$COUTD_6748_out0;
assign v$END60_15136_out0 = v$COUTD_6871_out0;
assign v$C3_15727_out0 = v$COUTD_6745_out0;
assign v$C3_15730_out0 = v$COUTD_6868_out0;
assign v$C5_15916_out0 = v$COUTD_6766_out0;
assign v$C5_15919_out0 = v$COUTD_6889_out0;
assign v$END23_16718_out0 = v$P$AD_762_out0;
assign v$END23_16721_out0 = v$P$AD_885_out0;
assign v$END25_17071_out0 = v$P$AD_740_out0;
assign v$END25_17074_out0 = v$P$AD_863_out0;
assign v$G$AD_17133_out0 = v$G4_11158_out0;
assign v$G$AD_17137_out0 = v$G4_11162_out0;
assign v$G$AD_17156_out0 = v$G4_11181_out0;
assign v$G$AD_17164_out0 = v$G4_11189_out0;
assign v$G$AD_17166_out0 = v$G4_11191_out0;
assign v$G$AD_17256_out0 = v$G4_11281_out0;
assign v$G$AD_17260_out0 = v$G4_11285_out0;
assign v$G$AD_17279_out0 = v$G4_11304_out0;
assign v$G$AD_17287_out0 = v$G4_11312_out0;
assign v$G$AD_17289_out0 = v$G4_11314_out0;
assign v$END16_217_out0 = v$G$AD_17166_out0;
assign v$END16_220_out0 = v$G$AD_17289_out0;
assign v$END14_275_out0 = v$G$AD_17137_out0;
assign v$END14_278_out0 = v$G$AD_17260_out0;
assign v$G$CD_981_out0 = v$G$AD_17164_out0;
assign v$G$CD_1104_out0 = v$G$AD_17287_out0;
assign v$C16_1270_out0 = v$COUTD_6805_out0;
assign {v$A7A_1658_out1,v$A7A_1658_out0 } = v$A5_6666_out0 + v$B5_18375_out0 + v$C4_1260_out0;
assign {v$A7A_1661_out1,v$A7A_1661_out0 } = v$A5_6669_out0 + v$B5_18378_out0 + v$C4_1263_out0;
assign v$C4_1877_out0 = v$C4_1260_out0;
assign v$C4_1880_out0 = v$C4_1263_out0;
assign {v$A6A_3122_out1,v$A6A_3122_out0 } = v$A6_309_out0 + v$B6_13299_out0 + v$C5_15916_out0;
assign {v$A6A_3125_out1,v$A6A_3125_out0 } = v$A6_312_out0 + v$B6_13302_out0 + v$C5_15919_out0;
assign v$OP1_3385_out0 = v$OP1_14191_out0;
assign v$G1_5579_out0 = v$P$AB_2058_out0 && v$P$CD_10511_out0;
assign v$G1_5586_out0 = v$P$AB_2065_out0 && v$P$CD_10518_out0;
assign v$G1_5590_out0 = v$P$AB_2069_out0 && v$P$CD_10522_out0;
assign v$G1_5593_out0 = v$P$AB_2072_out0 && v$P$CD_10525_out0;
assign v$G1_5601_out0 = v$P$AB_2080_out0 && v$P$CD_10533_out0;
assign v$G1_5702_out0 = v$P$AB_2181_out0 && v$P$CD_10634_out0;
assign v$G1_5709_out0 = v$P$AB_2188_out0 && v$P$CD_10641_out0;
assign v$G1_5713_out0 = v$P$AB_2192_out0 && v$P$CD_10645_out0;
assign v$G1_5716_out0 = v$P$AB_2195_out0 && v$P$CD_10648_out0;
assign v$G1_5724_out0 = v$P$AB_2203_out0 && v$P$CD_10656_out0;
assign v$C15_8145_out0 = v$COUTD_6802_out0;
assign v$C19_8162_out0 = v$COUTD_6813_out0;
assign v$CINA_8555_out0 = v$COUTD_6798_out0;
assign v$CINA_8574_out0 = v$COUTD_6798_out0;
assign v$G$AB_9180_out0 = v$G$AD_17156_out0;
assign v$G$AB_9189_out0 = v$G$AD_17156_out0;
assign v$G$AB_9190_out0 = v$G$AD_17133_out0;
assign v$G$AB_9201_out0 = v$G$AD_17156_out0;
assign v$G$AB_9203_out0 = v$G$AD_17156_out0;
assign v$G$AB_9210_out0 = v$G$AD_17156_out0;
assign v$G$AB_9211_out0 = v$G$AD_17133_out0;
assign v$G$AB_9303_out0 = v$G$AD_17279_out0;
assign v$G$AB_9312_out0 = v$G$AD_17279_out0;
assign v$G$AB_9313_out0 = v$G$AD_17256_out0;
assign v$G$AB_9324_out0 = v$G$AD_17279_out0;
assign v$G$AB_9326_out0 = v$G$AD_17279_out0;
assign v$G$AB_9333_out0 = v$G$AD_17279_out0;
assign v$G$AB_9334_out0 = v$G$AD_17256_out0;
assign v$G8_11442_out0 = v$CINA_8511_out0 && v$P$AB_2048_out0;
assign v$G8_11446_out0 = v$CINA_8515_out0 && v$P$AB_2052_out0;
assign v$G8_11465_out0 = v$CINA_8534_out0 && v$P$AB_2071_out0;
assign v$G8_11473_out0 = v$CINA_8542_out0 && v$P$AB_2079_out0;
assign v$G8_11475_out0 = v$CINA_8544_out0 && v$P$AB_2081_out0;
assign v$G8_11565_out0 = v$CINA_8634_out0 && v$P$AB_2171_out0;
assign v$G8_11569_out0 = v$CINA_8638_out0 && v$P$AB_2175_out0;
assign v$G8_11588_out0 = v$CINA_8657_out0 && v$P$AB_2194_out0;
assign v$G8_11596_out0 = v$CINA_8665_out0 && v$P$AB_2202_out0;
assign v$G8_11598_out0 = v$CINA_8667_out0 && v$P$AB_2204_out0;
assign v$C5_11687_out0 = v$C5_15916_out0;
assign v$C5_11690_out0 = v$C5_15919_out0;
assign v$END18_11947_out0 = v$G$AD_17133_out0;
assign v$END18_11950_out0 = v$G$AD_17256_out0;
assign v$SUM$6_12912_out0 = v$SEL10_1815_out0;
assign v$C20_15491_out0 = v$COUTD_6798_out0;
assign v$C3_15818_out0 = v$C3_15727_out0;
assign v$C3_15821_out0 = v$C3_15730_out0;
assign {v$A5A_16100_out1,v$A5A_16100_out0 } = v$A4_17499_out0 + v$B4_14664_out0 + v$C3_15727_out0;
assign {v$A5A_16103_out1,v$A5A_16103_out0 } = v$A4_17502_out0 + v$B4_14667_out0 + v$C3_15730_out0;
assign v$C18_16291_out0 = v$COUTD_6791_out0;
assign v$CIN_16818_out0 = v$CIN_3892_out0;
assign v$_18235_out0 = { v$_17750_out0,v$_1175_out0 };
assign v$_83_out0 = { v$A5A_16100_out0,v$A7A_1658_out0 };
assign v$_86_out0 = { v$A5A_16103_out0,v$A7A_1661_out0 };
assign v$P$AD_744_out0 = v$G1_5579_out0;
assign v$P$AD_751_out0 = v$G1_5586_out0;
assign v$P$AD_755_out0 = v$G1_5590_out0;
assign v$P$AD_758_out0 = v$G1_5593_out0;
assign v$P$AD_766_out0 = v$G1_5601_out0;
assign v$P$AD_867_out0 = v$G1_5702_out0;
assign v$P$AD_874_out0 = v$G1_5709_out0;
assign v$P$AD_878_out0 = v$G1_5713_out0;
assign v$P$AD_881_out0 = v$G1_5716_out0;
assign v$P$AD_889_out0 = v$G1_5724_out0;
assign v$_2454_out0 = { v$C4_1877_out0,v$C5_11687_out0 };
assign v$_2457_out0 = { v$C4_1880_out0,v$C5_11690_out0 };
assign v$END5_4144_out0 = v$A7A_1658_out1;
assign v$END5_4147_out0 = v$A7A_1661_out1;
assign v$G5_4563_out0 = v$G$AB_9180_out0 && v$P$CD_10498_out0;
assign v$G5_4572_out0 = v$G$AB_9189_out0 && v$P$CD_10507_out0;
assign v$G5_4573_out0 = v$G$AB_9190_out0 && v$P$CD_10508_out0;
assign v$G5_4584_out0 = v$G$AB_9201_out0 && v$P$CD_10519_out0;
assign v$G5_4586_out0 = v$G$AB_9203_out0 && v$P$CD_10521_out0;
assign v$G5_4593_out0 = v$G$AB_9210_out0 && v$P$CD_10528_out0;
assign v$G5_4594_out0 = v$G$AB_9211_out0 && v$P$CD_10529_out0;
assign v$G5_4686_out0 = v$G$AB_9303_out0 && v$P$CD_10621_out0;
assign v$G5_4695_out0 = v$G$AB_9312_out0 && v$P$CD_10630_out0;
assign v$G5_4696_out0 = v$G$AB_9313_out0 && v$P$CD_10631_out0;
assign v$G5_4707_out0 = v$G$AB_9324_out0 && v$P$CD_10642_out0;
assign v$G5_4709_out0 = v$G$AB_9326_out0 && v$P$CD_10644_out0;
assign v$G5_4716_out0 = v$G$AB_9333_out0 && v$P$CD_10651_out0;
assign v$G5_4717_out0 = v$G$AB_9334_out0 && v$P$CD_10652_out0;
assign v$END4_5247_out0 = v$A5A_16100_out1;
assign v$END4_5250_out0 = v$A5A_16103_out1;
assign v$G7_9682_out0 = v$G8_11442_out0 && v$P$CD_10501_out0;
assign v$G7_9686_out0 = v$G8_11446_out0 && v$P$CD_10505_out0;
assign v$G7_9705_out0 = v$G8_11465_out0 && v$P$CD_10524_out0;
assign v$G7_9713_out0 = v$G8_11473_out0 && v$P$CD_10532_out0;
assign v$G7_9715_out0 = v$G8_11475_out0 && v$P$CD_10534_out0;
assign v$G7_9805_out0 = v$G8_11565_out0 && v$P$CD_10624_out0;
assign v$G7_9809_out0 = v$G8_11569_out0 && v$P$CD_10628_out0;
assign v$G7_9828_out0 = v$G8_11588_out0 && v$P$CD_10647_out0;
assign v$G7_9836_out0 = v$G8_11596_out0 && v$P$CD_10655_out0;
assign v$G7_9838_out0 = v$G8_11598_out0 && v$P$CD_10657_out0;
assign v$G8_11486_out0 = v$CINA_8555_out0 && v$P$AB_2092_out0;
assign v$G8_11505_out0 = v$CINA_8574_out0 && v$P$AB_2111_out0;
assign v$C15_13133_out0 = v$C15_8145_out0;
assign v$C19_13835_out0 = v$C19_8162_out0;
assign v$C20_14980_out0 = v$C20_15491_out0;
assign v$_14999_out0 = { v$C2_18180_out0,v$C3_15818_out0 };
assign v$_15002_out0 = { v$C2_18183_out0,v$C3_15821_out0 };
assign v$C16_15159_out0 = v$C16_1270_out0;
assign v$END6_15250_out0 = v$A6A_3122_out1;
assign v$END6_15253_out0 = v$A6A_3125_out1;
assign {v$A14_15355_out1,v$A14_15355_out0 } = v$A16_13616_out0 + v$B16_16416_out0 + v$C15_8145_out0;
assign {v$A19_15910_out1,v$A19_15910_out0 } = v$A19_1215_out0 + v$B19_16791_out0 + v$C18_16291_out0;
assign {v$A24_16975_out1,v$A24_16975_out0 } = v$A21_2600_out0 + v$B21_18084_out0 + v$C20_15491_out0;
assign {v$A22_17490_out1,v$A22_17490_out0 } = v$A20_4438_out0 + v$B20_3945_out0 + v$C19_8162_out0;
assign v$SEL8_17657_out0 = v$OP1_3385_out0[23:1];
assign {v$A11_17876_out1,v$A11_17876_out0 } = v$A17_16724_out0 + v$B17_15537_out0 + v$C16_1270_out0;
assign v$C18_18007_out0 = v$C18_16291_out0;
assign v$END33_265_out0 = v$P$AD_758_out0;
assign v$END33_268_out0 = v$P$AD_881_out0;
assign v$G6_480_out0 = v$G4_11158_out0 || v$G7_9682_out0;
assign v$G6_484_out0 = v$G4_11162_out0 || v$G7_9686_out0;
assign v$G6_503_out0 = v$G4_11181_out0 || v$G7_9705_out0;
assign v$G6_511_out0 = v$G4_11189_out0 || v$G7_9713_out0;
assign v$G6_513_out0 = v$G4_11191_out0 || v$G7_9715_out0;
assign v$G6_603_out0 = v$G4_11281_out0 || v$G7_9805_out0;
assign v$G6_607_out0 = v$G4_11285_out0 || v$G7_9809_out0;
assign v$G6_626_out0 = v$G4_11304_out0 || v$G7_9828_out0;
assign v$G6_634_out0 = v$G4_11312_out0 || v$G7_9836_out0;
assign v$G6_636_out0 = v$G4_11314_out0 || v$G7_9838_out0;
assign v$_1201_out0 = { v$A15_13218_out0,v$A19_15910_out0 };
assign v$_1795_out0 = { v$A22_17490_out0,v$A24_16975_out0 };
assign v$P$AB_2051_out0 = v$P$AD_751_out0;
assign v$P$AB_2070_out0 = v$P$AD_751_out0;
assign v$P$AB_2174_out0 = v$P$AD_874_out0;
assign v$P$AB_2193_out0 = v$P$AD_874_out0;
assign v$END47_2680_out0 = v$P$AD_751_out0;
assign v$END47_2683_out0 = v$P$AD_874_out0;
assign v$_2842_out0 = { v$C14_327_out0,v$C15_13133_out0 };
assign v$ENDp_3191_out0 = v$A22_17490_out1;
assign v$ENDy_4116_out0 = v$A14_15355_out1;
assign v$ENDu_7031_out0 = v$A11_17876_out1;
assign v$_7254_out0 = { v$_8907_out0,v$_14999_out0 };
assign v$_7257_out0 = { v$_8910_out0,v$_15002_out0 };
assign v$_7870_out0 = { v$C16_15159_out0,v$C17_6068_out0 };
assign v$_8331_out0 = { v$C18_18007_out0,v$C19_13835_out0 };
assign v$G7_9726_out0 = v$G8_11486_out0 && v$P$CD_10545_out0;
assign v$G7_9745_out0 = v$G8_11505_out0 && v$P$CD_10564_out0;
assign v$G4_11155_out0 = v$G5_4563_out0 || v$G$CD_958_out0;
assign v$G4_11164_out0 = v$G5_4572_out0 || v$G$CD_967_out0;
assign v$G4_11165_out0 = v$G5_4573_out0 || v$G$CD_968_out0;
assign v$G4_11176_out0 = v$G5_4584_out0 || v$G$CD_979_out0;
assign v$G4_11178_out0 = v$G5_4586_out0 || v$G$CD_981_out0;
assign v$G4_11185_out0 = v$G5_4593_out0 || v$G$CD_988_out0;
assign v$G4_11186_out0 = v$G5_4594_out0 || v$G$CD_989_out0;
assign v$G4_11278_out0 = v$G5_4686_out0 || v$G$CD_1081_out0;
assign v$G4_11287_out0 = v$G5_4695_out0 || v$G$CD_1090_out0;
assign v$G4_11288_out0 = v$G5_4696_out0 || v$G$CD_1091_out0;
assign v$G4_11299_out0 = v$G5_4707_out0 || v$G$CD_1102_out0;
assign v$G4_11301_out0 = v$G5_4709_out0 || v$G$CD_1104_out0;
assign v$G4_11308_out0 = v$G5_4716_out0 || v$G$CD_1111_out0;
assign v$G4_11309_out0 = v$G5_4717_out0 || v$G$CD_1112_out0;
assign v$_13295_out0 = { v$A14_15355_out0,v$A11_17876_out0 };
assign v$END44_15666_out0 = v$P$AD_766_out0;
assign v$END44_15669_out0 = v$P$AD_889_out0;
assign v$ENDa_16566_out0 = v$A24_16975_out1;
assign v$_17999_out0 = { v$SEL8_17657_out0,v$CIN_16818_out0 };
assign v$END42_18312_out0 = v$P$AD_744_out0;
assign v$END42_18315_out0 = v$P$AD_867_out0;
assign v$END31_18521_out0 = v$P$AD_755_out0;
assign v$END31_18524_out0 = v$P$AD_878_out0;
assign v$ENDo_18694_out0 = v$A19_15910_out1;
assign v$G6_524_out0 = v$G4_11202_out0 || v$G7_9726_out0;
assign v$G6_543_out0 = v$G4_11221_out0 || v$G7_9745_out0;
assign v$_1244_out0 = { v$_10239_out0,v$_2842_out0 };
assign v$G1_5572_out0 = v$P$AB_2051_out0 && v$P$CD_10504_out0;
assign v$G1_5591_out0 = v$P$AB_2070_out0 && v$P$CD_10523_out0;
assign v$G1_5695_out0 = v$P$AB_2174_out0 && v$P$CD_10627_out0;
assign v$G1_5714_out0 = v$P$AB_2193_out0 && v$P$CD_10646_out0;
assign v$COUTD_6740_out0 = v$G6_480_out0;
assign v$COUTD_6744_out0 = v$G6_484_out0;
assign v$COUTD_6763_out0 = v$G6_503_out0;
assign v$COUTD_6771_out0 = v$G6_511_out0;
assign v$COUTD_6773_out0 = v$G6_513_out0;
assign v$COUTD_6863_out0 = v$G6_603_out0;
assign v$COUTD_6867_out0 = v$G6_607_out0;
assign v$COUTD_6886_out0 = v$G6_626_out0;
assign v$COUTD_6894_out0 = v$G6_634_out0;
assign v$COUTD_6896_out0 = v$G6_636_out0;
assign v$_10351_out0 = { v$_7870_out0,v$_8331_out0 };
assign {v$A1_15220_out1,v$A1_15220_out0 } = v$_17999_out0 + v$MUX1_8344_out0 + v$C6_11356_out0;
assign v$_16258_out0 = { v$_13295_out0,v$_1201_out0 };
assign v$G$AD_17130_out0 = v$G4_11155_out0;
assign v$G$AD_17139_out0 = v$G4_11164_out0;
assign v$G$AD_17140_out0 = v$G4_11165_out0;
assign v$G$AD_17151_out0 = v$G4_11176_out0;
assign v$G$AD_17153_out0 = v$G4_11178_out0;
assign v$G$AD_17160_out0 = v$G4_11185_out0;
assign v$G$AD_17161_out0 = v$G4_11186_out0;
assign v$G$AD_17253_out0 = v$G4_11278_out0;
assign v$G$AD_17262_out0 = v$G4_11287_out0;
assign v$G$AD_17263_out0 = v$G4_11288_out0;
assign v$G$AD_17274_out0 = v$G4_11299_out0;
assign v$G$AD_17276_out0 = v$G4_11301_out0;
assign v$G$AD_17283_out0 = v$G4_11308_out0;
assign v$G$AD_17284_out0 = v$G4_11309_out0;
assign v$END53_318_out0 = v$G$AD_17153_out0;
assign v$END53_321_out0 = v$G$AD_17276_out0;
assign v$P$AD_737_out0 = v$G1_5572_out0;
assign v$P$AD_756_out0 = v$G1_5591_out0;
assign v$P$AD_860_out0 = v$G1_5695_out0;
assign v$P$AD_879_out0 = v$G1_5714_out0;
assign v$END26_6436_out0 = v$G$AD_17160_out0;
assign v$END26_6439_out0 = v$G$AD_17283_out0;
assign v$COUTD_6784_out0 = v$G6_524_out0;
assign v$COUTD_6803_out0 = v$G6_543_out0;
assign v$C8_7431_out0 = v$COUTD_6740_out0;
assign v$C8_7434_out0 = v$COUTD_6863_out0;
assign v$COUT_8117_out0 = v$A1_15220_out1;
assign v$CINA_8508_out0 = v$COUTD_6763_out0;
assign v$CINA_8517_out0 = v$COUTD_6763_out0;
assign v$CINA_8518_out0 = v$COUTD_6740_out0;
assign v$CINA_8529_out0 = v$COUTD_6763_out0;
assign v$CINA_8531_out0 = v$COUTD_6763_out0;
assign v$CINA_8538_out0 = v$COUTD_6763_out0;
assign v$CINA_8539_out0 = v$COUTD_6740_out0;
assign v$CINA_8631_out0 = v$COUTD_6886_out0;
assign v$CINA_8640_out0 = v$COUTD_6886_out0;
assign v$CINA_8641_out0 = v$COUTD_6863_out0;
assign v$CINA_8652_out0 = v$COUTD_6886_out0;
assign v$CINA_8654_out0 = v$COUTD_6886_out0;
assign v$CINA_8661_out0 = v$COUTD_6886_out0;
assign v$CINA_8662_out0 = v$COUTD_6863_out0;
assign v$G$AB_9193_out0 = v$G$AD_17130_out0;
assign v$G$AB_9200_out0 = v$G$AD_17130_out0;
assign v$G$AB_9204_out0 = v$G$AD_17151_out0;
assign v$G$AB_9207_out0 = v$G$AD_17151_out0;
assign v$G$AB_9215_out0 = v$G$AD_17130_out0;
assign v$G$AB_9316_out0 = v$G$AD_17253_out0;
assign v$G$AB_9323_out0 = v$G$AD_17253_out0;
assign v$G$AB_9327_out0 = v$G$AD_17274_out0;
assign v$G$AB_9330_out0 = v$G$AD_17274_out0;
assign v$G$AB_9338_out0 = v$G$AD_17253_out0;
assign v$C6_9587_out0 = v$COUTD_6744_out0;
assign v$C6_9590_out0 = v$COUTD_6867_out0;
assign v$C7_10970_out0 = v$COUTD_6773_out0;
assign v$C7_10973_out0 = v$COUTD_6896_out0;
assign v$END20_13265_out0 = v$G$AD_17140_out0;
assign v$END20_13268_out0 = v$G$AD_17263_out0;
assign v$END28_13670_out0 = v$G$AD_17151_out0;
assign v$END28_13673_out0 = v$G$AD_17274_out0;
assign v$C11_14797_out0 = v$COUTD_6763_out0;
assign v$C11_14800_out0 = v$COUTD_6886_out0;
assign v$SUM_15172_out0 = v$A1_15220_out0;
assign v$END22_15485_out0 = v$G$AD_17161_out0;
assign v$END22_15488_out0 = v$G$AD_17284_out0;
assign v$END24_16404_out0 = v$G$AD_17139_out0;
assign v$END24_16407_out0 = v$G$AD_17262_out0;
assign v$_17355_out0 = { v$_18305_out0,v$_1244_out0 };
assign v$END61_17957_out0 = v$COUTD_6771_out0;
assign v$END61_17960_out0 = v$COUTD_6894_out0;
assign {v$A8A_1506_out1,v$A8A_1506_out0 } = v$A7_15308_out0 + v$B7_17041_out0 + v$C6_9587_out0;
assign {v$A8A_1509_out1,v$A8A_1509_out0 } = v$A7_15311_out0 + v$B7_17044_out0 + v$C6_9590_out0;
assign {v$A17A_2488_out1,v$A17A_2488_out0 } = v$A12_3139_out0 + v$B12_1951_out0 + v$C11_14797_out0;
assign {v$A17A_2491_out1,v$A17A_2491_out0 } = v$A12_3142_out0 + v$B12_1954_out0 + v$C11_14800_out0;
assign v$SUM_3472_out0 = v$SUM_15172_out0;
assign v$G5_4576_out0 = v$G$AB_9193_out0 && v$P$CD_10511_out0;
assign v$G5_4583_out0 = v$G$AB_9200_out0 && v$P$CD_10518_out0;
assign v$G5_4587_out0 = v$G$AB_9204_out0 && v$P$CD_10522_out0;
assign v$G5_4590_out0 = v$G$AB_9207_out0 && v$P$CD_10525_out0;
assign v$G5_4598_out0 = v$G$AB_9215_out0 && v$P$CD_10533_out0;
assign v$G5_4699_out0 = v$G$AB_9316_out0 && v$P$CD_10634_out0;
assign v$G5_4706_out0 = v$G$AB_9323_out0 && v$P$CD_10641_out0;
assign v$G5_4710_out0 = v$G$AB_9327_out0 && v$P$CD_10645_out0;
assign v$G5_4713_out0 = v$G$AB_9330_out0 && v$P$CD_10648_out0;
assign v$G5_4721_out0 = v$G$AB_9338_out0 && v$P$CD_10656_out0;
assign v$_4869_out0 = { v$_7792_out0,v$_17355_out0 };
assign v$C6_7056_out0 = v$C6_9587_out0;
assign v$C6_7059_out0 = v$C6_9590_out0;
assign v$C11_9511_out0 = v$C11_14797_out0;
assign v$C11_9514_out0 = v$C11_14800_out0;
assign {v$A9A_10412_out1,v$A9A_10412_out0 } = v$A8_18091_out0 + v$B8_13139_out0 + v$C7_10970_out0;
assign {v$A9A_10415_out1,v$A9A_10415_out0 } = v$A8_18094_out0 + v$B8_13142_out0 + v$C7_10973_out0;
assign v$COUT_10734_out0 = v$COUT_8117_out0;
assign v$C21_10769_out0 = v$COUTD_6803_out0;
assign v$C22_10983_out0 = v$COUTD_6784_out0;
assign v$G8_11439_out0 = v$CINA_8508_out0 && v$P$AB_2045_out0;
assign v$G8_11448_out0 = v$CINA_8517_out0 && v$P$AB_2054_out0;
assign v$G8_11449_out0 = v$CINA_8518_out0 && v$P$AB_2055_out0;
assign v$G8_11460_out0 = v$CINA_8529_out0 && v$P$AB_2066_out0;
assign v$G8_11462_out0 = v$CINA_8531_out0 && v$P$AB_2068_out0;
assign v$G8_11469_out0 = v$CINA_8538_out0 && v$P$AB_2075_out0;
assign v$G8_11470_out0 = v$CINA_8539_out0 && v$P$AB_2076_out0;
assign v$G8_11562_out0 = v$CINA_8631_out0 && v$P$AB_2168_out0;
assign v$G8_11571_out0 = v$CINA_8640_out0 && v$P$AB_2177_out0;
assign v$G8_11572_out0 = v$CINA_8641_out0 && v$P$AB_2178_out0;
assign v$G8_11583_out0 = v$CINA_8652_out0 && v$P$AB_2189_out0;
assign v$G8_11585_out0 = v$CINA_8654_out0 && v$P$AB_2191_out0;
assign v$G8_11592_out0 = v$CINA_8661_out0 && v$P$AB_2198_out0;
assign v$G8_11593_out0 = v$CINA_8662_out0 && v$P$AB_2199_out0;
assign v$END51_11677_out0 = v$P$AD_737_out0;
assign v$END51_11680_out0 = v$P$AD_860_out0;
assign {v$A10A_16003_out1,v$A10A_16003_out0 } = v$A9_3436_out0 + v$B9_4066_out0 + v$C8_7431_out0;
assign {v$A10A_16006_out1,v$A10A_16006_out0 } = v$A9_3439_out0 + v$B9_4069_out0 + v$C8_7434_out0;
assign v$C7_16431_out0 = v$C7_10970_out0;
assign v$C7_16434_out0 = v$C7_10973_out0;
assign v$END49_18451_out0 = v$P$AD_756_out0;
assign v$END49_18454_out0 = v$P$AD_879_out0;
assign v$C8_18498_out0 = v$C8_7431_out0;
assign v$C8_18501_out0 = v$C8_7434_out0;
assign v$SEL11_1500_out0 = v$SUM_3472_out0[0:0];
assign v$END7_3360_out0 = v$A8A_1506_out1;
assign v$END7_3363_out0 = v$A8A_1509_out1;
assign v$_3637_out0 = { v$A6A_3122_out0,v$A8A_1506_out0 };
assign v$_3640_out0 = { v$A6A_3125_out0,v$A8A_1509_out0 };
assign v$CIN_3888_out0 = v$COUT_10734_out0;
assign v$END8_3902_out0 = v$A9A_10412_out1;
assign v$END8_3905_out0 = v$A9A_10415_out1;
assign v$END9_4234_out0 = v$A10A_16003_out1;
assign v$END9_4237_out0 = v$A10A_16006_out1;
assign v$C21_6371_out0 = v$C21_10769_out0;
assign v$C22_8412_out0 = v$C22_10983_out0;
assign {v$A23_9548_out1,v$A23_9548_out0 } = v$A23_5065_out0 + v$B23_1285_out0 + v$C22_10983_out0;
assign v$ENDw_9552_out0 = v$A17A_2488_out1;
assign v$ENDw_9555_out0 = v$A17A_2491_out1;
assign v$G7_9679_out0 = v$G8_11439_out0 && v$P$CD_10498_out0;
assign v$G7_9688_out0 = v$G8_11448_out0 && v$P$CD_10507_out0;
assign v$G7_9689_out0 = v$G8_11449_out0 && v$P$CD_10508_out0;
assign v$G7_9700_out0 = v$G8_11460_out0 && v$P$CD_10519_out0;
assign v$G7_9702_out0 = v$G8_11462_out0 && v$P$CD_10521_out0;
assign v$G7_9709_out0 = v$G8_11469_out0 && v$P$CD_10528_out0;
assign v$G7_9710_out0 = v$G8_11470_out0 && v$P$CD_10529_out0;
assign v$G7_9802_out0 = v$G8_11562_out0 && v$P$CD_10621_out0;
assign v$G7_9811_out0 = v$G8_11571_out0 && v$P$CD_10630_out0;
assign v$G7_9812_out0 = v$G8_11572_out0 && v$P$CD_10631_out0;
assign v$G7_9823_out0 = v$G8_11583_out0 && v$P$CD_10642_out0;
assign v$G7_9825_out0 = v$G8_11585_out0 && v$P$CD_10644_out0;
assign v$G7_9832_out0 = v$G8_11592_out0 && v$P$CD_10651_out0;
assign v$G7_9833_out0 = v$G8_11593_out0 && v$P$CD_10652_out0;
assign v$G4_11168_out0 = v$G5_4576_out0 || v$G$CD_971_out0;
assign v$G4_11175_out0 = v$G5_4583_out0 || v$G$CD_978_out0;
assign v$G4_11179_out0 = v$G5_4587_out0 || v$G$CD_982_out0;
assign v$G4_11182_out0 = v$G5_4590_out0 || v$G$CD_985_out0;
assign v$G4_11190_out0 = v$G5_4598_out0 || v$G$CD_993_out0;
assign v$G4_11291_out0 = v$G5_4699_out0 || v$G$CD_1094_out0;
assign v$G4_11298_out0 = v$G5_4706_out0 || v$G$CD_1101_out0;
assign v$G4_11302_out0 = v$G5_4710_out0 || v$G$CD_1105_out0;
assign v$G4_11305_out0 = v$G5_4713_out0 || v$G$CD_1108_out0;
assign v$G4_11313_out0 = v$G5_4721_out0 || v$G$CD_1116_out0;
assign v$OP1_14187_out0 = v$SUM_3472_out0;
assign v$_15014_out0 = { v$A9A_10412_out0,v$A10A_16003_out0 };
assign v$_15017_out0 = { v$A9A_10415_out0,v$A10A_16006_out0 };
assign v$_16311_out0 = { v$C6_7056_out0,v$C7_16431_out0 };
assign v$_16314_out0 = { v$C6_7059_out0,v$C7_16434_out0 };
assign {v$A21_18570_out1,v$A21_18570_out0 } = v$A22_4426_out0 + v$B22_10807_out0 + v$C21_10769_out0;
assign v$G6_477_out0 = v$G4_11155_out0 || v$G7_9679_out0;
assign v$G6_486_out0 = v$G4_11164_out0 || v$G7_9688_out0;
assign v$G6_487_out0 = v$G4_11165_out0 || v$G7_9689_out0;
assign v$G6_498_out0 = v$G4_11176_out0 || v$G7_9700_out0;
assign v$G6_500_out0 = v$G4_11178_out0 || v$G7_9702_out0;
assign v$G6_507_out0 = v$G4_11185_out0 || v$G7_9709_out0;
assign v$G6_508_out0 = v$G4_11186_out0 || v$G7_9710_out0;
assign v$G6_600_out0 = v$G4_11278_out0 || v$G7_9802_out0;
assign v$G6_609_out0 = v$G4_11287_out0 || v$G7_9811_out0;
assign v$G6_610_out0 = v$G4_11288_out0 || v$G7_9812_out0;
assign v$G6_621_out0 = v$G4_11299_out0 || v$G7_9823_out0;
assign v$G6_623_out0 = v$G4_11301_out0 || v$G7_9825_out0;
assign v$G6_630_out0 = v$G4_11308_out0 || v$G7_9832_out0;
assign v$G6_631_out0 = v$G4_11309_out0 || v$G7_9833_out0;
assign v$_652_out0 = { v$C20_14980_out0,v$C21_6371_out0 };
assign v$_1578_out0 = { v$A21_18570_out0,v$A23_9548_out0 };
assign v$ENDs_3215_out0 = v$A21_18570_out1;
assign v$OP1_3381_out0 = v$OP1_14187_out0;
assign v$_7405_out0 = { v$_2454_out0,v$_16311_out0 };
assign v$_7408_out0 = { v$_2457_out0,v$_16314_out0 };
assign v$SUM$7_7743_out0 = v$SEL11_1500_out0;
assign v$ENDd_10834_out0 = v$A23_9548_out1;
assign v$_15710_out0 = { v$C22_8412_out0,v$C23_16151_out0 };
assign v$CIN_16814_out0 = v$CIN_3888_out0;
assign v$G$AD_17143_out0 = v$G4_11168_out0;
assign v$G$AD_17150_out0 = v$G4_11175_out0;
assign v$G$AD_17154_out0 = v$G4_11179_out0;
assign v$G$AD_17157_out0 = v$G4_11182_out0;
assign v$G$AD_17165_out0 = v$G4_11190_out0;
assign v$G$AD_17266_out0 = v$G4_11291_out0;
assign v$G$AD_17273_out0 = v$G4_11298_out0;
assign v$G$AD_17277_out0 = v$G4_11302_out0;
assign v$G$AD_17280_out0 = v$G4_11305_out0;
assign v$G$AD_17288_out0 = v$G4_11313_out0;
assign v$_17965_out0 = { v$_83_out0,v$_3637_out0 };
assign v$_17968_out0 = { v$_86_out0,v$_3640_out0 };
assign v$END32_2471_out0 = v$G$AD_17157_out0;
assign v$END32_2474_out0 = v$G$AD_17280_out0;
assign v$COUTD_6737_out0 = v$G6_477_out0;
assign v$COUTD_6746_out0 = v$G6_486_out0;
assign v$COUTD_6747_out0 = v$G6_487_out0;
assign v$COUTD_6758_out0 = v$G6_498_out0;
assign v$COUTD_6760_out0 = v$G6_500_out0;
assign v$COUTD_6767_out0 = v$G6_507_out0;
assign v$COUTD_6768_out0 = v$G6_508_out0;
assign v$COUTD_6860_out0 = v$G6_600_out0;
assign v$COUTD_6869_out0 = v$G6_609_out0;
assign v$COUTD_6870_out0 = v$G6_610_out0;
assign v$COUTD_6881_out0 = v$G6_621_out0;
assign v$COUTD_6883_out0 = v$G6_623_out0;
assign v$COUTD_6890_out0 = v$G6_630_out0;
assign v$COUTD_6891_out0 = v$G6_631_out0;
assign v$_7791_out0 = { v$_7254_out0,v$_7405_out0 };
assign v$_7794_out0 = { v$_7257_out0,v$_7408_out0 };
assign v$G$AB_9186_out0 = v$G$AD_17150_out0;
assign v$G$AB_9205_out0 = v$G$AD_17150_out0;
assign v$G$AB_9309_out0 = v$G$AD_17273_out0;
assign v$G$AB_9328_out0 = v$G$AD_17273_out0;
assign v$_9493_out0 = { v$_1795_out0,v$_1578_out0 };
assign v$END43_13193_out0 = v$G$AD_17165_out0;
assign v$END43_13196_out0 = v$G$AD_17288_out0;
assign v$_13734_out0 = { v$_652_out0,v$_15710_out0 };
assign v$END46_15046_out0 = v$G$AD_17150_out0;
assign v$END46_15049_out0 = v$G$AD_17273_out0;
assign v$END30_15714_out0 = v$G$AD_17154_out0;
assign v$END30_15717_out0 = v$G$AD_17277_out0;
assign v$END41_16666_out0 = v$G$AD_17143_out0;
assign v$END41_16669_out0 = v$G$AD_17266_out0;
assign v$SEL8_17653_out0 = v$OP1_3381_out0[23:1];
assign v$_17749_out0 = { v$_10356_out0,v$_17965_out0 };
assign v$_17752_out0 = { v$_10359_out0,v$_17968_out0 };
assign v$C14_280_out0 = v$COUTD_6758_out0;
assign v$C14_283_out0 = v$COUTD_6881_out0;
assign v$C17_2521_out0 = v$COUTD_6737_out0;
assign v$C17_2524_out0 = v$COUTD_6860_out0;
assign v$_4094_out0 = { v$_10351_out0,v$_13734_out0 };
assign v$G5_4569_out0 = v$G$AB_9186_out0 && v$P$CD_10504_out0;
assign v$G5_4588_out0 = v$G$AB_9205_out0 && v$P$CD_10523_out0;
assign v$G5_4692_out0 = v$G$AB_9309_out0 && v$P$CD_10627_out0;
assign v$G5_4711_out0 = v$G$AB_9328_out0 && v$P$CD_10646_out0;
assign v$C23_4844_out0 = v$COUTD_6760_out0;
assign v$C23_4847_out0 = v$COUTD_6883_out0;
assign v$C9_5938_out0 = v$COUTD_6747_out0;
assign v$C9_5941_out0 = v$COUTD_6870_out0;
assign v$_6660_out0 = { v$_16258_out0,v$_9493_out0 };
assign v$CINA_8521_out0 = v$COUTD_6737_out0;
assign v$CINA_8528_out0 = v$COUTD_6737_out0;
assign v$CINA_8532_out0 = v$COUTD_6758_out0;
assign v$CINA_8535_out0 = v$COUTD_6758_out0;
assign v$CINA_8543_out0 = v$COUTD_6737_out0;
assign v$CINA_8644_out0 = v$COUTD_6860_out0;
assign v$CINA_8651_out0 = v$COUTD_6860_out0;
assign v$CINA_8655_out0 = v$COUTD_6881_out0;
assign v$CINA_8658_out0 = v$COUTD_6881_out0;
assign v$CINA_8666_out0 = v$COUTD_6860_out0;
assign v$C13_11777_out0 = v$COUTD_6767_out0;
assign v$C13_11780_out0 = v$COUTD_6890_out0;
assign v$C10_12733_out0 = v$COUTD_6768_out0;
assign v$C10_12736_out0 = v$COUTD_6891_out0;
assign v$C12_13521_out0 = v$COUTD_6746_out0;
assign v$C12_13524_out0 = v$COUTD_6869_out0;
assign v$_17995_out0 = { v$SEL8_17653_out0,v$CIN_16814_out0 };
assign v$C14_326_out0 = v$C14_280_out0;
assign v$C14_329_out0 = v$C14_283_out0;
assign v$C10_1941_out0 = v$C10_12733_out0;
assign v$C10_1944_out0 = v$C10_12736_out0;
assign v$_3761_out0 = { v$_4869_out0,v$_4094_out0 };
assign {v$A12A_4446_out1,v$A12A_4446_out0 } = v$A11_9963_out0 + v$B11_9117_out0 + v$C10_12733_out0;
assign {v$A12A_4449_out1,v$A12A_4449_out0 } = v$A11_9966_out0 + v$B11_9120_out0 + v$C10_12736_out0;
assign v$C17_6067_out0 = v$C17_2521_out0;
assign v$C17_6070_out0 = v$C17_2524_out0;
assign {v$A13_7241_out1,v$A13_7241_out0 } = v$A15_17319_out0 + v$B15_10022_out0 + v$C14_280_out0;
assign {v$A13_7244_out1,v$A13_7244_out0 } = v$A15_17322_out0 + v$B15_10025_out0 + v$C14_283_out0;
assign v$C12_9395_out0 = v$C12_13521_out0;
assign v$C12_9398_out0 = v$C12_13524_out0;
assign v$_9908_out0 = { v$_18235_out0,v$_6660_out0 };
assign {v$A18_10033_out1,v$A18_10033_out0 } = v$A13_13863_out0 + v$B13_8676_out0 + v$C12_13521_out0;
assign {v$A18_10036_out1,v$A18_10036_out0 } = v$A13_13866_out0 + v$B13_8679_out0 + v$C12_13524_out0;
assign v$G4_11161_out0 = v$G5_4569_out0 || v$G$CD_964_out0;
assign v$G4_11180_out0 = v$G5_4588_out0 || v$G$CD_983_out0;
assign v$G4_11284_out0 = v$G5_4692_out0 || v$G$CD_1087_out0;
assign v$G4_11303_out0 = v$G5_4711_out0 || v$G$CD_1106_out0;
assign v$G8_11452_out0 = v$CINA_8521_out0 && v$P$AB_2058_out0;
assign v$G8_11459_out0 = v$CINA_8528_out0 && v$P$AB_2065_out0;
assign v$G8_11463_out0 = v$CINA_8532_out0 && v$P$AB_2069_out0;
assign v$G8_11466_out0 = v$CINA_8535_out0 && v$P$AB_2072_out0;
assign v$G8_11474_out0 = v$CINA_8543_out0 && v$P$AB_2080_out0;
assign v$G8_11575_out0 = v$CINA_8644_out0 && v$P$AB_2181_out0;
assign v$G8_11582_out0 = v$CINA_8651_out0 && v$P$AB_2188_out0;
assign v$G8_11586_out0 = v$CINA_8655_out0 && v$P$AB_2192_out0;
assign v$G8_11589_out0 = v$CINA_8658_out0 && v$P$AB_2195_out0;
assign v$G8_11597_out0 = v$CINA_8666_out0 && v$P$AB_2203_out0;
assign v$C9_12156_out0 = v$C9_5938_out0;
assign v$C9_12159_out0 = v$C9_5941_out0;
assign {v$A15_13217_out1,v$A15_13217_out0 } = v$A18_17696_out0 + v$B18_10868_out0 + v$C17_2521_out0;
assign {v$A15_13220_out1,v$A15_13220_out0 } = v$A18_17699_out0 + v$B18_10871_out0 + v$C17_2524_out0;
assign {v$A16A_14560_out1,v$A16A_14560_out0 } = v$A10_1549_out0 + v$B10_9878_out0 + v$C9_5938_out0;
assign {v$A16A_14563_out1,v$A16A_14563_out0 } = v$A10_1552_out0 + v$B10_9881_out0 + v$C9_5941_out0;
assign {v$A1_15216_out1,v$A1_15216_out0 } = v$_17995_out0 + v$MUX1_8340_out0 + v$C6_11352_out0;
assign v$C23_16150_out0 = v$C23_4844_out0;
assign v$C23_16153_out0 = v$C23_4847_out0;
assign {v$A20_16375_out1,v$A20_16375_out0 } = v$A14_677_out0 + v$B14_4003_out0 + v$C13_11777_out0;
assign {v$A20_16378_out1,v$A20_16378_out0 } = v$A14_680_out0 + v$B14_4006_out0 + v$C13_11780_out0;
assign v$C13_18590_out0 = v$C13_11777_out0;
assign v$C13_18593_out0 = v$C13_11780_out0;
assign v$ENDq_1459_out0 = v$A12A_4446_out1;
assign v$ENDq_1462_out0 = v$A12A_4449_out1;
assign v$_5897_out0 = { v$A17A_2488_out0,v$A18_10033_out0 };
assign v$_5900_out0 = { v$A17A_2491_out0,v$A18_10036_out0 };
assign v$CARRY_6333_out0 = v$C23_16150_out0;
assign v$CARRY_6336_out0 = v$C23_16153_out0;
assign v$ENDr_7523_out0 = v$A20_16375_out1;
assign v$ENDr_7526_out0 = v$A20_16378_out1;
assign v$_7553_out0 = { v$C8_18498_out0,v$C9_12156_out0 };
assign v$_7556_out0 = { v$C8_18501_out0,v$C9_12159_out0 };
assign v$COUT_8113_out0 = v$A1_15216_out1;
assign v$ENDi_8683_out0 = v$A15_13217_out1;
assign v$ENDi_8686_out0 = v$A15_13220_out1;
assign v$END0_9353_out0 = v$A16A_14560_out1;
assign v$END0_9356_out0 = v$A16A_14563_out1;
assign v$SUM_9364_out0 = v$_9908_out0;
assign v$G7_9692_out0 = v$G8_11452_out0 && v$P$CD_10511_out0;
assign v$G7_9699_out0 = v$G8_11459_out0 && v$P$CD_10518_out0;
assign v$G7_9703_out0 = v$G8_11463_out0 && v$P$CD_10522_out0;
assign v$G7_9706_out0 = v$G8_11466_out0 && v$P$CD_10525_out0;
assign v$G7_9714_out0 = v$G8_11474_out0 && v$P$CD_10533_out0;
assign v$G7_9815_out0 = v$G8_11575_out0 && v$P$CD_10634_out0;
assign v$G7_9822_out0 = v$G8_11582_out0 && v$P$CD_10641_out0;
assign v$G7_9826_out0 = v$G8_11586_out0 && v$P$CD_10645_out0;
assign v$G7_9829_out0 = v$G8_11589_out0 && v$P$CD_10648_out0;
assign v$G7_9837_out0 = v$G8_11597_out0 && v$P$CD_10656_out0;
assign v$_10238_out0 = { v$C12_9395_out0,v$C13_18590_out0 };
assign v$_10241_out0 = { v$C12_9398_out0,v$C13_18593_out0 };
assign v$ENDt_10259_out0 = v$A13_7241_out1;
assign v$ENDt_10262_out0 = v$A13_7244_out1;
assign v$_10959_out0 = { v$A16A_14560_out0,v$A12A_4446_out0 };
assign v$_10962_out0 = { v$A16A_14563_out0,v$A12A_4449_out0 };
assign v$SUM1_12829_out0 = v$_3761_out0;
assign v$_14837_out0 = { v$C10_1941_out0,v$C11_9511_out0 };
assign v$_14840_out0 = { v$C10_1944_out0,v$C11_9514_out0 };
assign v$SUM_15168_out0 = v$A1_15216_out0;
assign v$G$AD_17136_out0 = v$G4_11161_out0;
assign v$G$AD_17155_out0 = v$G4_11180_out0;
assign v$G$AD_17259_out0 = v$G4_11284_out0;
assign v$G$AD_17278_out0 = v$G4_11303_out0;
assign v$_17457_out0 = { v$A20_16375_out0,v$A13_7241_out0 };
assign v$_17460_out0 = { v$A20_16378_out0,v$A13_7244_out0 };
assign v$ENDe_17893_out0 = v$A18_10033_out1;
assign v$ENDe_17896_out0 = v$A18_10036_out1;
assign v$G6_490_out0 = v$G4_11168_out0 || v$G7_9692_out0;
assign v$G6_497_out0 = v$G4_11175_out0 || v$G7_9699_out0;
assign v$G6_501_out0 = v$G4_11179_out0 || v$G7_9703_out0;
assign v$G6_504_out0 = v$G4_11182_out0 || v$G7_9706_out0;
assign v$G6_512_out0 = v$G4_11190_out0 || v$G7_9714_out0;
assign v$G6_613_out0 = v$G4_11291_out0 || v$G7_9815_out0;
assign v$G6_620_out0 = v$G4_11298_out0 || v$G7_9822_out0;
assign v$G6_624_out0 = v$G4_11302_out0 || v$G7_9826_out0;
assign v$G6_627_out0 = v$G4_11305_out0 || v$G7_9829_out0;
assign v$G6_635_out0 = v$G4_11313_out0 || v$G7_9837_out0;
assign v$_1558_out0 = { v$_15014_out0,v$_10959_out0 };
assign v$_1561_out0 = { v$_15017_out0,v$_10962_out0 };
assign v$SUM_3468_out0 = v$SUM_15168_out0;
assign v$END50_7414_out0 = v$G$AD_17136_out0;
assign v$END50_7417_out0 = v$G$AD_17259_out0;
assign v$SEL4_7557_out0 = v$SUM_9364_out0[23:1];
assign v$END48_10366_out0 = v$G$AD_17155_out0;
assign v$END48_10369_out0 = v$G$AD_17278_out0;
assign v$COUT_10730_out0 = v$COUT_8113_out0;
assign v$IGNORE_12634_out0 = v$SUM1_12829_out0;
assign v$_14294_out0 = { v$_5897_out0,v$_17457_out0 };
assign v$_14297_out0 = { v$_5900_out0,v$_17460_out0 };
assign v$OVERFLOW_14976_out0 = v$CARRY_6333_out0;
assign v$OVERFLOW_14977_out0 = v$CARRY_6336_out0;
assign v$_18304_out0 = { v$_7553_out0,v$_14837_out0 };
assign v$_18307_out0 = { v$_7556_out0,v$_14840_out0 };
assign v$COUT$HALF_72_out0 = v$COUT_10730_out0;
assign v$OVERFLOW_426_out0 = v$OVERFLOW_14976_out0;
assign v$OVERFLOW_427_out0 = v$OVERFLOW_14977_out0;
assign v$_1174_out0 = { v$_1558_out0,v$_14294_out0 };
assign v$_1177_out0 = { v$_1561_out0,v$_14297_out0 };
assign v$SUM$HALF_2883_out0 = v$SUM_3468_out0;
assign v$SEL13_3883_out0 = v$SUM_3468_out0[0:0];
assign v$COUTD_6750_out0 = v$G6_490_out0;
assign v$COUTD_6757_out0 = v$G6_497_out0;
assign v$COUTD_6761_out0 = v$G6_501_out0;
assign v$COUTD_6764_out0 = v$G6_504_out0;
assign v$COUTD_6772_out0 = v$G6_512_out0;
assign v$COUTD_6873_out0 = v$G6_613_out0;
assign v$COUTD_6880_out0 = v$G6_620_out0;
assign v$COUTD_6884_out0 = v$G6_624_out0;
assign v$COUTD_6887_out0 = v$G6_627_out0;
assign v$COUTD_6895_out0 = v$G6_635_out0;
assign v$_7380_out0 = { v$SEL4_7557_out0,v$CARRY_6334_out0 };
assign v$C16_1269_out0 = v$COUTD_6764_out0;
assign v$C16_1272_out0 = v$COUTD_6887_out0;
assign v$FINAL$RESULT_2572_out0 = v$_7380_out0;
assign v$OVERFLOW_3630_out0 = v$OVERFLOW_426_out0;
assign v$OVERFLOW_3631_out0 = v$OVERFLOW_427_out0;
assign v$CIN_3890_out0 = v$COUT$HALF_72_out0;
assign v$C15_8144_out0 = v$COUTD_6761_out0;
assign v$C15_8147_out0 = v$COUTD_6884_out0;
assign v$C19_8161_out0 = v$COUTD_6772_out0;
assign v$C19_8164_out0 = v$COUTD_6895_out0;
assign v$CINA_8514_out0 = v$COUTD_6757_out0;
assign v$CINA_8533_out0 = v$COUTD_6757_out0;
assign v$CINA_8637_out0 = v$COUTD_6880_out0;
assign v$CINA_8656_out0 = v$COUTD_6880_out0;
assign v$OP1_14189_out0 = v$SUM$HALF_2883_out0;
assign v$C20_15490_out0 = v$COUTD_6757_out0;
assign v$C20_15493_out0 = v$COUTD_6880_out0;
assign v$SUM$8_15776_out0 = v$SEL13_3883_out0;
assign v$C18_16290_out0 = v$COUTD_6750_out0;
assign v$C18_16293_out0 = v$COUTD_6873_out0;
assign v$_18234_out0 = { v$_17749_out0,v$_1174_out0 };
assign v$_18237_out0 = { v$_17752_out0,v$_1177_out0 };
assign v$OP1_3383_out0 = v$OP1_14189_out0;
assign v$MULTIPLIER$OUT_9343_out0 = v$FINAL$RESULT_2572_out0;
assign v$G8_11445_out0 = v$CINA_8514_out0 && v$P$AB_2051_out0;
assign v$G8_11464_out0 = v$CINA_8533_out0 && v$P$AB_2070_out0;
assign v$G8_11568_out0 = v$CINA_8637_out0 && v$P$AB_2174_out0;
assign v$G8_11587_out0 = v$CINA_8656_out0 && v$P$AB_2193_out0;
assign v$C15_13132_out0 = v$C15_8144_out0;
assign v$C15_13135_out0 = v$C15_8147_out0;
assign v$C19_13834_out0 = v$C19_8161_out0;
assign v$C19_13837_out0 = v$C19_8164_out0;
assign v$C20_14979_out0 = v$C20_15490_out0;
assign v$C20_14982_out0 = v$C20_15493_out0;
assign v$C16_15158_out0 = v$C16_1269_out0;
assign v$C16_15161_out0 = v$C16_1272_out0;
assign {v$A14_15354_out1,v$A14_15354_out0 } = v$A16_13615_out0 + v$B16_16415_out0 + v$C15_8144_out0;
assign {v$A14_15357_out1,v$A14_15357_out0 } = v$A16_13618_out0 + v$B16_16418_out0 + v$C15_8147_out0;
assign {v$A19_15909_out1,v$A19_15909_out0 } = v$A19_1214_out0 + v$B19_16790_out0 + v$C18_16290_out0;
assign {v$A19_15912_out1,v$A19_15912_out0 } = v$A19_1217_out0 + v$B19_16793_out0 + v$C18_16293_out0;
assign v$CIN_16816_out0 = v$CIN_3890_out0;
assign {v$A24_16974_out1,v$A24_16974_out0 } = v$A21_2599_out0 + v$B21_18083_out0 + v$C20_15490_out0;
assign {v$A24_16977_out1,v$A24_16977_out0 } = v$A21_2602_out0 + v$B21_18086_out0 + v$C20_15493_out0;
assign {v$A22_17489_out1,v$A22_17489_out0 } = v$A20_4437_out0 + v$B20_3944_out0 + v$C19_8161_out0;
assign {v$A22_17492_out1,v$A22_17492_out0 } = v$A20_4440_out0 + v$B20_3947_out0 + v$C19_8164_out0;
assign {v$A11_17875_out1,v$A11_17875_out0 } = v$A17_16723_out0 + v$B17_15536_out0 + v$C16_1269_out0;
assign {v$A11_17878_out1,v$A11_17878_out0 } = v$A17_16726_out0 + v$B17_15539_out0 + v$C16_1272_out0;
assign v$C18_18006_out0 = v$C18_16290_out0;
assign v$C18_18009_out0 = v$C18_16293_out0;
assign v$OVERFLOW_18455_out0 = v$OVERFLOW_3630_out0;
assign v$OVERFLOW_18456_out0 = v$OVERFLOW_3631_out0;
assign v$OVERFLOW_18525_out0 = v$OVERFLOW_3630_out0;
assign v$OVERFLOW_18526_out0 = v$OVERFLOW_3631_out0;
assign v$_1200_out0 = { v$A15_13217_out0,v$A19_15909_out0 };
assign v$_1203_out0 = { v$A15_13220_out0,v$A19_15912_out0 };
assign v$_1794_out0 = { v$A22_17489_out0,v$A24_16974_out0 };
assign v$_1797_out0 = { v$A22_17492_out0,v$A24_16977_out0 };
assign v$_2841_out0 = { v$C14_326_out0,v$C15_13132_out0 };
assign v$_2844_out0 = { v$C14_329_out0,v$C15_13135_out0 };
assign v$ENDp_3190_out0 = v$A22_17489_out1;
assign v$ENDp_3193_out0 = v$A22_17492_out1;
assign v$ENDy_4115_out0 = v$A14_15354_out1;
assign v$ENDy_4118_out0 = v$A14_15357_out1;
assign v$ENDu_7030_out0 = v$A11_17875_out1;
assign v$ENDu_7033_out0 = v$A11_17878_out1;
assign v$_7869_out0 = { v$C16_15158_out0,v$C17_6067_out0 };
assign v$_7872_out0 = { v$C16_15161_out0,v$C17_6070_out0 };
assign v$_8330_out0 = { v$C18_18006_out0,v$C19_13834_out0 };
assign v$_8333_out0 = { v$C18_18009_out0,v$C19_13837_out0 };
assign v$G7_9685_out0 = v$G8_11445_out0 && v$P$CD_10504_out0;
assign v$G7_9704_out0 = v$G8_11464_out0 && v$P$CD_10523_out0;
assign v$G7_9808_out0 = v$G8_11568_out0 && v$P$CD_10627_out0;
assign v$G7_9827_out0 = v$G8_11587_out0 && v$P$CD_10646_out0;
assign v$IN_11071_out0 = v$MULTIPLIER$OUT_9343_out0;
assign v$IN_11072_out0 = v$MULTIPLIER$OUT_9343_out0;
assign {v$A1_11802_out1,v$A1_11802_out0 } = v$C1_7424_out0 + v$EXPONENT_16011_out0 + v$OVERFLOW_18525_out0;
assign {v$A1_11803_out1,v$A1_11803_out0 } = v$C1_7425_out0 + v$EXPONENT_16012_out0 + v$OVERFLOW_18526_out0;
assign v$_13294_out0 = { v$A14_15354_out0,v$A11_17875_out0 };
assign v$_13297_out0 = { v$A14_15357_out0,v$A11_17878_out0 };
assign {v$A1_15763_out1,v$A1_15763_out0 } = v$C1_13991_out0 + v$EXPONENT_13686_out0 + v$OVERFLOW_18455_out0;
assign {v$A1_15764_out1,v$A1_15764_out0 } = v$C1_13992_out0 + v$EXPONENT_13687_out0 + v$OVERFLOW_18456_out0;
assign v$ENDa_16565_out0 = v$A24_16974_out1;
assign v$ENDa_16568_out0 = v$A24_16977_out1;
assign v$SEL8_17655_out0 = v$OP1_3383_out0[23:1];
assign v$ENDo_18693_out0 = v$A19_15909_out1;
assign v$ENDo_18696_out0 = v$A19_15912_out1;
assign v$OUT_170_out0 = v$A1_11802_out0;
assign v$OUT_171_out0 = v$A1_11803_out0;
assign v$G6_483_out0 = v$G4_11161_out0 || v$G7_9685_out0;
assign v$G6_502_out0 = v$G4_11180_out0 || v$G7_9704_out0;
assign v$G6_606_out0 = v$G4_11284_out0 || v$G7_9808_out0;
assign v$G6_625_out0 = v$G4_11303_out0 || v$G7_9827_out0;
assign v$_1243_out0 = { v$_10238_out0,v$_2841_out0 };
assign v$_1246_out0 = { v$_10241_out0,v$_2844_out0 };
assign v$NOT$USED_2891_out0 = v$A1_11802_out1;
assign v$NOT$USED_2892_out0 = v$A1_11803_out1;
assign v$NOT$USED_5449_out0 = v$A1_15763_out1;
assign v$NOT$USED_5450_out0 = v$A1_15764_out1;
assign v$_10350_out0 = { v$_7869_out0,v$_8330_out0 };
assign v$_10353_out0 = { v$_7872_out0,v$_8333_out0 };
assign v$IN_11642_out0 = v$IN_11071_out0;
assign v$IN_11643_out0 = v$IN_11072_out0;
assign v$OUT_14778_out0 = v$A1_15763_out0;
assign v$OUT_14779_out0 = v$A1_15764_out0;
assign v$_16257_out0 = { v$_13294_out0,v$_1200_out0 };
assign v$_16260_out0 = { v$_13297_out0,v$_1203_out0 };
assign v$_17997_out0 = { v$SEL8_17655_out0,v$CIN_16816_out0 };
assign v$COUTD_6743_out0 = v$G6_483_out0;
assign v$COUTD_6762_out0 = v$G6_502_out0;
assign v$COUTD_6866_out0 = v$G6_606_out0;
assign v$COUTD_6885_out0 = v$G6_625_out0;
assign v$IN_8294_out0 = v$IN_11642_out0;
assign v$IN_8295_out0 = v$IN_11643_out0;
assign v$IN_13562_out0 = v$IN_11642_out0;
assign v$IN_13564_out0 = v$IN_11643_out0;
assign {v$A1_15218_out1,v$A1_15218_out0 } = v$_17997_out0 + v$MUX1_8342_out0 + v$C6_11354_out0;
assign v$_17354_out0 = { v$_18304_out0,v$_1243_out0 };
assign v$_17357_out0 = { v$_18307_out0,v$_1246_out0 };
assign v$IN_18262_out0 = v$IN_11642_out0;
assign v$IN_18263_out0 = v$IN_11643_out0;
assign v$IN_4190_out0 = v$IN_8294_out0;
assign v$IN_4191_out0 = v$IN_8295_out0;
assign v$_4868_out0 = { v$_7791_out0,v$_17354_out0 };
assign v$_4871_out0 = { v$_7794_out0,v$_17357_out0 };
assign v$IN_5162_out0 = v$IN_18262_out0;
assign v$IN_5172_out0 = v$IN_18263_out0;
assign v$SEL2_6393_out0 = v$IN_13562_out0[23:8];
assign v$SEL2_6394_out0 = v$IN_13564_out0[23:8];
assign v$COUT_8115_out0 = v$A1_15218_out1;
assign v$C21_10768_out0 = v$COUTD_6762_out0;
assign v$C21_10771_out0 = v$COUTD_6885_out0;
assign v$C22_10982_out0 = v$COUTD_6743_out0;
assign v$C22_10985_out0 = v$COUTD_6866_out0;
assign v$SUM_15170_out0 = v$A1_15218_out0;
assign v$SEL1_16684_out0 = v$IN_13562_out0[7:0];
assign v$SEL1_16686_out0 = v$IN_13564_out0[7:0];
assign v$SUM_3470_out0 = v$SUM_15170_out0;
assign v$IN_3859_out0 = v$IN_5162_out0;
assign v$IN_3862_out0 = v$IN_5172_out0;
assign v$SEL15_4886_out0 = v$IN_4190_out0[9:9];
assign v$SEL15_4887_out0 = v$IN_4191_out0[9:9];
assign v$C21_6370_out0 = v$C21_10768_out0;
assign v$C21_6373_out0 = v$C21_10771_out0;
assign v$SEL13_6924_out0 = v$IN_4190_out0[11:11];
assign v$SEL13_6925_out0 = v$IN_4191_out0[11:11];
assign v$SEL1_7088_out0 = v$IN_4190_out0[23:23];
assign v$SEL1_7089_out0 = v$IN_4191_out0[23:23];
assign v$SEL11_7225_out0 = v$IN_4190_out0[13:13];
assign v$SEL11_7226_out0 = v$IN_4191_out0[13:13];
assign v$SEL4_7321_out0 = v$IN_4190_out0[20:20];
assign v$SEL4_7322_out0 = v$IN_4191_out0[20:20];
assign v$SEL22_7397_out0 = v$IN_4190_out0[2:2];
assign v$SEL22_7398_out0 = v$IN_4191_out0[2:2];
assign v$SEL23_7617_out0 = v$IN_4190_out0[1:1];
assign v$SEL23_7618_out0 = v$IN_4191_out0[1:1];
assign v$SEL20_8174_out0 = v$IN_4190_out0[4:4];
assign v$SEL20_8175_out0 = v$IN_4191_out0[4:4];
assign v$C22_8411_out0 = v$C22_10982_out0;
assign v$C22_8414_out0 = v$C22_10985_out0;
assign v$SEL10_9506_out0 = v$IN_4190_out0[16:16];
assign v$SEL10_9507_out0 = v$IN_4191_out0[16:16];
assign {v$A23_9547_out1,v$A23_9547_out0 } = v$A23_5064_out0 + v$B23_1284_out0 + v$C22_10982_out0;
assign {v$A23_9550_out1,v$A23_9550_out0 } = v$A23_5067_out0 + v$B23_1287_out0 + v$C22_10985_out0;
assign v$SEL9_10263_out0 = v$IN_4190_out0[14:14];
assign v$SEL9_10264_out0 = v$IN_4191_out0[14:14];
assign v$COUT_10732_out0 = v$COUT_8115_out0;
assign v$SEL21_11048_out0 = v$IN_4190_out0[3:3];
assign v$SEL21_11049_out0 = v$IN_4191_out0[3:3];
assign v$SEL18_11379_out0 = v$IN_4190_out0[6:6];
assign v$SEL18_11380_out0 = v$IN_4191_out0[6:6];
assign v$SEL3_11729_out0 = v$IN_4190_out0[21:21];
assign v$SEL3_11730_out0 = v$IN_4191_out0[21:21];
assign v$SEL6_12472_out0 = v$IN_4190_out0[18:18];
assign v$SEL6_12473_out0 = v$IN_4191_out0[18:18];
assign v$SEL19_12815_out0 = v$IN_4190_out0[5:5];
assign v$SEL19_12816_out0 = v$IN_4191_out0[5:5];
assign v$SEL2_13321_out0 = v$IN_4190_out0[22:22];
assign v$SEL2_13322_out0 = v$IN_4191_out0[22:22];
assign v$IN_13563_out0 = v$SEL2_6393_out0;
assign v$IN_13565_out0 = v$SEL2_6394_out0;
assign v$SEL12_13844_out0 = v$IN_4190_out0[12:12];
assign v$SEL12_13845_out0 = v$IN_4191_out0[12:12];
assign v$SEL7_14332_out0 = v$IN_4190_out0[17:17];
assign v$SEL7_14333_out0 = v$IN_4191_out0[17:17];
assign v$IN_14857_out0 = v$SEL1_16684_out0;
assign v$IN_14858_out0 = v$SEL1_16686_out0;
assign v$SEL5_15451_out0 = v$IN_4190_out0[19:19];
assign v$SEL5_15452_out0 = v$IN_4191_out0[19:19];
assign v$SEL17_16069_out0 = v$IN_4190_out0[7:7];
assign v$SEL17_16070_out0 = v$IN_4191_out0[7:7];
assign v$SEL14_16347_out0 = v$IN_4190_out0[10:10];
assign v$SEL14_16348_out0 = v$IN_4191_out0[10:10];
assign v$SEL16_16894_out0 = v$IN_4190_out0[8:8];
assign v$SEL16_16895_out0 = v$IN_4191_out0[8:8];
assign v$SEL24_16922_out0 = v$IN_4190_out0[0:0];
assign v$SEL24_16923_out0 = v$IN_4191_out0[0:0];
assign v$SEL8_17683_out0 = v$IN_4190_out0[15:15];
assign v$SEL8_17684_out0 = v$IN_4191_out0[15:15];
assign {v$A21_18569_out1,v$A21_18569_out0 } = v$A22_4425_out0 + v$B22_10806_out0 + v$C21_10768_out0;
assign {v$A21_18572_out1,v$A21_18572_out0 } = v$A22_4428_out0 + v$B22_10809_out0 + v$C21_10771_out0;
assign v$_651_out0 = { v$C20_14979_out0,v$C21_6370_out0 };
assign v$_654_out0 = { v$C20_14982_out0,v$C21_6373_out0 };
assign v$SEL12_1516_out0 = v$SUM_3470_out0[0:0];
assign v$_1577_out0 = { v$A21_18569_out0,v$A23_9547_out0 };
assign v$_1580_out0 = { v$A21_18572_out0,v$A23_9550_out0 };
assign v$SEL2_3027_out0 = v$IN_14857_out0[7:4];
assign v$SEL2_3028_out0 = v$IN_14858_out0[7:4];
assign v$ENDs_3214_out0 = v$A21_18569_out1;
assign v$ENDs_3217_out0 = v$A21_18572_out1;
assign v$SEL4_3368_out0 = v$IN_13563_out0[15:12];
assign v$SEL4_3369_out0 = v$IN_13565_out0[15:12];
assign v$CIN_3889_out0 = v$COUT_10732_out0;
assign v$SEL3_7364_out0 = v$IN_13563_out0[11:8];
assign v$SEL3_7365_out0 = v$IN_13565_out0[11:8];
assign v$SEL1_8710_out0 = v$IN_3859_out0[23:1];
assign v$SEL1_8720_out0 = v$IN_3862_out0[23:1];
assign v$ENDd_10833_out0 = v$A23_9547_out1;
assign v$ENDd_10836_out0 = v$A23_9550_out1;
assign v$SEL2_13850_out0 = v$IN_13563_out0[7:4];
assign v$SEL2_13851_out0 = v$IN_13565_out0[7:4];
assign v$OP1_14188_out0 = v$SUM_3470_out0;
assign v$SEL1_15401_out0 = v$IN_3859_out0[22:0];
assign v$SEL1_15411_out0 = v$IN_3862_out0[22:0];
assign v$_15709_out0 = { v$C22_8411_out0,v$C23_16150_out0 };
assign v$_15712_out0 = { v$C22_8414_out0,v$C23_16153_out0 };
assign v$SEL1_16458_out0 = v$IN_14857_out0[3:0];
assign v$SEL1_16459_out0 = v$IN_14858_out0[3:0];
assign v$SEL1_16685_out0 = v$IN_13563_out0[3:0];
assign v$SEL1_16687_out0 = v$IN_13565_out0[3:0];
assign v$MUX24_18056_out0 = v$EQ24_2536_out0 ? v$SEL24_16922_out0 : v$C1_15720_out0;
assign v$MUX24_18057_out0 = v$EQ24_2537_out0 ? v$SEL24_16923_out0 : v$C1_15721_out0;
assign v$SUM$9_197_out0 = v$SEL12_1516_out0;
assign v$OP1_3382_out0 = v$OP1_14188_out0;
assign v$_4260_out0 = { v$C2_118_out0,v$SEL1_15401_out0 };
assign v$_4270_out0 = { v$C2_128_out0,v$SEL1_15411_out0 };
assign v$_8995_out0 = { v$SEL1_8710_out0,v$C1_5976_out0 };
assign v$_9005_out0 = { v$SEL1_8720_out0,v$C1_5986_out0 };
assign v$_9492_out0 = { v$_1794_out0,v$_1577_out0 };
assign v$_9495_out0 = { v$_1797_out0,v$_1580_out0 };
assign v$_13733_out0 = { v$_651_out0,v$_15709_out0 };
assign v$_13736_out0 = { v$_654_out0,v$_15712_out0 };
assign v$IN_15063_out0 = v$SEL3_7364_out0;
assign v$IN_15064_out0 = v$SEL1_16685_out0;
assign v$IN_15065_out0 = v$SEL2_13850_out0;
assign v$IN_15066_out0 = v$SEL4_3368_out0;
assign v$IN_15067_out0 = v$SEL1_16458_out0;
assign v$IN_15068_out0 = v$SEL2_3027_out0;
assign v$IN_15069_out0 = v$SEL3_7365_out0;
assign v$IN_15070_out0 = v$SEL1_16687_out0;
assign v$IN_15071_out0 = v$SEL2_13851_out0;
assign v$IN_15072_out0 = v$SEL4_3369_out0;
assign v$IN_15073_out0 = v$SEL1_16459_out0;
assign v$IN_15074_out0 = v$SEL2_3028_out0;
assign v$MUX23_16223_out0 = v$EQ23_3194_out0 ? v$SEL23_7617_out0 : v$MUX24_18056_out0;
assign v$MUX23_16224_out0 = v$EQ23_3195_out0 ? v$SEL23_7618_out0 : v$MUX24_18057_out0;
assign v$CIN_16815_out0 = v$CIN_3889_out0;
assign v$SEL3_2300_out0 = v$IN_15063_out0[2:2];
assign v$SEL3_2301_out0 = v$IN_15064_out0[2:2];
assign v$SEL3_2302_out0 = v$IN_15065_out0[2:2];
assign v$SEL3_2303_out0 = v$IN_15066_out0[2:2];
assign v$SEL3_2304_out0 = v$IN_15067_out0[2:2];
assign v$SEL3_2305_out0 = v$IN_15068_out0[2:2];
assign v$SEL3_2306_out0 = v$IN_15069_out0[2:2];
assign v$SEL3_2307_out0 = v$IN_15070_out0[2:2];
assign v$SEL3_2308_out0 = v$IN_15071_out0[2:2];
assign v$SEL3_2309_out0 = v$IN_15072_out0[2:2];
assign v$SEL3_2310_out0 = v$IN_15073_out0[2:2];
assign v$SEL3_2311_out0 = v$IN_15074_out0[2:2];
assign v$MUX1_2364_out0 = v$LEFT$SHIT_3056_out0 ? v$_4260_out0 : v$_8995_out0;
assign v$MUX1_2374_out0 = v$LEFT$SHIT_3066_out0 ? v$_4270_out0 : v$_9005_out0;
assign v$_4093_out0 = { v$_10350_out0,v$_13733_out0 };
assign v$_4096_out0 = { v$_10353_out0,v$_13736_out0 };
assign v$SEL4_6085_out0 = v$IN_15063_out0[3:3];
assign v$SEL4_6086_out0 = v$IN_15064_out0[3:3];
assign v$SEL4_6087_out0 = v$IN_15065_out0[3:3];
assign v$SEL4_6088_out0 = v$IN_15066_out0[3:3];
assign v$SEL4_6089_out0 = v$IN_15067_out0[3:3];
assign v$SEL4_6090_out0 = v$IN_15068_out0[3:3];
assign v$SEL4_6091_out0 = v$IN_15069_out0[3:3];
assign v$SEL4_6092_out0 = v$IN_15070_out0[3:3];
assign v$SEL4_6093_out0 = v$IN_15071_out0[3:3];
assign v$SEL4_6094_out0 = v$IN_15072_out0[3:3];
assign v$SEL4_6095_out0 = v$IN_15073_out0[3:3];
assign v$SEL4_6096_out0 = v$IN_15074_out0[3:3];
assign v$_6659_out0 = { v$_16257_out0,v$_9492_out0 };
assign v$_6662_out0 = { v$_16260_out0,v$_9495_out0 };
assign v$SEL2_7676_out0 = v$IN_15063_out0[1:1];
assign v$SEL2_7677_out0 = v$IN_15064_out0[1:1];
assign v$SEL2_7678_out0 = v$IN_15065_out0[1:1];
assign v$SEL2_7679_out0 = v$IN_15066_out0[1:1];
assign v$SEL2_7680_out0 = v$IN_15067_out0[1:1];
assign v$SEL2_7681_out0 = v$IN_15068_out0[1:1];
assign v$SEL2_7682_out0 = v$IN_15069_out0[1:1];
assign v$SEL2_7683_out0 = v$IN_15070_out0[1:1];
assign v$SEL2_7684_out0 = v$IN_15071_out0[1:1];
assign v$SEL2_7685_out0 = v$IN_15072_out0[1:1];
assign v$SEL2_7686_out0 = v$IN_15073_out0[1:1];
assign v$SEL2_7687_out0 = v$IN_15074_out0[1:1];
assign v$SEL1_13465_out0 = v$IN_15063_out0[0:0];
assign v$SEL1_13466_out0 = v$IN_15064_out0[0:0];
assign v$SEL1_13467_out0 = v$IN_15065_out0[0:0];
assign v$SEL1_13468_out0 = v$IN_15066_out0[0:0];
assign v$SEL1_13469_out0 = v$IN_15067_out0[0:0];
assign v$SEL1_13470_out0 = v$IN_15068_out0[0:0];
assign v$SEL1_13471_out0 = v$IN_15069_out0[0:0];
assign v$SEL1_13472_out0 = v$IN_15070_out0[0:0];
assign v$SEL1_13473_out0 = v$IN_15071_out0[0:0];
assign v$SEL1_13474_out0 = v$IN_15072_out0[0:0];
assign v$SEL1_13475_out0 = v$IN_15073_out0[0:0];
assign v$SEL1_13476_out0 = v$IN_15074_out0[0:0];
assign v$MUX22_16464_out0 = v$EQ22_2836_out0 ? v$SEL22_7397_out0 : v$MUX23_16223_out0;
assign v$MUX22_16465_out0 = v$EQ22_2837_out0 ? v$SEL22_7398_out0 : v$MUX23_16224_out0;
assign v$SEL8_17654_out0 = v$OP1_3382_out0[23:1];
assign v$G10_1386_out0 = !(v$SEL1_13465_out0 || v$SEL2_7676_out0);
assign v$G10_1387_out0 = !(v$SEL1_13466_out0 || v$SEL2_7677_out0);
assign v$G10_1388_out0 = !(v$SEL1_13467_out0 || v$SEL2_7678_out0);
assign v$G10_1389_out0 = !(v$SEL1_13468_out0 || v$SEL2_7679_out0);
assign v$G10_1390_out0 = !(v$SEL1_13469_out0 || v$SEL2_7680_out0);
assign v$G10_1391_out0 = !(v$SEL1_13470_out0 || v$SEL2_7681_out0);
assign v$G10_1392_out0 = !(v$SEL1_13471_out0 || v$SEL2_7682_out0);
assign v$G10_1393_out0 = !(v$SEL1_13472_out0 || v$SEL2_7683_out0);
assign v$G10_1394_out0 = !(v$SEL1_13473_out0 || v$SEL2_7684_out0);
assign v$G10_1395_out0 = !(v$SEL1_13474_out0 || v$SEL2_7685_out0);
assign v$G10_1396_out0 = !(v$SEL1_13475_out0 || v$SEL2_7686_out0);
assign v$G10_1397_out0 = !(v$SEL1_13476_out0 || v$SEL2_7687_out0);
assign v$G6_3561_out0 = ! v$SEL2_7676_out0;
assign v$G6_3562_out0 = ! v$SEL2_7677_out0;
assign v$G6_3563_out0 = ! v$SEL2_7678_out0;
assign v$G6_3564_out0 = ! v$SEL2_7679_out0;
assign v$G6_3565_out0 = ! v$SEL2_7680_out0;
assign v$G6_3566_out0 = ! v$SEL2_7681_out0;
assign v$G6_3567_out0 = ! v$SEL2_7682_out0;
assign v$G6_3568_out0 = ! v$SEL2_7683_out0;
assign v$G6_3569_out0 = ! v$SEL2_7684_out0;
assign v$G6_3570_out0 = ! v$SEL2_7685_out0;
assign v$G6_3571_out0 = ! v$SEL2_7686_out0;
assign v$G6_3572_out0 = ! v$SEL2_7687_out0;
assign v$_3760_out0 = { v$_4868_out0,v$_4093_out0 };
assign v$_3763_out0 = { v$_4871_out0,v$_4096_out0 };
assign v$MUX21_4902_out0 = v$EQ21_3324_out0 ? v$SEL21_11048_out0 : v$MUX22_16464_out0;
assign v$MUX21_4903_out0 = v$EQ21_3325_out0 ? v$SEL21_11049_out0 : v$MUX22_16465_out0;
assign v$G5_5837_out0 = ! v$SEL4_6085_out0;
assign v$G5_5838_out0 = ! v$SEL4_6086_out0;
assign v$G5_5839_out0 = ! v$SEL4_6087_out0;
assign v$G5_5840_out0 = ! v$SEL4_6088_out0;
assign v$G5_5841_out0 = ! v$SEL4_6089_out0;
assign v$G5_5842_out0 = ! v$SEL4_6090_out0;
assign v$G5_5843_out0 = ! v$SEL4_6091_out0;
assign v$G5_5844_out0 = ! v$SEL4_6092_out0;
assign v$G5_5845_out0 = ! v$SEL4_6093_out0;
assign v$G5_5846_out0 = ! v$SEL4_6094_out0;
assign v$G5_5847_out0 = ! v$SEL4_6095_out0;
assign v$G5_5848_out0 = ! v$SEL4_6096_out0;
assign v$G11_8848_out0 = !(v$SEL3_2300_out0 || v$SEL4_6085_out0);
assign v$G11_8849_out0 = !(v$SEL3_2301_out0 || v$SEL4_6086_out0);
assign v$G11_8850_out0 = !(v$SEL3_2302_out0 || v$SEL4_6087_out0);
assign v$G11_8851_out0 = !(v$SEL3_2303_out0 || v$SEL4_6088_out0);
assign v$G11_8852_out0 = !(v$SEL3_2304_out0 || v$SEL4_6089_out0);
assign v$G11_8853_out0 = !(v$SEL3_2305_out0 || v$SEL4_6090_out0);
assign v$G11_8854_out0 = !(v$SEL3_2306_out0 || v$SEL4_6091_out0);
assign v$G11_8855_out0 = !(v$SEL3_2307_out0 || v$SEL4_6092_out0);
assign v$G11_8856_out0 = !(v$SEL3_2308_out0 || v$SEL4_6093_out0);
assign v$G11_8857_out0 = !(v$SEL3_2309_out0 || v$SEL4_6094_out0);
assign v$G11_8858_out0 = !(v$SEL3_2310_out0 || v$SEL4_6095_out0);
assign v$G11_8859_out0 = !(v$SEL3_2311_out0 || v$SEL4_6096_out0);
assign v$_9907_out0 = { v$_18234_out0,v$_6659_out0 };
assign v$_9910_out0 = { v$_18237_out0,v$_6662_out0 };
assign v$G8_11996_out0 = ! v$SEL3_2300_out0;
assign v$G8_11997_out0 = ! v$SEL3_2301_out0;
assign v$G8_11998_out0 = ! v$SEL3_2302_out0;
assign v$G8_11999_out0 = ! v$SEL3_2303_out0;
assign v$G8_12000_out0 = ! v$SEL3_2304_out0;
assign v$G8_12001_out0 = ! v$SEL3_2305_out0;
assign v$G8_12002_out0 = ! v$SEL3_2306_out0;
assign v$G8_12003_out0 = ! v$SEL3_2307_out0;
assign v$G8_12004_out0 = ! v$SEL3_2308_out0;
assign v$G8_12005_out0 = ! v$SEL3_2309_out0;
assign v$G8_12006_out0 = ! v$SEL3_2310_out0;
assign v$G8_12007_out0 = ! v$SEL3_2311_out0;
assign v$_17996_out0 = { v$SEL8_17654_out0,v$CIN_16815_out0 };
assign v$SUM_9363_out0 = v$_9907_out0;
assign v$SUM_9366_out0 = v$_9910_out0;
assign v$MUX20_11364_out0 = v$EQ20_9946_out0 ? v$SEL20_8174_out0 : v$MUX21_4902_out0;
assign v$MUX20_11365_out0 = v$EQ20_9947_out0 ? v$SEL20_8175_out0 : v$MUX21_4903_out0;
assign v$G3_12668_out0 = v$G10_1386_out0 && v$G11_8848_out0;
assign v$G3_12669_out0 = v$G10_1387_out0 && v$G11_8849_out0;
assign v$G3_12670_out0 = v$G10_1388_out0 && v$G11_8850_out0;
assign v$G3_12671_out0 = v$G10_1389_out0 && v$G11_8851_out0;
assign v$G3_12672_out0 = v$G10_1390_out0 && v$G11_8852_out0;
assign v$G3_12673_out0 = v$G10_1391_out0 && v$G11_8853_out0;
assign v$G3_12674_out0 = v$G10_1392_out0 && v$G11_8854_out0;
assign v$G3_12675_out0 = v$G10_1393_out0 && v$G11_8855_out0;
assign v$G3_12676_out0 = v$G10_1394_out0 && v$G11_8856_out0;
assign v$G3_12677_out0 = v$G10_1395_out0 && v$G11_8857_out0;
assign v$G3_12678_out0 = v$G10_1396_out0 && v$G11_8858_out0;
assign v$G3_12679_out0 = v$G10_1397_out0 && v$G11_8859_out0;
assign v$SUM1_12828_out0 = v$_3760_out0;
assign v$SUM1_12831_out0 = v$_3763_out0;
assign {v$A1_15217_out1,v$A1_15217_out0 } = v$_17996_out0 + v$MUX1_8341_out0 + v$C6_11353_out0;
assign v$G9_17594_out0 = v$G8_11996_out0 && v$G5_5837_out0;
assign v$G9_17595_out0 = v$G8_11997_out0 && v$G5_5838_out0;
assign v$G9_17596_out0 = v$G8_11998_out0 && v$G5_5839_out0;
assign v$G9_17597_out0 = v$G8_11999_out0 && v$G5_5840_out0;
assign v$G9_17598_out0 = v$G8_12000_out0 && v$G5_5841_out0;
assign v$G9_17599_out0 = v$G8_12001_out0 && v$G5_5842_out0;
assign v$G9_17600_out0 = v$G8_12002_out0 && v$G5_5843_out0;
assign v$G9_17601_out0 = v$G8_12003_out0 && v$G5_5844_out0;
assign v$G9_17602_out0 = v$G8_12004_out0 && v$G5_5845_out0;
assign v$G9_17603_out0 = v$G8_12005_out0 && v$G5_5846_out0;
assign v$G9_17604_out0 = v$G8_12006_out0 && v$G5_5847_out0;
assign v$G9_17605_out0 = v$G8_12007_out0 && v$G5_5848_out0;
assign v$G7_18137_out0 = v$G6_3561_out0 || v$SEL3_2300_out0;
assign v$G7_18138_out0 = v$G6_3562_out0 || v$SEL3_2301_out0;
assign v$G7_18139_out0 = v$G6_3563_out0 || v$SEL3_2302_out0;
assign v$G7_18140_out0 = v$G6_3564_out0 || v$SEL3_2303_out0;
assign v$G7_18141_out0 = v$G6_3565_out0 || v$SEL3_2304_out0;
assign v$G7_18142_out0 = v$G6_3566_out0 || v$SEL3_2305_out0;
assign v$G7_18143_out0 = v$G6_3567_out0 || v$SEL3_2306_out0;
assign v$G7_18144_out0 = v$G6_3568_out0 || v$SEL3_2307_out0;
assign v$G7_18145_out0 = v$G6_3569_out0 || v$SEL3_2308_out0;
assign v$G7_18146_out0 = v$G6_3570_out0 || v$SEL3_2309_out0;
assign v$G7_18147_out0 = v$G6_3571_out0 || v$SEL3_2310_out0;
assign v$G7_18148_out0 = v$G6_3572_out0 || v$SEL3_2311_out0;
assign v$SUM_1905_out0 = v$SUM_9363_out0;
assign v$SUM_1906_out0 = v$SUM_9366_out0;
assign v$MUX19_6374_out0 = v$EQ19_5442_out0 ? v$SEL19_12815_out0 : v$MUX20_11364_out0;
assign v$MUX19_6375_out0 = v$EQ19_5443_out0 ? v$SEL19_12816_out0 : v$MUX20_11365_out0;
assign v$COUT_8114_out0 = v$A1_15217_out1;
assign v$END1_9929_out0 = v$SUM1_12828_out0;
assign v$END1_9930_out0 = v$SUM1_12831_out0;
assign v$Z_12559_out0 = v$G3_12668_out0;
assign v$Z_12560_out0 = v$G3_12669_out0;
assign v$Z_12561_out0 = v$G3_12670_out0;
assign v$Z_12562_out0 = v$G3_12671_out0;
assign v$Z_12563_out0 = v$G3_12672_out0;
assign v$Z_12564_out0 = v$G3_12673_out0;
assign v$Z_12565_out0 = v$G3_12674_out0;
assign v$Z_12566_out0 = v$G3_12675_out0;
assign v$Z_12567_out0 = v$G3_12676_out0;
assign v$Z_12568_out0 = v$G3_12677_out0;
assign v$Z_12569_out0 = v$G3_12678_out0;
assign v$Z_12570_out0 = v$G3_12679_out0;
assign v$SEL1_14363_out0 = v$SUM_9363_out0[23:1];
assign v$SEL1_14364_out0 = v$SUM_9366_out0[23:1];
assign v$SUM_15169_out0 = v$A1_15217_out0;
assign v$G4_17529_out0 = v$G7_18137_out0 && v$G5_5837_out0;
assign v$G4_17530_out0 = v$G7_18138_out0 && v$G5_5838_out0;
assign v$G4_17531_out0 = v$G7_18139_out0 && v$G5_5839_out0;
assign v$G4_17532_out0 = v$G7_18140_out0 && v$G5_5840_out0;
assign v$G4_17533_out0 = v$G7_18141_out0 && v$G5_5841_out0;
assign v$G4_17534_out0 = v$G7_18142_out0 && v$G5_5842_out0;
assign v$G4_17535_out0 = v$G7_18143_out0 && v$G5_5843_out0;
assign v$G4_17536_out0 = v$G7_18144_out0 && v$G5_5844_out0;
assign v$G4_17537_out0 = v$G7_18145_out0 && v$G5_5845_out0;
assign v$G4_17538_out0 = v$G7_18146_out0 && v$G5_5846_out0;
assign v$G4_17539_out0 = v$G7_18147_out0 && v$G5_5847_out0;
assign v$G4_17540_out0 = v$G7_18148_out0 && v$G5_5848_out0;
assign v$Z2_182_out0 = v$Z_12563_out0;
assign v$Z2_183_out0 = v$Z_12569_out0;
assign v$_1510_out0 = { v$SEL1_14363_out0,v$C4_3754_out0 };
assign v$_1511_out0 = { v$SEL1_14364_out0,v$C4_3755_out0 };
assign v$SUM_3469_out0 = v$SUM_15169_out0;
assign v$MUX18_4858_out0 = v$EQ18_12806_out0 ? v$SEL18_11379_out0 : v$MUX19_6374_out0;
assign v$MUX18_4859_out0 = v$EQ18_12807_out0 ? v$SEL18_11380_out0 : v$MUX19_6375_out0;
assign v$XOR1_5399_out0 = v$SUM_1905_out0 ^ v$C9_15264_out0;
assign v$XOR1_5400_out0 = v$SUM_1906_out0 ^ v$C9_15265_out0;
assign v$Z1_5767_out0 = v$Z_12564_out0;
assign v$Z1_5768_out0 = v$Z_12570_out0;
assign v$_6272_out0 = { v$G4_17529_out0,v$G9_17594_out0 };
assign v$_6273_out0 = { v$G4_17530_out0,v$G9_17595_out0 };
assign v$_6274_out0 = { v$G4_17531_out0,v$G9_17596_out0 };
assign v$_6275_out0 = { v$G4_17532_out0,v$G9_17597_out0 };
assign v$_6276_out0 = { v$G4_17533_out0,v$G9_17598_out0 };
assign v$_6277_out0 = { v$G4_17534_out0,v$G9_17599_out0 };
assign v$_6278_out0 = { v$G4_17535_out0,v$G9_17600_out0 };
assign v$_6279_out0 = { v$G4_17536_out0,v$G9_17601_out0 };
assign v$_6280_out0 = { v$G4_17537_out0,v$G9_17602_out0 };
assign v$_6281_out0 = { v$G4_17538_out0,v$G9_17603_out0 };
assign v$_6282_out0 = { v$G4_17539_out0,v$G9_17604_out0 };
assign v$_6283_out0 = { v$G4_17540_out0,v$G9_17605_out0 };
assign v$Z2_6321_out0 = v$Z_12561_out0;
assign v$Z2_6323_out0 = v$Z_12567_out0;
assign v$Z4_7919_out0 = v$Z_12562_out0;
assign v$Z4_7920_out0 = v$Z_12568_out0;
assign v$COUT_10731_out0 = v$COUT_8114_out0;
assign v$Z1_16995_out0 = v$Z_12560_out0;
assign v$Z1_16997_out0 = v$Z_12566_out0;
assign v$Z3_17777_out0 = v$Z_12559_out0;
assign v$Z3_17778_out0 = v$Z_12565_out0;
assign v$MUX7_3280_out0 = v$OVERFLOW_14976_out0 ? v$_1510_out0 : v$SUM_1905_out0;
assign v$MUX7_3281_out0 = v$OVERFLOW_14977_out0 ? v$_1511_out0 : v$SUM_1906_out0;
assign v$CIN_3891_out0 = v$COUT_10731_out0;
assign v$SEL14_4815_out0 = v$SUM_3469_out0[0:0];
assign v$G4_6053_out0 = ! v$Z4_7919_out0;
assign v$G4_6054_out0 = ! v$Z4_7920_out0;
assign v$G6_6170_out0 = ! v$Z2_6321_out0;
assign v$G6_6172_out0 = ! v$Z2_6323_out0;
assign v$Y_6489_out0 = v$_6272_out0;
assign v$Y_6490_out0 = v$_6273_out0;
assign v$Y_6491_out0 = v$_6274_out0;
assign v$Y_6492_out0 = v$_6275_out0;
assign v$Y_6493_out0 = v$_6276_out0;
assign v$Y_6494_out0 = v$_6277_out0;
assign v$Y_6495_out0 = v$_6278_out0;
assign v$Y_6496_out0 = v$_6279_out0;
assign v$Y_6497_out0 = v$_6280_out0;
assign v$Y_6498_out0 = v$_6281_out0;
assign v$Y_6499_out0 = v$_6282_out0;
assign v$Y_6500_out0 = v$_6283_out0;
assign v$A1_13595_out0 = v$XOR1_5399_out0;
assign v$A1_13598_out0 = v$XOR1_5400_out0;
assign v$OP1_14190_out0 = v$SUM_3469_out0;
assign v$G1_14594_out0 = v$Z1_5767_out0 && v$Z2_182_out0;
assign v$G1_14595_out0 = v$Z1_5768_out0 && v$Z2_183_out0;
assign v$G9_15199_out0 = v$Z1_16995_out0 && v$Z2_6321_out0;
assign v$G9_15201_out0 = v$Z1_16997_out0 && v$Z2_6323_out0;
assign v$MUX17_16536_out0 = v$EQ17_5879_out0 ? v$SEL17_16069_out0 : v$MUX18_4858_out0;
assign v$MUX17_16537_out0 = v$EQ17_5880_out0 ? v$SEL17_16070_out0 : v$MUX18_4859_out0;
assign v$G5_17507_out0 = ! v$Z3_17777_out0;
assign v$G5_17508_out0 = ! v$Z3_17778_out0;
assign v$OP1_3384_out0 = v$OP1_14190_out0;
assign v$_3977_out0 = { v$Y_6492_out0,v$C3_3302_out0 };
assign v$_3978_out0 = { v$Y_6498_out0,v$C3_3303_out0 };
assign v$_5090_out0 = { v$Y_6491_out0,v$C5_16909_out0 };
assign v$_5092_out0 = { v$Y_6497_out0,v$C5_16911_out0 };
assign v$_5469_out0 = { v$Y_6494_out0,v$C1_17669_out0 };
assign v$_5470_out0 = { v$Y_6500_out0,v$C1_17670_out0 };
assign v$_7539_out0 = v$A1_13595_out0[11:0];
assign v$_7539_out1 = v$A1_13595_out0[23:12];
assign v$_7542_out0 = v$A1_13598_out0[11:0];
assign v$_7542_out1 = v$A1_13598_out0[23:12];
assign v$_8151_out0 = { v$Y_6493_out0,v$C2_7627_out0 };
assign v$_8152_out0 = { v$Y_6499_out0,v$C2_7628_out0 };
assign v$_8781_out0 = { v$Y_6490_out0,v$C6_6535_out0 };
assign v$_8783_out0 = { v$Y_6496_out0,v$C6_6537_out0 };
assign v$_8896_out0 = { v$Y_6489_out0,v$C4_16509_out0 };
assign v$_8897_out0 = { v$Y_6495_out0,v$C4_16510_out0 };
assign v$G7_9851_out0 = v$G9_15199_out0 && v$Z3_17777_out0;
assign v$G7_9852_out0 = v$G9_15201_out0 && v$Z3_17778_out0;
assign v$Z_10332_out0 = v$G1_14594_out0;
assign v$Z_10333_out0 = v$G1_14595_out0;
assign v$SEL3_14249_out0 = v$MUX7_3280_out0[22:0];
assign v$SEL3_14250_out0 = v$MUX7_3281_out0[22:0];
assign v$SUM$10_14308_out0 = v$SEL14_4815_out0;
assign v$MUX16_16762_out0 = v$EQ16_8286_out0 ? v$SEL16_16894_out0 : v$MUX17_16536_out0;
assign v$MUX16_16763_out0 = v$EQ16_8287_out0 ? v$SEL16_16895_out0 : v$MUX17_16537_out0;
assign v$CIN_16817_out0 = v$CIN_3891_out0;
assign v$MUX5_4054_out0 = v$G6_6170_out0 ? v$_5090_out0 : v$_8781_out0;
assign v$MUX5_4056_out0 = v$G6_6172_out0 ? v$_5092_out0 : v$_8783_out0;
assign v$LOWER$PART_6314_out0 = v$MUX16_16762_out0;
assign v$LOWER$PART_6315_out0 = v$MUX16_16763_out0;
assign v$MUX1_14696_out0 = v$Z1_5767_out0 ? v$_8151_out0 : v$_5469_out0;
assign v$MUX1_14697_out0 = v$Z1_5768_out0 ? v$_8152_out0 : v$_5470_out0;
assign v$_16111_out0 = v$_7539_out0[5:0];
assign v$_16111_out1 = v$_7539_out0[11:6];
assign v$_16114_out0 = v$_7542_out0[5:0];
assign v$_16114_out1 = v$_7542_out0[11:6];
assign v$G1_16141_out0 = v$G7_9851_out0 && v$Z4_7919_out0;
assign v$G1_16142_out0 = v$G7_9852_out0 && v$Z4_7920_out0;
assign v$Z1_16994_out0 = v$Z_10332_out0;
assign v$Z1_16996_out0 = v$Z_10333_out0;
assign v$_17028_out0 = v$_7539_out1[5:0];
assign v$_17028_out1 = v$_7539_out1[11:6];
assign v$_17031_out0 = v$_7542_out1[5:0];
assign v$_17031_out1 = v$_7542_out1[11:6];
assign v$SEL8_17656_out0 = v$OP1_3384_out0[23:1];
assign v$MUX15_1317_out0 = v$EQ15_15965_out0 ? v$SEL15_4886_out0 : v$LOWER$PART_6314_out0;
assign v$MUX15_1318_out0 = v$EQ15_15966_out0 ? v$SEL15_4887_out0 : v$LOWER$PART_6315_out0;
assign v$_1863_out0 = v$_17028_out1[2:0];
assign v$_1863_out1 = v$_17028_out1[5:3];
assign v$_1866_out0 = v$_17031_out1[2:0];
assign v$_1866_out1 = v$_17031_out1[5:3];
assign v$Z_2552_out0 = v$G1_16141_out0;
assign v$Z_2554_out0 = v$G1_16142_out0;
assign v$MUX4_2871_out0 = v$G5_17507_out0 ? v$_8896_out0 : v$MUX5_4054_out0;
assign v$MUX4_2872_out0 = v$G5_17508_out0 ? v$_8897_out0 : v$MUX5_4056_out0;
assign v$Y_7759_out0 = v$MUX1_14696_out0;
assign v$Y_7760_out0 = v$MUX1_14697_out0;
assign v$_10048_out0 = v$_17028_out0[2:0];
assign v$_10048_out1 = v$_17028_out0[5:3];
assign v$_10051_out0 = v$_17031_out0[2:0];
assign v$_10051_out1 = v$_17031_out0[5:3];
assign v$_13770_out0 = v$_16111_out0[2:0];
assign v$_13770_out1 = v$_16111_out0[5:3];
assign v$_13773_out0 = v$_16114_out0[2:0];
assign v$_13773_out1 = v$_16114_out0[5:3];
assign v$_17998_out0 = { v$SEL8_17656_out0,v$CIN_16817_out0 };
assign v$_18420_out0 = v$_16111_out1[2:0];
assign v$_18420_out1 = v$_16111_out1[5:3];
assign v$_18423_out0 = v$_16114_out1[2:0];
assign v$_18423_out1 = v$_16114_out1[5:3];
assign v$_1302_out0 = v$_18420_out0[0:0];
assign v$_1302_out1 = v$_18420_out0[2:2];
assign v$_1305_out0 = v$_18423_out0[0:0];
assign v$_1305_out1 = v$_18423_out0[2:2];
assign v$_1353_out0 = v$_13770_out1[0:0];
assign v$_1353_out1 = v$_13770_out1[2:2];
assign v$_1356_out0 = v$_13773_out1[0:0];
assign v$_1356_out1 = v$_13773_out1[2:2];
assign v$_1854_out0 = v$_1863_out1[0:0];
assign v$_1854_out1 = v$_1863_out1[2:2];
assign v$_1857_out0 = v$_1866_out1[0:0];
assign v$_1857_out1 = v$_1866_out1[2:2];
assign v$MUX14_4919_out0 = v$EQ14_5401_out0 ? v$SEL14_16347_out0 : v$MUX15_1317_out0;
assign v$MUX14_4920_out0 = v$EQ14_5402_out0 ? v$SEL14_16348_out0 : v$MUX15_1318_out0;
assign v$Z2_6320_out0 = v$Z_2552_out0;
assign v$Z2_6322_out0 = v$Z_2554_out0;
assign v$_7067_out0 = v$_13770_out0[0:0];
assign v$_7067_out1 = v$_13770_out0[2:2];
assign v$_7070_out0 = v$_13773_out0[0:0];
assign v$_7070_out1 = v$_13773_out0[2:2];
assign v$_8780_out0 = { v$Y_7759_out0,v$C6_6534_out0 };
assign v$_8782_out0 = { v$Y_7760_out0,v$C6_6536_out0 };
assign v$_10446_out0 = v$_10048_out0[0:0];
assign v$_10446_out1 = v$_10048_out0[2:2];
assign v$_10449_out0 = v$_10051_out0[0:0];
assign v$_10449_out1 = v$_10051_out0[2:2];
assign v$_10910_out0 = v$_18420_out1[0:0];
assign v$_10910_out1 = v$_18420_out1[2:2];
assign v$_10913_out0 = v$_18423_out1[0:0];
assign v$_10913_out1 = v$_18423_out1[2:2];
assign v$_11099_out0 = v$_1863_out0[0:0];
assign v$_11099_out1 = v$_1863_out0[2:2];
assign v$_11102_out0 = v$_1866_out0[0:0];
assign v$_11102_out1 = v$_1866_out0[2:2];
assign {v$A1_15219_out1,v$A1_15219_out0 } = v$_17998_out0 + v$MUX1_8343_out0 + v$C6_11355_out0;
assign v$_16130_out0 = v$_10048_out1[0:0];
assign v$_16130_out1 = v$_10048_out1[2:2];
assign v$_16133_out0 = v$_10051_out1[0:0];
assign v$_16133_out1 = v$_10051_out1[2:2];
assign v$MUX3_17470_out0 = v$G4_6053_out0 ? v$_3977_out0 : v$MUX4_2871_out0;
assign v$MUX3_17471_out0 = v$G4_6054_out0 ? v$_3978_out0 : v$MUX4_2872_out0;
assign v$A6_308_out0 = v$_1302_out0;
assign v$A6_311_out0 = v$_1305_out0;
assign v$A21_2598_out0 = v$_1854_out0;
assign v$A21_2601_out0 = v$_1857_out0;
assign v$A12_3138_out0 = v$_10446_out0;
assign v$A12_3141_out0 = v$_10449_out0;
assign v$A9_3435_out0 = v$_10910_out0;
assign v$A9_3438_out0 = v$_10913_out0;
assign v$A0_4308_out0 = v$_7067_out0;
assign v$A0_4311_out0 = v$_7070_out0;
assign v$_5948_out0 = v$_16130_out1[0:0];
assign v$_5948_out1 = v$_16130_out1[1:1];
assign v$_5951_out0 = v$_16133_out1[0:0];
assign v$_5951_out1 = v$_16133_out1[1:1];
assign v$G6_6169_out0 = ! v$Z2_6320_out0;
assign v$G6_6171_out0 = ! v$Z2_6322_out0;
assign v$_7358_out0 = v$_1353_out1[0:0];
assign v$_7358_out1 = v$_1353_out1[1:1];
assign v$_7361_out0 = v$_1356_out1[0:0];
assign v$_7361_out1 = v$_1356_out1[1:1];
assign v$COUT_8116_out0 = v$A1_15219_out1;
assign v$OUT_8952_out0 = v$MUX3_17470_out0;
assign v$OUT_8954_out0 = v$MUX3_17471_out0;
assign v$_10284_out0 = v$_1854_out1[0:0];
assign v$_10284_out1 = v$_1854_out1[1:1];
assign v$_10287_out0 = v$_1857_out1[0:0];
assign v$_10287_out1 = v$_1857_out1[1:1];
assign v$_11618_out0 = v$_7067_out1[0:0];
assign v$_11618_out1 = v$_7067_out1[1:1];
assign v$_11621_out0 = v$_7070_out1[0:0];
assign v$_11621_out1 = v$_7070_out1[1:1];
assign v$MUX13_13682_out0 = v$EQ13_9515_out0 ? v$SEL13_6924_out0 : v$MUX14_4919_out0;
assign v$MUX13_13683_out0 = v$EQ13_9516_out0 ? v$SEL13_6925_out0 : v$MUX14_4920_out0;
assign v$A3_14607_out0 = v$_1353_out0;
assign v$A3_14610_out0 = v$_1356_out0;
assign v$SUM_15171_out0 = v$A1_15219_out0;
assign v$G9_15198_out0 = v$Z1_16994_out0 && v$Z2_6320_out0;
assign v$G9_15200_out0 = v$Z1_16996_out0 && v$Z2_6322_out0;
assign v$_15741_out0 = v$_1302_out1[0:0];
assign v$_15741_out1 = v$_1302_out1[1:1];
assign v$_15744_out0 = v$_1305_out1[0:0];
assign v$_15744_out1 = v$_1305_out1[1:1];
assign v$_16182_out0 = v$_10446_out1[0:0];
assign v$_16182_out1 = v$_10446_out1[1:1];
assign v$_16185_out0 = v$_10449_out1[0:0];
assign v$_16185_out1 = v$_10449_out1[1:1];
assign v$_16704_out0 = v$_11099_out1[0:0];
assign v$_16704_out1 = v$_11099_out1[1:1];
assign v$_16707_out0 = v$_11102_out1[0:0];
assign v$_16707_out1 = v$_11102_out1[1:1];
assign v$A15_17318_out0 = v$_16130_out0;
assign v$A15_17321_out0 = v$_16133_out0;
assign v$A18_17695_out0 = v$_11099_out0;
assign v$A18_17698_out0 = v$_11102_out0;
assign v$_17755_out0 = v$_10910_out1[0:0];
assign v$_17755_out1 = v$_10910_out1[1:1];
assign v$_17758_out0 = v$_10913_out1[0:0];
assign v$_17758_out1 = v$_10913_out1[1:1];
assign v$A14_676_out0 = v$_16182_out1;
assign v$A14_679_out0 = v$_16185_out1;
assign v$A19_1213_out0 = v$_16704_out0;
assign v$A19_1216_out0 = v$_16707_out0;
assign v$A10_1548_out0 = v$_17755_out0;
assign v$A10_1551_out0 = v$_17758_out0;
assign v$A1_1710_out0 = v$_11618_out0;
assign v$A1_1713_out0 = v$_11621_out0;
assign v$Z_2551_out0 = v$G9_15198_out0;
assign v$Z_2553_out0 = v$G9_15200_out0;
assign v$SUM_3471_out0 = v$SUM_15171_out0;
assign v$A22_4424_out0 = v$_10284_out0;
assign v$A22_4427_out0 = v$_10287_out0;
assign v$A20_4436_out0 = v$_16704_out1;
assign v$A20_4439_out0 = v$_16707_out1;
assign v$A23_5063_out0 = v$_10284_out1;
assign v$A23_5066_out0 = v$_10287_out1;
assign v$_5089_out0 = { v$OUT_8952_out0,v$C5_16908_out0 };
assign v$_5091_out0 = { v$OUT_8954_out0,v$C5_16910_out0 };
assign v$A5_6665_out0 = v$_7358_out1;
assign v$A5_6668_out0 = v$_7361_out1;
assign v$A_7101_out0 = v$A6_308_out0;
assign v$A_7102_out0 = v$A3_14607_out0;
assign v$A_7103_out0 = v$A21_2598_out0;
assign v$A_7104_out0 = v$A9_3435_out0;
assign v$A_7105_out0 = v$A15_17318_out0;
assign v$A_7109_out0 = v$A12_3138_out0;
assign v$A_7113_out0 = v$A0_4308_out0;
assign v$A_7118_out0 = v$A18_17695_out0;
assign v$A_7173_out0 = v$A6_311_out0;
assign v$A_7174_out0 = v$A3_14610_out0;
assign v$A_7175_out0 = v$A21_2601_out0;
assign v$A_7176_out0 = v$A9_3438_out0;
assign v$A_7177_out0 = v$A15_17321_out0;
assign v$A_7181_out0 = v$A12_3141_out0;
assign v$A_7185_out0 = v$A0_4311_out0;
assign v$A_7190_out0 = v$A18_17698_out0;
assign v$A11_9962_out0 = v$_17755_out1;
assign v$A11_9965_out0 = v$_17758_out1;
assign v$COUT_10733_out0 = v$COUT_8116_out0;
assign {v$A1A_11660_out1,v$A1A_11660_out0 } = v$A0_4308_out0 + v$B0_3200_out0 + v$C1_4464_out0;
assign {v$A1A_11663_out1,v$A1A_11663_out0 } = v$A0_4311_out0 + v$B0_3203_out0 + v$C1_4467_out0;
assign v$A16_13614_out0 = v$_5948_out0;
assign v$A16_13617_out0 = v$_5951_out0;
assign v$A13_13862_out0 = v$_16182_out0;
assign v$A13_13865_out0 = v$_16185_out0;
assign v$A7_15307_out0 = v$_15741_out0;
assign v$A7_15310_out0 = v$_15744_out0;
assign v$A17_16722_out0 = v$_5948_out1;
assign v$A17_16725_out0 = v$_5951_out1;
assign v$A4_17498_out0 = v$_7358_out0;
assign v$A4_17501_out0 = v$_7361_out0;
assign v$MUX12_17813_out0 = v$EQ12_13838_out0 ? v$SEL12_13844_out0 : v$MUX13_13682_out0;
assign v$MUX12_17814_out0 = v$EQ12_13839_out0 ? v$SEL12_13845_out0 : v$MUX13_13683_out0;
assign v$A8_18090_out0 = v$_15741_out1;
assign v$A8_18093_out0 = v$_15744_out1;
assign v$A2_18266_out0 = v$_11618_out1;
assign v$A2_18269_out0 = v$_11621_out1;
assign v$SUM_892_out0 = v$SUM_3471_out0;
assign v$CIN_3886_out0 = v$COUT_10733_out0;
assign v$MUX5_4053_out0 = v$G6_6169_out0 ? v$_5089_out0 : v$_8780_out0;
assign v$MUX5_4055_out0 = v$G6_6171_out0 ? v$_5091_out0 : v$_8782_out0;
assign v$COUT_5015_out0 = v$COUT_10733_out0;
assign v$G2_5261_out0 = ((v$A_7101_out0 && !v$B_2696_out0) || (!v$A_7101_out0) && v$B_2696_out0);
assign v$G2_5262_out0 = ((v$A_7102_out0 && !v$B_2697_out0) || (!v$A_7102_out0) && v$B_2697_out0);
assign v$G2_5263_out0 = ((v$A_7103_out0 && !v$B_2698_out0) || (!v$A_7103_out0) && v$B_2698_out0);
assign v$G2_5264_out0 = ((v$A_7104_out0 && !v$B_2699_out0) || (!v$A_7104_out0) && v$B_2699_out0);
assign v$G2_5265_out0 = ((v$A_7105_out0 && !v$B_2700_out0) || (!v$A_7105_out0) && v$B_2700_out0);
assign v$G2_5269_out0 = ((v$A_7109_out0 && !v$B_2704_out0) || (!v$A_7109_out0) && v$B_2704_out0);
assign v$G2_5273_out0 = ((v$A_7113_out0 && !v$B_2708_out0) || (!v$A_7113_out0) && v$B_2708_out0);
assign v$G2_5278_out0 = ((v$A_7118_out0 && !v$B_2713_out0) || (!v$A_7118_out0) && v$B_2713_out0);
assign v$G2_5333_out0 = ((v$A_7173_out0 && !v$B_2768_out0) || (!v$A_7173_out0) && v$B_2768_out0);
assign v$G2_5334_out0 = ((v$A_7174_out0 && !v$B_2769_out0) || (!v$A_7174_out0) && v$B_2769_out0);
assign v$G2_5335_out0 = ((v$A_7175_out0 && !v$B_2770_out0) || (!v$A_7175_out0) && v$B_2770_out0);
assign v$G2_5336_out0 = ((v$A_7176_out0 && !v$B_2771_out0) || (!v$A_7176_out0) && v$B_2771_out0);
assign v$G2_5337_out0 = ((v$A_7177_out0 && !v$B_2772_out0) || (!v$A_7177_out0) && v$B_2772_out0);
assign v$G2_5341_out0 = ((v$A_7181_out0 && !v$B_2776_out0) || (!v$A_7181_out0) && v$B_2776_out0);
assign v$G2_5345_out0 = ((v$A_7185_out0 && !v$B_2780_out0) || (!v$A_7185_out0) && v$B_2780_out0);
assign v$G2_5350_out0 = ((v$A_7190_out0 && !v$B_2785_out0) || (!v$A_7190_out0) && v$B_2785_out0);
assign v$A_7106_out0 = v$A7_15307_out0;
assign v$A_7107_out0 = v$A1_1710_out0;
assign v$A_7108_out0 = v$A14_676_out0;
assign v$A_7110_out0 = v$A8_18090_out0;
assign v$A_7111_out0 = v$A17_16722_out0;
assign v$A_7112_out0 = v$A23_5063_out0;
assign v$A_7114_out0 = v$A13_13862_out0;
assign v$A_7115_out0 = v$A4_17498_out0;
assign v$A_7116_out0 = v$A19_1213_out0;
assign v$A_7117_out0 = v$A22_4424_out0;
assign v$A_7119_out0 = v$A10_1548_out0;
assign v$A_7120_out0 = v$A20_4436_out0;
assign v$A_7121_out0 = v$A2_18266_out0;
assign v$A_7122_out0 = v$A11_9962_out0;
assign v$A_7123_out0 = v$A5_6665_out0;
assign v$A_7124_out0 = v$A16_13614_out0;
assign v$A_7178_out0 = v$A7_15310_out0;
assign v$A_7179_out0 = v$A1_1713_out0;
assign v$A_7180_out0 = v$A14_679_out0;
assign v$A_7182_out0 = v$A8_18093_out0;
assign v$A_7183_out0 = v$A17_16725_out0;
assign v$A_7184_out0 = v$A23_5066_out0;
assign v$A_7186_out0 = v$A13_13865_out0;
assign v$A_7187_out0 = v$A4_17501_out0;
assign v$A_7188_out0 = v$A19_1216_out0;
assign v$A_7189_out0 = v$A22_4427_out0;
assign v$A_7191_out0 = v$A10_1551_out0;
assign v$A_7192_out0 = v$A20_4439_out0;
assign v$A_7193_out0 = v$A2_18269_out0;
assign v$A_7194_out0 = v$A11_9965_out0;
assign v$A_7195_out0 = v$A5_6668_out0;
assign v$A_7196_out0 = v$A16_13617_out0;
assign v$SEL15_9438_out0 = v$SUM_3471_out0[0:0];
assign v$G1_12335_out0 = v$A_7101_out0 && v$B_2696_out0;
assign v$G1_12336_out0 = v$A_7102_out0 && v$B_2697_out0;
assign v$G1_12337_out0 = v$A_7103_out0 && v$B_2698_out0;
assign v$G1_12338_out0 = v$A_7104_out0 && v$B_2699_out0;
assign v$G1_12339_out0 = v$A_7105_out0 && v$B_2700_out0;
assign v$G1_12343_out0 = v$A_7109_out0 && v$B_2704_out0;
assign v$G1_12347_out0 = v$A_7113_out0 && v$B_2708_out0;
assign v$G1_12352_out0 = v$A_7118_out0 && v$B_2713_out0;
assign v$G1_12407_out0 = v$A_7173_out0 && v$B_2768_out0;
assign v$G1_12408_out0 = v$A_7174_out0 && v$B_2769_out0;
assign v$G1_12409_out0 = v$A_7175_out0 && v$B_2770_out0;
assign v$G1_12410_out0 = v$A_7176_out0 && v$B_2771_out0;
assign v$G1_12411_out0 = v$A_7177_out0 && v$B_2772_out0;
assign v$G1_12415_out0 = v$A_7181_out0 && v$B_2776_out0;
assign v$G1_12419_out0 = v$A_7185_out0 && v$B_2780_out0;
assign v$G1_12424_out0 = v$A_7190_out0 && v$B_2785_out0;
assign v$OP1_14185_out0 = v$SUM_3471_out0;
assign v$Z_15808_out0 = v$Z_2551_out0;
assign v$Z_15809_out0 = v$Z_2553_out0;
assign v$MUX11_17933_out0 = v$EQ11_6143_out0 ? v$SEL11_7225_out0 : v$MUX12_17813_out0;
assign v$MUX11_17934_out0 = v$EQ11_6144_out0 ? v$SEL11_7226_out0 : v$MUX12_17814_out0;
assign v$END_18272_out0 = v$A1A_11660_out1;
assign v$END_18275_out0 = v$A1A_11663_out1;
assign v$MUX8_2945_out0 = v$EQ9_13775_out0 ? v$SEL9_10263_out0 : v$MUX11_17933_out0;
assign v$MUX8_2946_out0 = v$EQ9_13776_out0 ? v$SEL9_10264_out0 : v$MUX11_17934_out0;
assign v$OP1_3379_out0 = v$OP1_14185_out0;
assign v$G2_5266_out0 = ((v$A_7106_out0 && !v$B_2701_out0) || (!v$A_7106_out0) && v$B_2701_out0);
assign v$G2_5267_out0 = ((v$A_7107_out0 && !v$B_2702_out0) || (!v$A_7107_out0) && v$B_2702_out0);
assign v$G2_5268_out0 = ((v$A_7108_out0 && !v$B_2703_out0) || (!v$A_7108_out0) && v$B_2703_out0);
assign v$G2_5270_out0 = ((v$A_7110_out0 && !v$B_2705_out0) || (!v$A_7110_out0) && v$B_2705_out0);
assign v$G2_5271_out0 = ((v$A_7111_out0 && !v$B_2706_out0) || (!v$A_7111_out0) && v$B_2706_out0);
assign v$G2_5272_out0 = ((v$A_7112_out0 && !v$B_2707_out0) || (!v$A_7112_out0) && v$B_2707_out0);
assign v$G2_5274_out0 = ((v$A_7114_out0 && !v$B_2709_out0) || (!v$A_7114_out0) && v$B_2709_out0);
assign v$G2_5275_out0 = ((v$A_7115_out0 && !v$B_2710_out0) || (!v$A_7115_out0) && v$B_2710_out0);
assign v$G2_5276_out0 = ((v$A_7116_out0 && !v$B_2711_out0) || (!v$A_7116_out0) && v$B_2711_out0);
assign v$G2_5277_out0 = ((v$A_7117_out0 && !v$B_2712_out0) || (!v$A_7117_out0) && v$B_2712_out0);
assign v$G2_5279_out0 = ((v$A_7119_out0 && !v$B_2714_out0) || (!v$A_7119_out0) && v$B_2714_out0);
assign v$G2_5280_out0 = ((v$A_7120_out0 && !v$B_2715_out0) || (!v$A_7120_out0) && v$B_2715_out0);
assign v$G2_5281_out0 = ((v$A_7121_out0 && !v$B_2716_out0) || (!v$A_7121_out0) && v$B_2716_out0);
assign v$G2_5282_out0 = ((v$A_7122_out0 && !v$B_2717_out0) || (!v$A_7122_out0) && v$B_2717_out0);
assign v$G2_5283_out0 = ((v$A_7123_out0 && !v$B_2718_out0) || (!v$A_7123_out0) && v$B_2718_out0);
assign v$G2_5284_out0 = ((v$A_7124_out0 && !v$B_2719_out0) || (!v$A_7124_out0) && v$B_2719_out0);
assign v$G2_5338_out0 = ((v$A_7178_out0 && !v$B_2773_out0) || (!v$A_7178_out0) && v$B_2773_out0);
assign v$G2_5339_out0 = ((v$A_7179_out0 && !v$B_2774_out0) || (!v$A_7179_out0) && v$B_2774_out0);
assign v$G2_5340_out0 = ((v$A_7180_out0 && !v$B_2775_out0) || (!v$A_7180_out0) && v$B_2775_out0);
assign v$G2_5342_out0 = ((v$A_7182_out0 && !v$B_2777_out0) || (!v$A_7182_out0) && v$B_2777_out0);
assign v$G2_5343_out0 = ((v$A_7183_out0 && !v$B_2778_out0) || (!v$A_7183_out0) && v$B_2778_out0);
assign v$G2_5344_out0 = ((v$A_7184_out0 && !v$B_2779_out0) || (!v$A_7184_out0) && v$B_2779_out0);
assign v$G2_5346_out0 = ((v$A_7186_out0 && !v$B_2781_out0) || (!v$A_7186_out0) && v$B_2781_out0);
assign v$G2_5347_out0 = ((v$A_7187_out0 && !v$B_2782_out0) || (!v$A_7187_out0) && v$B_2782_out0);
assign v$G2_5348_out0 = ((v$A_7188_out0 && !v$B_2783_out0) || (!v$A_7188_out0) && v$B_2783_out0);
assign v$G2_5349_out0 = ((v$A_7189_out0 && !v$B_2784_out0) || (!v$A_7189_out0) && v$B_2784_out0);
assign v$G2_5351_out0 = ((v$A_7191_out0 && !v$B_2786_out0) || (!v$A_7191_out0) && v$B_2786_out0);
assign v$G2_5352_out0 = ((v$A_7192_out0 && !v$B_2787_out0) || (!v$A_7192_out0) && v$B_2787_out0);
assign v$G2_5353_out0 = ((v$A_7193_out0 && !v$B_2788_out0) || (!v$A_7193_out0) && v$B_2788_out0);
assign v$G2_5354_out0 = ((v$A_7194_out0 && !v$B_2789_out0) || (!v$A_7194_out0) && v$B_2789_out0);
assign v$G2_5355_out0 = ((v$A_7195_out0 && !v$B_2790_out0) || (!v$A_7195_out0) && v$B_2790_out0);
assign v$G2_5356_out0 = ((v$A_7196_out0 && !v$B_2791_out0) || (!v$A_7196_out0) && v$B_2791_out0);
assign v$OUT_8951_out0 = v$MUX5_4053_out0;
assign v$OUT_8953_out0 = v$MUX5_4055_out0;
assign v$G_10055_out0 = v$G1_12335_out0;
assign v$G_10056_out0 = v$G1_12336_out0;
assign v$G_10057_out0 = v$G1_12337_out0;
assign v$G_10058_out0 = v$G1_12338_out0;
assign v$G_10059_out0 = v$G1_12339_out0;
assign v$G_10063_out0 = v$G1_12343_out0;
assign v$G_10067_out0 = v$G1_12347_out0;
assign v$G_10072_out0 = v$G1_12352_out0;
assign v$G_10127_out0 = v$G1_12407_out0;
assign v$G_10128_out0 = v$G1_12408_out0;
assign v$G_10129_out0 = v$G1_12409_out0;
assign v$G_10130_out0 = v$G1_12410_out0;
assign v$G_10131_out0 = v$G1_12411_out0;
assign v$G_10135_out0 = v$G1_12415_out0;
assign v$G_10139_out0 = v$G1_12419_out0;
assign v$G_10144_out0 = v$G1_12424_out0;
assign v$_10453_out0 = { v$SUM_892_out0,v$COUT_5015_out0 };
assign v$G1_12340_out0 = v$A_7106_out0 && v$B_2701_out0;
assign v$G1_12341_out0 = v$A_7107_out0 && v$B_2702_out0;
assign v$G1_12342_out0 = v$A_7108_out0 && v$B_2703_out0;
assign v$G1_12344_out0 = v$A_7110_out0 && v$B_2705_out0;
assign v$G1_12345_out0 = v$A_7111_out0 && v$B_2706_out0;
assign v$G1_12346_out0 = v$A_7112_out0 && v$B_2707_out0;
assign v$G1_12348_out0 = v$A_7114_out0 && v$B_2709_out0;
assign v$G1_12349_out0 = v$A_7115_out0 && v$B_2710_out0;
assign v$G1_12350_out0 = v$A_7116_out0 && v$B_2711_out0;
assign v$G1_12351_out0 = v$A_7117_out0 && v$B_2712_out0;
assign v$G1_12353_out0 = v$A_7119_out0 && v$B_2714_out0;
assign v$G1_12354_out0 = v$A_7120_out0 && v$B_2715_out0;
assign v$G1_12355_out0 = v$A_7121_out0 && v$B_2716_out0;
assign v$G1_12356_out0 = v$A_7122_out0 && v$B_2717_out0;
assign v$G1_12357_out0 = v$A_7123_out0 && v$B_2718_out0;
assign v$G1_12358_out0 = v$A_7124_out0 && v$B_2719_out0;
assign v$G1_12412_out0 = v$A_7178_out0 && v$B_2773_out0;
assign v$G1_12413_out0 = v$A_7179_out0 && v$B_2774_out0;
assign v$G1_12414_out0 = v$A_7180_out0 && v$B_2775_out0;
assign v$G1_12416_out0 = v$A_7182_out0 && v$B_2777_out0;
assign v$G1_12417_out0 = v$A_7183_out0 && v$B_2778_out0;
assign v$G1_12418_out0 = v$A_7184_out0 && v$B_2779_out0;
assign v$G1_12420_out0 = v$A_7186_out0 && v$B_2781_out0;
assign v$G1_12421_out0 = v$A_7187_out0 && v$B_2782_out0;
assign v$G1_12422_out0 = v$A_7188_out0 && v$B_2783_out0;
assign v$G1_12423_out0 = v$A_7189_out0 && v$B_2784_out0;
assign v$G1_12425_out0 = v$A_7191_out0 && v$B_2786_out0;
assign v$G1_12426_out0 = v$A_7192_out0 && v$B_2787_out0;
assign v$G1_12427_out0 = v$A_7193_out0 && v$B_2788_out0;
assign v$G1_12428_out0 = v$A_7194_out0 && v$B_2789_out0;
assign v$G1_12429_out0 = v$A_7195_out0 && v$B_2790_out0;
assign v$G1_12430_out0 = v$A_7196_out0 && v$B_2791_out0;
assign v$P_13868_out0 = v$G2_5261_out0;
assign v$P_13869_out0 = v$G2_5262_out0;
assign v$P_13870_out0 = v$G2_5263_out0;
assign v$P_13871_out0 = v$G2_5264_out0;
assign v$P_13872_out0 = v$G2_5265_out0;
assign v$P_13876_out0 = v$G2_5269_out0;
assign v$P_13880_out0 = v$G2_5273_out0;
assign v$P_13885_out0 = v$G2_5278_out0;
assign v$P_13940_out0 = v$G2_5333_out0;
assign v$P_13941_out0 = v$G2_5334_out0;
assign v$P_13942_out0 = v$G2_5335_out0;
assign v$P_13943_out0 = v$G2_5336_out0;
assign v$P_13944_out0 = v$G2_5337_out0;
assign v$P_13948_out0 = v$G2_5341_out0;
assign v$P_13952_out0 = v$G2_5345_out0;
assign v$P_13957_out0 = v$G2_5350_out0;
assign v$CIN_16812_out0 = v$CIN_3886_out0;
assign v$SUM$11_17033_out0 = v$SEL15_9438_out0;
assign v$P12_235_out0 = v$P_13876_out0;
assign v$P12_238_out0 = v$P_13948_out0;
assign v$P21_4769_out0 = v$P_13870_out0;
assign v$P21_4772_out0 = v$P_13942_out0;
assign v$P0_4810_out0 = v$P_13880_out0;
assign v$P0_4813_out0 = v$P_13952_out0;
assign v$_4910_out0 = { v$SUM$11_17033_out0,v$_10453_out0 };
assign v$P15_6904_out0 = v$P_13872_out0;
assign v$P15_6907_out0 = v$P_13944_out0;
assign v$G12_7042_out0 = v$G_10063_out0;
assign v$G12_7045_out0 = v$G_10135_out0;
assign v$P6_8104_out0 = v$P_13868_out0;
assign v$P6_8107_out0 = v$P_13940_out0;
assign v$G9_8925_out0 = v$G_10058_out0;
assign v$G9_8928_out0 = v$G_10130_out0;
assign v$AMOUNT$OF$SHIFT_9459_out0 = v$OUT_8951_out0;
assign v$AMOUNT$OF$SHIFT_9460_out0 = v$OUT_8953_out0;
assign v$G_10060_out0 = v$G1_12340_out0;
assign v$G_10061_out0 = v$G1_12341_out0;
assign v$G_10062_out0 = v$G1_12342_out0;
assign v$G_10064_out0 = v$G1_12344_out0;
assign v$G_10065_out0 = v$G1_12345_out0;
assign v$G_10066_out0 = v$G1_12346_out0;
assign v$G_10068_out0 = v$G1_12348_out0;
assign v$G_10069_out0 = v$G1_12349_out0;
assign v$G_10070_out0 = v$G1_12350_out0;
assign v$G_10071_out0 = v$G1_12351_out0;
assign v$G_10073_out0 = v$G1_12353_out0;
assign v$G_10074_out0 = v$G1_12354_out0;
assign v$G_10075_out0 = v$G1_12355_out0;
assign v$G_10076_out0 = v$G1_12356_out0;
assign v$G_10077_out0 = v$G1_12357_out0;
assign v$G_10078_out0 = v$G1_12358_out0;
assign v$G_10132_out0 = v$G1_12412_out0;
assign v$G_10133_out0 = v$G1_12413_out0;
assign v$G_10134_out0 = v$G1_12414_out0;
assign v$G_10136_out0 = v$G1_12416_out0;
assign v$G_10137_out0 = v$G1_12417_out0;
assign v$G_10138_out0 = v$G1_12418_out0;
assign v$G_10140_out0 = v$G1_12420_out0;
assign v$G_10141_out0 = v$G1_12421_out0;
assign v$G_10142_out0 = v$G1_12422_out0;
assign v$G_10143_out0 = v$G1_12423_out0;
assign v$G_10145_out0 = v$G1_12425_out0;
assign v$G_10146_out0 = v$G1_12426_out0;
assign v$G_10147_out0 = v$G1_12427_out0;
assign v$G_10148_out0 = v$G1_12428_out0;
assign v$G_10149_out0 = v$G1_12429_out0;
assign v$G_10150_out0 = v$G1_12430_out0;
assign v$G15_11030_out0 = v$G_10059_out0;
assign v$G15_11033_out0 = v$G_10131_out0;
assign v$G3_11104_out0 = v$G_10056_out0;
assign v$G3_11107_out0 = v$G_10128_out0;
assign v$P18_11722_out0 = v$P_13885_out0;
assign v$P18_11725_out0 = v$P_13957_out0;
assign v$G18_12938_out0 = v$G_10072_out0;
assign v$G18_12941_out0 = v$G_10144_out0;
assign v$P_13873_out0 = v$G2_5266_out0;
assign v$P_13874_out0 = v$G2_5267_out0;
assign v$P_13875_out0 = v$G2_5268_out0;
assign v$P_13877_out0 = v$G2_5270_out0;
assign v$P_13878_out0 = v$G2_5271_out0;
assign v$P_13879_out0 = v$G2_5272_out0;
assign v$P_13881_out0 = v$G2_5274_out0;
assign v$P_13882_out0 = v$G2_5275_out0;
assign v$P_13883_out0 = v$G2_5276_out0;
assign v$P_13884_out0 = v$G2_5277_out0;
assign v$P_13886_out0 = v$G2_5279_out0;
assign v$P_13887_out0 = v$G2_5280_out0;
assign v$P_13888_out0 = v$G2_5281_out0;
assign v$P_13889_out0 = v$G2_5282_out0;
assign v$P_13890_out0 = v$G2_5283_out0;
assign v$P_13891_out0 = v$G2_5284_out0;
assign v$P_13945_out0 = v$G2_5338_out0;
assign v$P_13946_out0 = v$G2_5339_out0;
assign v$P_13947_out0 = v$G2_5340_out0;
assign v$P_13949_out0 = v$G2_5342_out0;
assign v$P_13950_out0 = v$G2_5343_out0;
assign v$P_13951_out0 = v$G2_5344_out0;
assign v$P_13953_out0 = v$G2_5346_out0;
assign v$P_13954_out0 = v$G2_5347_out0;
assign v$P_13955_out0 = v$G2_5348_out0;
assign v$P_13956_out0 = v$G2_5349_out0;
assign v$P_13958_out0 = v$G2_5351_out0;
assign v$P_13959_out0 = v$G2_5352_out0;
assign v$P_13960_out0 = v$G2_5353_out0;
assign v$P_13961_out0 = v$G2_5354_out0;
assign v$P_13962_out0 = v$G2_5355_out0;
assign v$P_13963_out0 = v$G2_5356_out0;
assign v$G21_14017_out0 = v$G_10057_out0;
assign v$G21_14020_out0 = v$G_10129_out0;
assign v$P3_15335_out0 = v$P_13869_out0;
assign v$P3_15338_out0 = v$P_13941_out0;
assign v$MUX10_15672_out0 = v$EQ10_5892_out0 ? v$SEL8_17683_out0 : v$MUX8_2945_out0;
assign v$MUX10_15673_out0 = v$EQ10_5893_out0 ? v$SEL8_17684_out0 : v$MUX8_2946_out0;
assign v$G0_15942_out0 = v$G_10067_out0;
assign v$G0_15945_out0 = v$G_10139_out0;
assign v$G6_16353_out0 = v$G_10055_out0;
assign v$G6_16356_out0 = v$G_10127_out0;
assign v$SEL8_17651_out0 = v$OP1_3379_out0[23:1];
assign v$P9_18445_out0 = v$P_13871_out0;
assign v$P9_18448_out0 = v$P_13943_out0;
assign v$P5_221_out0 = v$P_13890_out0;
assign v$P5_224_out0 = v$P_13962_out0;
assign v$P10_344_out0 = v$P_13886_out0;
assign v$P10_347_out0 = v$P_13958_out0;
assign v$G$CD_924_out0 = v$G6_16353_out0;
assign v$G$CD_925_out0 = v$G3_11104_out0;
assign v$G$CD_926_out0 = v$G12_7042_out0;
assign v$G$CD_927_out0 = v$G9_8925_out0;
assign v$G$CD_930_out0 = v$G18_12938_out0;
assign v$G$CD_941_out0 = v$G15_11030_out0;
assign v$G$CD_942_out0 = v$G21_14017_out0;
assign v$G$CD_1047_out0 = v$G6_16356_out0;
assign v$G$CD_1048_out0 = v$G3_11107_out0;
assign v$G$CD_1049_out0 = v$G12_7045_out0;
assign v$G$CD_1050_out0 = v$G9_8928_out0;
assign v$G$CD_1053_out0 = v$G18_12941_out0;
assign v$G$CD_1064_out0 = v$G15_11033_out0;
assign v$G$CD_1065_out0 = v$G21_14020_out0;
assign v$G7_1691_out0 = v$G_10060_out0;
assign v$G7_1694_out0 = v$G_10132_out0;
assign v$P8_1703_out0 = v$P_13877_out0;
assign v$P8_1706_out0 = v$P_13949_out0;
assign v$G10_1833_out0 = v$G_10073_out0;
assign v$G10_1836_out0 = v$G_10145_out0;
assign v$SEL4_1845_out0 = v$AMOUNT$OF$SHIFT_9459_out0[3:3];
assign v$SEL4_1846_out0 = v$AMOUNT$OF$SHIFT_9460_out0[3:3];
assign v$G19_1881_out0 = v$G_10070_out0;
assign v$G19_1884_out0 = v$G_10142_out0;
assign v$P$AB_2005_out0 = v$P0_4810_out0;
assign v$P$AB_2008_out0 = v$P18_11722_out0;
assign v$P$AB_2009_out0 = v$P21_4769_out0;
assign v$P$AB_2021_out0 = v$P12_235_out0;
assign v$P$AB_2023_out0 = v$P15_6904_out0;
assign v$P$AB_2026_out0 = v$P6_8104_out0;
assign v$P$AB_2032_out0 = v$P3_15335_out0;
assign v$P$AB_2037_out0 = v$P9_18445_out0;
assign v$P$AB_2128_out0 = v$P0_4813_out0;
assign v$P$AB_2131_out0 = v$P18_11725_out0;
assign v$P$AB_2132_out0 = v$P21_4772_out0;
assign v$P$AB_2144_out0 = v$P12_238_out0;
assign v$P$AB_2146_out0 = v$P15_6907_out0;
assign v$P$AB_2149_out0 = v$P6_8107_out0;
assign v$P$AB_2155_out0 = v$P3_15338_out0;
assign v$P$AB_2160_out0 = v$P9_18448_out0;
assign v$P2_2219_out0 = v$P_13888_out0;
assign v$P2_2222_out0 = v$P_13960_out0;
assign v$G8_2577_out0 = v$G_10064_out0;
assign v$G8_2580_out0 = v$G_10136_out0;
assign v$G13_2828_out0 = v$G_10068_out0;
assign v$G13_2831_out0 = v$G_10140_out0;
assign v$P1_2959_out0 = v$P_13874_out0;
assign v$P1_2962_out0 = v$P_13946_out0;
assign v$P13_3032_out0 = v$P_13881_out0;
assign v$P13_3035_out0 = v$P_13953_out0;
assign v$P14_3151_out0 = v$P_13875_out0;
assign v$P14_3154_out0 = v$P_13947_out0;
assign v$P22_4734_out0 = v$P_13884_out0;
assign v$P22_4737_out0 = v$P_13956_out0;
assign v$G1_5053_out0 = v$G_10061_out0;
assign v$G1_5056_out0 = v$G_10133_out0;
assign v$G4_5735_out0 = v$G_10069_out0;
assign v$G4_5738_out0 = v$G_10141_out0;
assign v$P23_6386_out0 = v$P_13879_out0;
assign v$P23_6389_out0 = v$P_13951_out0;
assign v$P16_6962_out0 = v$P_13891_out0;
assign v$P16_6965_out0 = v$P_13963_out0;
assign v$G20_8225_out0 = v$G_10074_out0;
assign v$G20_8228_out0 = v$G_10146_out0;
assign v$MUX9_8243_out0 = v$EQ8_14414_out0 ? v$SEL10_9506_out0 : v$MUX10_15672_out0;
assign v$MUX9_8244_out0 = v$EQ8_14415_out0 ? v$SEL10_9507_out0 : v$MUX10_15673_out0;
assign v$G$AB_9140_out0 = v$G0_15942_out0;
assign v$G$AB_9143_out0 = v$G18_12938_out0;
assign v$G$AB_9144_out0 = v$G21_14017_out0;
assign v$G$AB_9156_out0 = v$G12_7042_out0;
assign v$G$AB_9158_out0 = v$G15_11030_out0;
assign v$G$AB_9161_out0 = v$G6_16353_out0;
assign v$G$AB_9167_out0 = v$G3_11104_out0;
assign v$G$AB_9172_out0 = v$G9_8925_out0;
assign v$G$AB_9263_out0 = v$G0_15945_out0;
assign v$G$AB_9266_out0 = v$G18_12941_out0;
assign v$G$AB_9267_out0 = v$G21_14020_out0;
assign v$G$AB_9279_out0 = v$G12_7045_out0;
assign v$G$AB_9281_out0 = v$G15_11033_out0;
assign v$G$AB_9284_out0 = v$G6_16356_out0;
assign v$G$AB_9290_out0 = v$G3_11107_out0;
assign v$G$AB_9295_out0 = v$G9_8928_out0;
assign v$G17_9346_out0 = v$G_10065_out0;
assign v$G17_9349_out0 = v$G_10137_out0;
assign v$P11_9611_out0 = v$P_13889_out0;
assign v$P11_9614_out0 = v$P_13961_out0;
assign v$P$CD_10464_out0 = v$P6_8104_out0;
assign v$P$CD_10465_out0 = v$P3_15335_out0;
assign v$P$CD_10466_out0 = v$P12_235_out0;
assign v$P$CD_10467_out0 = v$P9_18445_out0;
assign v$P$CD_10470_out0 = v$P18_11722_out0;
assign v$P$CD_10481_out0 = v$P15_6904_out0;
assign v$P$CD_10482_out0 = v$P21_4769_out0;
assign v$P$CD_10587_out0 = v$P6_8107_out0;
assign v$P$CD_10588_out0 = v$P3_15338_out0;
assign v$P$CD_10589_out0 = v$P12_238_out0;
assign v$P$CD_10590_out0 = v$P9_18448_out0;
assign v$P$CD_10593_out0 = v$P18_11725_out0;
assign v$P$CD_10604_out0 = v$P15_6907_out0;
assign v$P$CD_10605_out0 = v$P21_4772_out0;
assign v$P20_10659_out0 = v$P_13887_out0;
assign v$P20_10662_out0 = v$P_13959_out0;
assign v$G5_10676_out0 = v$G_10077_out0;
assign v$G5_10679_out0 = v$G_10149_out0;
assign v$G11_11063_out0 = v$G_10076_out0;
assign v$G11_11066_out0 = v$G_10148_out0;
assign v$SEL5_11667_out0 = v$AMOUNT$OF$SHIFT_9459_out0[4:4];
assign v$SEL5_11668_out0 = v$AMOUNT$OF$SHIFT_9460_out0[4:4];
assign v$P17_11759_out0 = v$P_13878_out0;
assign v$P17_11762_out0 = v$P_13950_out0;
assign v$P7_11769_out0 = v$P_13873_out0;
assign v$P7_11772_out0 = v$P_13945_out0;
assign v$G22_12510_out0 = v$G_10071_out0;
assign v$G22_12513_out0 = v$G_10143_out0;
assign v$SEL1_13355_out0 = v$AMOUNT$OF$SHIFT_9459_out0[0:0];
assign v$SEL1_13356_out0 = v$AMOUNT$OF$SHIFT_9460_out0[0:0];
assign v$P4_13636_out0 = v$P_13882_out0;
assign v$P4_13639_out0 = v$P_13954_out0;
assign v$_13990_out0 = { v$SUM$10_14308_out0,v$_4910_out0 };
assign v$SEL3_14006_out0 = v$AMOUNT$OF$SHIFT_9459_out0[2:2];
assign v$SEL3_14007_out0 = v$AMOUNT$OF$SHIFT_9460_out0[2:2];
assign v$G23_14317_out0 = v$G_10066_out0;
assign v$G23_14320_out0 = v$G_10138_out0;
assign v$GATE2_15756_out0 = v$CIN_16106_out0 && v$P0_4810_out0;
assign v$GATE2_15759_out0 = v$CIN_16109_out0 && v$P0_4813_out0;
assign v$G2_15960_out0 = v$G_10075_out0;
assign v$G2_15963_out0 = v$G_10147_out0;
assign v$P19_16317_out0 = v$P_13883_out0;
assign v$P19_16320_out0 = v$P_13955_out0;
assign v$G16_16448_out0 = v$G_10078_out0;
assign v$G16_16451_out0 = v$G_10150_out0;
assign v$G14_17976_out0 = v$G_10062_out0;
assign v$G14_17979_out0 = v$G_10134_out0;
assign v$_17993_out0 = { v$SEL8_17651_out0,v$CIN_16812_out0 };
assign v$SEL2_18502_out0 = v$AMOUNT$OF$SHIFT_9459_out0[1:1];
assign v$SEL2_18503_out0 = v$AMOUNT$OF$SHIFT_9460_out0[1:1];
assign v$GATE1_659_out0 = v$GATE2_15756_out0 || v$G0_15942_out0;
assign v$GATE1_662_out0 = v$GATE2_15759_out0 || v$G0_15945_out0;
assign v$G$CD_915_out0 = v$G14_17976_out0;
assign v$G$CD_916_out0 = v$G8_2577_out0;
assign v$G$CD_918_out0 = v$G1_5053_out0;
assign v$G$CD_921_out0 = v$G19_1881_out0;
assign v$G$CD_922_out0 = v$G22_12510_out0;
assign v$G$CD_929_out0 = v$G23_14317_out0;
assign v$G$CD_931_out0 = v$G2_15960_out0;
assign v$G$CD_932_out0 = v$G5_10676_out0;
assign v$G$CD_934_out0 = v$G13_2828_out0;
assign v$G$CD_935_out0 = v$G17_9346_out0;
assign v$G$CD_936_out0 = v$G16_16448_out0;
assign v$G$CD_939_out0 = v$G7_1691_out0;
assign v$G$CD_945_out0 = v$G4_5735_out0;
assign v$G$CD_949_out0 = v$G20_8225_out0;
assign v$G$CD_950_out0 = v$G10_1833_out0;
assign v$G$CD_954_out0 = v$G11_11063_out0;
assign v$G$CD_1038_out0 = v$G14_17979_out0;
assign v$G$CD_1039_out0 = v$G8_2580_out0;
assign v$G$CD_1041_out0 = v$G1_5056_out0;
assign v$G$CD_1044_out0 = v$G19_1884_out0;
assign v$G$CD_1045_out0 = v$G22_12513_out0;
assign v$G$CD_1052_out0 = v$G23_14320_out0;
assign v$G$CD_1054_out0 = v$G2_15963_out0;
assign v$G$CD_1055_out0 = v$G5_10679_out0;
assign v$G$CD_1057_out0 = v$G13_2831_out0;
assign v$G$CD_1058_out0 = v$G17_9349_out0;
assign v$G$CD_1059_out0 = v$G16_16451_out0;
assign v$G$CD_1062_out0 = v$G7_1694_out0;
assign v$G$CD_1068_out0 = v$G4_5738_out0;
assign v$G$CD_1072_out0 = v$G20_8228_out0;
assign v$G$CD_1073_out0 = v$G10_1836_out0;
assign v$G$CD_1077_out0 = v$G11_11066_out0;
assign v$MUX7_1227_out0 = v$EQ7_4085_out0 ? v$SEL7_14332_out0 : v$MUX9_8243_out0;
assign v$MUX7_1228_out0 = v$EQ7_4086_out0 ? v$SEL7_14333_out0 : v$MUX9_8244_out0;
assign v$EN_1337_out0 = v$SEL4_1845_out0;
assign v$EN_1340_out0 = v$SEL4_1846_out0;
assign v$EN_3875_out0 = v$SEL1_13355_out0;
assign v$EN_3876_out0 = v$SEL1_13356_out0;
assign v$EN_4754_out0 = v$SEL3_14006_out0;
assign v$EN_4756_out0 = v$SEL3_14007_out0;
assign v$EN_5213_out0 = v$SEL5_11667_out0;
assign v$EN_5215_out0 = v$SEL5_11668_out0;
assign v$EN_7876_out0 = v$SEL2_18502_out0;
assign v$EN_7878_out0 = v$SEL2_18503_out0;
assign v$_10037_out0 = { v$SUM$9_197_out0,v$_13990_out0 };
assign v$P$CD_10455_out0 = v$P14_3151_out0;
assign v$P$CD_10456_out0 = v$P8_1703_out0;
assign v$P$CD_10458_out0 = v$P1_2959_out0;
assign v$P$CD_10461_out0 = v$P19_16317_out0;
assign v$P$CD_10462_out0 = v$P22_4734_out0;
assign v$P$CD_10469_out0 = v$P23_6386_out0;
assign v$P$CD_10471_out0 = v$P2_2219_out0;
assign v$P$CD_10472_out0 = v$P5_221_out0;
assign v$P$CD_10474_out0 = v$P13_3032_out0;
assign v$P$CD_10475_out0 = v$P17_11759_out0;
assign v$P$CD_10476_out0 = v$P16_6962_out0;
assign v$P$CD_10479_out0 = v$P7_11769_out0;
assign v$P$CD_10485_out0 = v$P4_13636_out0;
assign v$P$CD_10489_out0 = v$P20_10659_out0;
assign v$P$CD_10490_out0 = v$P10_344_out0;
assign v$P$CD_10494_out0 = v$P11_9611_out0;
assign v$P$CD_10578_out0 = v$P14_3154_out0;
assign v$P$CD_10579_out0 = v$P8_1706_out0;
assign v$P$CD_10581_out0 = v$P1_2962_out0;
assign v$P$CD_10584_out0 = v$P19_16320_out0;
assign v$P$CD_10585_out0 = v$P22_4737_out0;
assign v$P$CD_10592_out0 = v$P23_6389_out0;
assign v$P$CD_10594_out0 = v$P2_2222_out0;
assign v$P$CD_10595_out0 = v$P5_224_out0;
assign v$P$CD_10597_out0 = v$P13_3035_out0;
assign v$P$CD_10598_out0 = v$P17_11762_out0;
assign v$P$CD_10599_out0 = v$P16_6965_out0;
assign v$P$CD_10602_out0 = v$P7_11772_out0;
assign v$P$CD_10608_out0 = v$P4_13639_out0;
assign v$P$CD_10612_out0 = v$P20_10662_out0;
assign v$P$CD_10613_out0 = v$P10_347_out0;
assign v$P$CD_10617_out0 = v$P11_9614_out0;
assign v$G8_11399_out0 = v$CINA_8468_out0 && v$P$AB_2005_out0;
assign v$G8_11402_out0 = v$CINA_8471_out0 && v$P$AB_2008_out0;
assign v$G8_11403_out0 = v$CINA_8472_out0 && v$P$AB_2009_out0;
assign v$G8_11415_out0 = v$CINA_8484_out0 && v$P$AB_2021_out0;
assign v$G8_11417_out0 = v$CINA_8486_out0 && v$P$AB_2023_out0;
assign v$G8_11420_out0 = v$CINA_8489_out0 && v$P$AB_2026_out0;
assign v$G8_11426_out0 = v$CINA_8495_out0 && v$P$AB_2032_out0;
assign v$G8_11431_out0 = v$CINA_8500_out0 && v$P$AB_2037_out0;
assign v$G8_11522_out0 = v$CINA_8591_out0 && v$P$AB_2128_out0;
assign v$G8_11525_out0 = v$CINA_8594_out0 && v$P$AB_2131_out0;
assign v$G8_11526_out0 = v$CINA_8595_out0 && v$P$AB_2132_out0;
assign v$G8_11538_out0 = v$CINA_8607_out0 && v$P$AB_2144_out0;
assign v$G8_11540_out0 = v$CINA_8609_out0 && v$P$AB_2146_out0;
assign v$G8_11543_out0 = v$CINA_8612_out0 && v$P$AB_2149_out0;
assign v$G8_11549_out0 = v$CINA_8618_out0 && v$P$AB_2155_out0;
assign v$G8_11554_out0 = v$CINA_8623_out0 && v$P$AB_2160_out0;
assign {v$A1_15214_out1,v$A1_15214_out0 } = v$_17993_out0 + v$MUX1_8338_out0 + v$C6_11350_out0;
assign v$G5_4523_out0 = v$G$AB_9140_out0 && v$P$CD_10458_out0;
assign v$G5_4526_out0 = v$G$AB_9143_out0 && v$P$CD_10461_out0;
assign v$G5_4527_out0 = v$G$AB_9144_out0 && v$P$CD_10462_out0;
assign v$G5_4539_out0 = v$G$AB_9156_out0 && v$P$CD_10474_out0;
assign v$G5_4541_out0 = v$G$AB_9158_out0 && v$P$CD_10476_out0;
assign v$G5_4544_out0 = v$G$AB_9161_out0 && v$P$CD_10479_out0;
assign v$G5_4550_out0 = v$G$AB_9167_out0 && v$P$CD_10485_out0;
assign v$G5_4555_out0 = v$G$AB_9172_out0 && v$P$CD_10490_out0;
assign v$G5_4646_out0 = v$G$AB_9263_out0 && v$P$CD_10581_out0;
assign v$G5_4649_out0 = v$G$AB_9266_out0 && v$P$CD_10584_out0;
assign v$G5_4650_out0 = v$G$AB_9267_out0 && v$P$CD_10585_out0;
assign v$G5_4662_out0 = v$G$AB_9279_out0 && v$P$CD_10597_out0;
assign v$G5_4664_out0 = v$G$AB_9281_out0 && v$P$CD_10599_out0;
assign v$G5_4667_out0 = v$G$AB_9284_out0 && v$P$CD_10602_out0;
assign v$G5_4673_out0 = v$G$AB_9290_out0 && v$P$CD_10608_out0;
assign v$G5_4678_out0 = v$G$AB_9295_out0 && v$P$CD_10613_out0;
assign v$G1_5526_out0 = v$P$AB_2005_out0 && v$P$CD_10458_out0;
assign v$G1_5529_out0 = v$P$AB_2008_out0 && v$P$CD_10461_out0;
assign v$G1_5530_out0 = v$P$AB_2009_out0 && v$P$CD_10462_out0;
assign v$G1_5542_out0 = v$P$AB_2021_out0 && v$P$CD_10474_out0;
assign v$G1_5544_out0 = v$P$AB_2023_out0 && v$P$CD_10476_out0;
assign v$G1_5547_out0 = v$P$AB_2026_out0 && v$P$CD_10479_out0;
assign v$G1_5553_out0 = v$P$AB_2032_out0 && v$P$CD_10485_out0;
assign v$G1_5558_out0 = v$P$AB_2037_out0 && v$P$CD_10490_out0;
assign v$G1_5649_out0 = v$P$AB_2128_out0 && v$P$CD_10581_out0;
assign v$G1_5652_out0 = v$P$AB_2131_out0 && v$P$CD_10584_out0;
assign v$G1_5653_out0 = v$P$AB_2132_out0 && v$P$CD_10585_out0;
assign v$G1_5665_out0 = v$P$AB_2144_out0 && v$P$CD_10597_out0;
assign v$G1_5667_out0 = v$P$AB_2146_out0 && v$P$CD_10599_out0;
assign v$G1_5670_out0 = v$P$AB_2149_out0 && v$P$CD_10602_out0;
assign v$G1_5676_out0 = v$P$AB_2155_out0 && v$P$CD_10608_out0;
assign v$G1_5681_out0 = v$P$AB_2160_out0 && v$P$CD_10613_out0;
assign v$COUT_8111_out0 = v$A1_15214_out1;
assign v$G7_9639_out0 = v$G8_11399_out0 && v$P$CD_10458_out0;
assign v$G7_9642_out0 = v$G8_11402_out0 && v$P$CD_10461_out0;
assign v$G7_9643_out0 = v$G8_11403_out0 && v$P$CD_10462_out0;
assign v$G7_9655_out0 = v$G8_11415_out0 && v$P$CD_10474_out0;
assign v$G7_9657_out0 = v$G8_11417_out0 && v$P$CD_10476_out0;
assign v$G7_9660_out0 = v$G8_11420_out0 && v$P$CD_10479_out0;
assign v$G7_9666_out0 = v$G8_11426_out0 && v$P$CD_10485_out0;
assign v$G7_9671_out0 = v$G8_11431_out0 && v$P$CD_10490_out0;
assign v$G7_9762_out0 = v$G8_11522_out0 && v$P$CD_10581_out0;
assign v$G7_9765_out0 = v$G8_11525_out0 && v$P$CD_10584_out0;
assign v$G7_9766_out0 = v$G8_11526_out0 && v$P$CD_10585_out0;
assign v$G7_9778_out0 = v$G8_11538_out0 && v$P$CD_10597_out0;
assign v$G7_9780_out0 = v$G8_11540_out0 && v$P$CD_10599_out0;
assign v$G7_9783_out0 = v$G8_11543_out0 && v$P$CD_10602_out0;
assign v$G7_9789_out0 = v$G8_11549_out0 && v$P$CD_10608_out0;
assign v$G7_9794_out0 = v$G8_11554_out0 && v$P$CD_10613_out0;
assign v$C0_10692_out0 = v$GATE1_659_out0;
assign v$C0_10695_out0 = v$GATE1_662_out0;
assign v$MUX2_14827_out0 = v$EN_3875_out0 ? v$MUX1_2364_out0 : v$IN_3859_out0;
assign v$MUX2_14828_out0 = v$EN_3876_out0 ? v$MUX1_2374_out0 : v$IN_3862_out0;
assign v$_15111_out0 = { v$SUM$8_15776_out0,v$_10037_out0 };
assign v$SUM_15166_out0 = v$A1_15214_out0;
assign v$MUX6_16285_out0 = v$EQ6_5425_out0 ? v$SEL6_12472_out0 : v$MUX7_1227_out0;
assign v$MUX6_16286_out0 = v$EQ6_5426_out0 ? v$SEL6_12473_out0 : v$MUX7_1228_out0;
assign v$P$AD_691_out0 = v$G1_5526_out0;
assign v$P$AD_694_out0 = v$G1_5529_out0;
assign v$P$AD_695_out0 = v$G1_5530_out0;
assign v$P$AD_707_out0 = v$G1_5542_out0;
assign v$P$AD_709_out0 = v$G1_5544_out0;
assign v$P$AD_712_out0 = v$G1_5547_out0;
assign v$P$AD_718_out0 = v$G1_5553_out0;
assign v$P$AD_723_out0 = v$G1_5558_out0;
assign v$P$AD_814_out0 = v$G1_5649_out0;
assign v$P$AD_817_out0 = v$G1_5652_out0;
assign v$P$AD_818_out0 = v$G1_5653_out0;
assign v$P$AD_830_out0 = v$G1_5665_out0;
assign v$P$AD_832_out0 = v$G1_5667_out0;
assign v$P$AD_835_out0 = v$G1_5670_out0;
assign v$P$AD_841_out0 = v$G1_5676_out0;
assign v$P$AD_846_out0 = v$G1_5681_out0;
assign {v$A2A_1631_out1,v$A2A_1631_out0 } = v$A1_1710_out0 + v$B1_8123_out0 + v$C0_10692_out0;
assign {v$A2A_1634_out1,v$A2A_1634_out0 } = v$A1_1713_out0 + v$B1_8126_out0 + v$C0_10695_out0;
assign v$_1971_out0 = { v$SUM$7_7743_out0,v$_15111_out0 };
assign v$SUM_3466_out0 = v$SUM_15166_out0;
assign v$MUX5_6928_out0 = v$EQ5_3315_out0 ? v$SEL5_15451_out0 : v$MUX6_16285_out0;
assign v$MUX5_6929_out0 = v$EQ5_3316_out0 ? v$SEL5_15452_out0 : v$MUX6_16286_out0;
assign v$C0_9374_out0 = v$C0_10692_out0;
assign v$C0_9377_out0 = v$C0_10695_out0;
assign v$COUT_10728_out0 = v$COUT_8111_out0;
assign v$G4_11115_out0 = v$G5_4523_out0 || v$G$CD_918_out0;
assign v$G4_11118_out0 = v$G5_4526_out0 || v$G$CD_921_out0;
assign v$G4_11119_out0 = v$G5_4527_out0 || v$G$CD_922_out0;
assign v$G4_11131_out0 = v$G5_4539_out0 || v$G$CD_934_out0;
assign v$G4_11133_out0 = v$G5_4541_out0 || v$G$CD_936_out0;
assign v$G4_11136_out0 = v$G5_4544_out0 || v$G$CD_939_out0;
assign v$G4_11142_out0 = v$G5_4550_out0 || v$G$CD_945_out0;
assign v$G4_11147_out0 = v$G5_4555_out0 || v$G$CD_950_out0;
assign v$G4_11238_out0 = v$G5_4646_out0 || v$G$CD_1041_out0;
assign v$G4_11241_out0 = v$G5_4649_out0 || v$G$CD_1044_out0;
assign v$G4_11242_out0 = v$G5_4650_out0 || v$G$CD_1045_out0;
assign v$G4_11254_out0 = v$G5_4662_out0 || v$G$CD_1057_out0;
assign v$G4_11256_out0 = v$G5_4664_out0 || v$G$CD_1059_out0;
assign v$G4_11259_out0 = v$G5_4667_out0 || v$G$CD_1062_out0;
assign v$G4_11265_out0 = v$G5_4673_out0 || v$G$CD_1068_out0;
assign v$G4_11270_out0 = v$G5_4678_out0 || v$G$CD_1073_out0;
assign v$OUT_14916_out0 = v$MUX2_14827_out0;
assign v$OUT_14926_out0 = v$MUX2_14828_out0;
assign v$G6_437_out0 = v$G4_11115_out0 || v$G7_9639_out0;
assign v$G6_440_out0 = v$G4_11118_out0 || v$G7_9642_out0;
assign v$G6_441_out0 = v$G4_11119_out0 || v$G7_9643_out0;
assign v$G6_453_out0 = v$G4_11131_out0 || v$G7_9655_out0;
assign v$G6_455_out0 = v$G4_11133_out0 || v$G7_9657_out0;
assign v$G6_458_out0 = v$G4_11136_out0 || v$G7_9660_out0;
assign v$G6_464_out0 = v$G4_11142_out0 || v$G7_9666_out0;
assign v$G6_469_out0 = v$G4_11147_out0 || v$G7_9671_out0;
assign v$G6_560_out0 = v$G4_11238_out0 || v$G7_9762_out0;
assign v$G6_563_out0 = v$G4_11241_out0 || v$G7_9765_out0;
assign v$G6_564_out0 = v$G4_11242_out0 || v$G7_9766_out0;
assign v$G6_576_out0 = v$G4_11254_out0 || v$G7_9778_out0;
assign v$G6_578_out0 = v$G4_11256_out0 || v$G7_9780_out0;
assign v$G6_581_out0 = v$G4_11259_out0 || v$G7_9783_out0;
assign v$G6_587_out0 = v$G4_11265_out0 || v$G7_9789_out0;
assign v$G6_592_out0 = v$G4_11270_out0 || v$G7_9794_out0;
assign v$END1_1543_out0 = v$A2A_1631_out1;
assign v$END1_1546_out0 = v$A2A_1634_out1;
assign v$COUT$EXEC1_1594_out0 = v$COUT_10728_out0;
assign v$P$AB_2002_out0 = v$P$AD_707_out0;
assign v$P$AB_2003_out0 = v$P$AD_712_out0;
assign v$P$AB_2016_out0 = v$P$AD_695_out0;
assign v$P$AB_2018_out0 = v$P$AD_691_out0;
assign v$P$AB_2019_out0 = v$P$AD_718_out0;
assign v$P$AB_2022_out0 = v$P$AD_709_out0;
assign v$P$AB_2036_out0 = v$P$AD_694_out0;
assign v$P$AB_2041_out0 = v$P$AD_723_out0;
assign v$P$AB_2125_out0 = v$P$AD_830_out0;
assign v$P$AB_2126_out0 = v$P$AD_835_out0;
assign v$P$AB_2139_out0 = v$P$AD_818_out0;
assign v$P$AB_2141_out0 = v$P$AD_814_out0;
assign v$P$AB_2142_out0 = v$P$AD_841_out0;
assign v$P$AB_2145_out0 = v$P$AD_832_out0;
assign v$P$AB_2159_out0 = v$P$AD_817_out0;
assign v$P$AB_2164_out0 = v$P$AD_846_out0;
assign v$IN_5166_out0 = v$OUT_14916_out0;
assign v$IN_5176_out0 = v$OUT_14926_out0;
assign v$MUX4_7799_out0 = v$EQ4_18599_out0 ? v$SEL4_7321_out0 : v$MUX5_6928_out0;
assign v$MUX4_7800_out0 = v$EQ4_18600_out0 ? v$SEL4_7322_out0 : v$MUX5_6929_out0;
assign v$P$CD_10459_out0 = v$P$AD_718_out0;
assign v$P$CD_10463_out0 = v$P$AD_695_out0;
assign v$P$CD_10484_out0 = v$P$AD_709_out0;
assign v$P$CD_10487_out0 = v$P$AD_707_out0;
assign v$P$CD_10488_out0 = v$P$AD_723_out0;
assign v$P$CD_10492_out0 = v$P$AD_694_out0;
assign v$P$CD_10493_out0 = v$P$AD_712_out0;
assign v$P$CD_10582_out0 = v$P$AD_841_out0;
assign v$P$CD_10586_out0 = v$P$AD_818_out0;
assign v$P$CD_10607_out0 = v$P$AD_832_out0;
assign v$P$CD_10610_out0 = v$P$AD_830_out0;
assign v$P$CD_10611_out0 = v$P$AD_846_out0;
assign v$P$CD_10615_out0 = v$P$AD_817_out0;
assign v$P$CD_10616_out0 = v$P$AD_835_out0;
assign v$_12651_out0 = { v$SUM$6_12912_out0,v$_1971_out0 };
assign v$_13437_out0 = { v$A1A_11660_out0,v$A2A_1631_out0 };
assign v$_13440_out0 = { v$A1A_11663_out0,v$A2A_1634_out0 };
assign v$G$AD_17090_out0 = v$G4_11115_out0;
assign v$G$AD_17093_out0 = v$G4_11118_out0;
assign v$G$AD_17094_out0 = v$G4_11119_out0;
assign v$G$AD_17106_out0 = v$G4_11131_out0;
assign v$G$AD_17108_out0 = v$G4_11133_out0;
assign v$G$AD_17111_out0 = v$G4_11136_out0;
assign v$G$AD_17117_out0 = v$G4_11142_out0;
assign v$G$AD_17122_out0 = v$G4_11147_out0;
assign v$G$AD_17213_out0 = v$G4_11238_out0;
assign v$G$AD_17216_out0 = v$G4_11241_out0;
assign v$G$AD_17217_out0 = v$G4_11242_out0;
assign v$G$AD_17229_out0 = v$G4_11254_out0;
assign v$G$AD_17231_out0 = v$G4_11256_out0;
assign v$G$AD_17234_out0 = v$G4_11259_out0;
assign v$G$AD_17240_out0 = v$G4_11265_out0;
assign v$G$AD_17245_out0 = v$G4_11270_out0;
assign v$SUM$EXEC1_18543_out0 = v$SUM_3466_out0;
assign v$G$CD_919_out0 = v$G$AD_17117_out0;
assign v$G$CD_923_out0 = v$G$AD_17094_out0;
assign v$G$CD_944_out0 = v$G$AD_17108_out0;
assign v$G$CD_947_out0 = v$G$AD_17106_out0;
assign v$G$CD_948_out0 = v$G$AD_17122_out0;
assign v$G$CD_952_out0 = v$G$AD_17093_out0;
assign v$G$CD_953_out0 = v$G$AD_17111_out0;
assign v$G$CD_1042_out0 = v$G$AD_17240_out0;
assign v$G$CD_1046_out0 = v$G$AD_17217_out0;
assign v$G$CD_1067_out0 = v$G$AD_17231_out0;
assign v$G$CD_1070_out0 = v$G$AD_17229_out0;
assign v$G$CD_1071_out0 = v$G$AD_17245_out0;
assign v$G$CD_1075_out0 = v$G$AD_17216_out0;
assign v$G$CD_1076_out0 = v$G$AD_17234_out0;
assign v$_5491_out0 = { v$SUM$5_7817_out0,v$_12651_out0 };
assign v$G1_5523_out0 = v$P$AB_2002_out0 && v$P$CD_10455_out0;
assign v$G1_5524_out0 = v$P$AB_2003_out0 && v$P$CD_10456_out0;
assign v$G1_5537_out0 = v$P$AB_2016_out0 && v$P$CD_10469_out0;
assign v$G1_5539_out0 = v$P$AB_2018_out0 && v$P$CD_10471_out0;
assign v$G1_5540_out0 = v$P$AB_2019_out0 && v$P$CD_10472_out0;
assign v$G1_5543_out0 = v$P$AB_2022_out0 && v$P$CD_10475_out0;
assign v$G1_5557_out0 = v$P$AB_2036_out0 && v$P$CD_10489_out0;
assign v$G1_5562_out0 = v$P$AB_2041_out0 && v$P$CD_10494_out0;
assign v$G1_5646_out0 = v$P$AB_2125_out0 && v$P$CD_10578_out0;
assign v$G1_5647_out0 = v$P$AB_2126_out0 && v$P$CD_10579_out0;
assign v$G1_5660_out0 = v$P$AB_2139_out0 && v$P$CD_10592_out0;
assign v$G1_5662_out0 = v$P$AB_2141_out0 && v$P$CD_10594_out0;
assign v$G1_5663_out0 = v$P$AB_2142_out0 && v$P$CD_10595_out0;
assign v$G1_5666_out0 = v$P$AB_2145_out0 && v$P$CD_10598_out0;
assign v$G1_5680_out0 = v$P$AB_2159_out0 && v$P$CD_10612_out0;
assign v$G1_5685_out0 = v$P$AB_2164_out0 && v$P$CD_10617_out0;
assign v$COUTD_6697_out0 = v$G6_437_out0;
assign v$COUTD_6700_out0 = v$G6_440_out0;
assign v$COUTD_6701_out0 = v$G6_441_out0;
assign v$COUTD_6713_out0 = v$G6_453_out0;
assign v$COUTD_6715_out0 = v$G6_455_out0;
assign v$COUTD_6718_out0 = v$G6_458_out0;
assign v$COUTD_6724_out0 = v$G6_464_out0;
assign v$COUTD_6729_out0 = v$G6_469_out0;
assign v$COUTD_6820_out0 = v$G6_560_out0;
assign v$COUTD_6823_out0 = v$G6_563_out0;
assign v$COUTD_6824_out0 = v$G6_564_out0;
assign v$COUTD_6836_out0 = v$G6_576_out0;
assign v$COUTD_6838_out0 = v$G6_578_out0;
assign v$COUTD_6841_out0 = v$G6_581_out0;
assign v$COUTD_6847_out0 = v$G6_587_out0;
assign v$COUTD_6852_out0 = v$G6_592_out0;
assign v$MUX3_7600_out0 = v$EQ3_1816_out0 ? v$SEL3_11729_out0 : v$MUX4_7799_out0;
assign v$MUX3_7601_out0 = v$EQ3_1817_out0 ? v$SEL3_11730_out0 : v$MUX4_7800_out0;
assign v$G$AB_9137_out0 = v$G$AD_17106_out0;
assign v$G$AB_9138_out0 = v$G$AD_17111_out0;
assign v$G$AB_9151_out0 = v$G$AD_17094_out0;
assign v$G$AB_9153_out0 = v$G$AD_17090_out0;
assign v$G$AB_9154_out0 = v$G$AD_17117_out0;
assign v$G$AB_9157_out0 = v$G$AD_17108_out0;
assign v$G$AB_9171_out0 = v$G$AD_17093_out0;
assign v$G$AB_9176_out0 = v$G$AD_17122_out0;
assign v$G$AB_9260_out0 = v$G$AD_17229_out0;
assign v$G$AB_9261_out0 = v$G$AD_17234_out0;
assign v$G$AB_9274_out0 = v$G$AD_17217_out0;
assign v$G$AB_9276_out0 = v$G$AD_17213_out0;
assign v$G$AB_9277_out0 = v$G$AD_17240_out0;
assign v$G$AB_9280_out0 = v$G$AD_17231_out0;
assign v$G$AB_9294_out0 = v$G$AD_17216_out0;
assign v$G$AB_9299_out0 = v$G$AD_17245_out0;
assign v$IN_11784_out0 = v$IN_5166_out0;
assign v$IN_11786_out0 = v$IN_5176_out0;
assign v$_18087_out0 = { v$SUM$11_17033_out0,v$SUM$EXEC1_18543_out0 };
assign v$P$AD_688_out0 = v$G1_5523_out0;
assign v$P$AD_689_out0 = v$G1_5524_out0;
assign v$P$AD_702_out0 = v$G1_5537_out0;
assign v$P$AD_704_out0 = v$G1_5539_out0;
assign v$P$AD_705_out0 = v$G1_5540_out0;
assign v$P$AD_708_out0 = v$G1_5543_out0;
assign v$P$AD_722_out0 = v$G1_5557_out0;
assign v$P$AD_727_out0 = v$G1_5562_out0;
assign v$P$AD_811_out0 = v$G1_5646_out0;
assign v$P$AD_812_out0 = v$G1_5647_out0;
assign v$P$AD_825_out0 = v$G1_5660_out0;
assign v$P$AD_827_out0 = v$G1_5662_out0;
assign v$P$AD_828_out0 = v$G1_5663_out0;
assign v$P$AD_831_out0 = v$G1_5666_out0;
assign v$P$AD_845_out0 = v$G1_5680_out0;
assign v$P$AD_850_out0 = v$G1_5685_out0;
assign v$G5_4520_out0 = v$G$AB_9137_out0 && v$P$CD_10455_out0;
assign v$G5_4521_out0 = v$G$AB_9138_out0 && v$P$CD_10456_out0;
assign v$G5_4534_out0 = v$G$AB_9151_out0 && v$P$CD_10469_out0;
assign v$G5_4536_out0 = v$G$AB_9153_out0 && v$P$CD_10471_out0;
assign v$G5_4537_out0 = v$G$AB_9154_out0 && v$P$CD_10472_out0;
assign v$G5_4540_out0 = v$G$AB_9157_out0 && v$P$CD_10475_out0;
assign v$G5_4554_out0 = v$G$AB_9171_out0 && v$P$CD_10489_out0;
assign v$G5_4559_out0 = v$G$AB_9176_out0 && v$P$CD_10494_out0;
assign v$G5_4643_out0 = v$G$AB_9260_out0 && v$P$CD_10578_out0;
assign v$G5_4644_out0 = v$G$AB_9261_out0 && v$P$CD_10579_out0;
assign v$G5_4657_out0 = v$G$AB_9274_out0 && v$P$CD_10592_out0;
assign v$G5_4659_out0 = v$G$AB_9276_out0 && v$P$CD_10594_out0;
assign v$G5_4660_out0 = v$G$AB_9277_out0 && v$P$CD_10595_out0;
assign v$G5_4663_out0 = v$G$AB_9280_out0 && v$P$CD_10598_out0;
assign v$G5_4677_out0 = v$G$AB_9294_out0 && v$P$CD_10612_out0;
assign v$G5_4682_out0 = v$G$AB_9299_out0 && v$P$CD_10617_out0;
assign v$CINA_8465_out0 = v$COUTD_6713_out0;
assign v$CINA_8466_out0 = v$COUTD_6718_out0;
assign v$CINA_8479_out0 = v$COUTD_6701_out0;
assign v$CINA_8481_out0 = v$COUTD_6697_out0;
assign v$CINA_8482_out0 = v$COUTD_6724_out0;
assign v$CINA_8485_out0 = v$COUTD_6715_out0;
assign v$CINA_8499_out0 = v$COUTD_6700_out0;
assign v$CINA_8504_out0 = v$COUTD_6729_out0;
assign v$CINA_8588_out0 = v$COUTD_6836_out0;
assign v$CINA_8589_out0 = v$COUTD_6841_out0;
assign v$CINA_8602_out0 = v$COUTD_6824_out0;
assign v$CINA_8604_out0 = v$COUTD_6820_out0;
assign v$CINA_8605_out0 = v$COUTD_6847_out0;
assign v$CINA_8608_out0 = v$COUTD_6838_out0;
assign v$CINA_8622_out0 = v$COUTD_6823_out0;
assign v$CINA_8627_out0 = v$COUTD_6852_out0;
assign v$SEL1_8714_out0 = v$IN_11784_out0[23:2];
assign v$SEL1_8724_out0 = v$IN_11786_out0[23:2];
assign v$_9488_out0 = { v$SUM$4_15246_out0,v$_5491_out0 };
assign v$_11764_out0 = { v$SUM$10_14308_out0,v$_18087_out0 };
assign v$MUX2_13608_out0 = v$EQ2_14208_out0 ? v$SEL2_13321_out0 : v$MUX3_7600_out0;
assign v$MUX2_13609_out0 = v$EQ2_14209_out0 ? v$SEL2_13322_out0 : v$MUX3_7601_out0;
assign v$SEL1_15405_out0 = v$IN_11784_out0[21:0];
assign v$SEL1_15415_out0 = v$IN_11786_out0[21:0];
assign v$C1_16781_out0 = v$COUTD_6697_out0;
assign v$C1_16784_out0 = v$COUTD_6820_out0;
assign v$P$AB_2001_out0 = v$P$AD_689_out0;
assign v$P$AB_2006_out0 = v$P$AD_704_out0;
assign v$P$AB_2012_out0 = v$P$AD_704_out0;
assign v$P$AB_2015_out0 = v$P$AD_722_out0;
assign v$P$AB_2020_out0 = v$P$AD_688_out0;
assign v$P$AB_2033_out0 = v$P$AD_704_out0;
assign v$P$AB_2124_out0 = v$P$AD_812_out0;
assign v$P$AB_2129_out0 = v$P$AD_827_out0;
assign v$P$AB_2135_out0 = v$P$AD_827_out0;
assign v$P$AB_2138_out0 = v$P$AD_845_out0;
assign v$P$AB_2143_out0 = v$P$AD_811_out0;
assign v$P$AB_2156_out0 = v$P$AD_827_out0;
assign v$MUX1_2865_out0 = v$EQ1_13414_out0 ? v$SEL1_7088_out0 : v$MUX2_13608_out0;
assign v$MUX1_2866_out0 = v$EQ1_13415_out0 ? v$SEL1_7089_out0 : v$MUX2_13609_out0;
assign v$_4264_out0 = { v$C2_122_out0,v$SEL1_15405_out0 };
assign v$_4274_out0 = { v$C2_132_out0,v$SEL1_15415_out0 };
assign v$_7621_out0 = { v$SUM$9_197_out0,v$_11764_out0 };
assign v$_8999_out0 = { v$SEL1_8714_out0,v$C1_5980_out0 };
assign v$_9009_out0 = { v$SEL1_8724_out0,v$C1_5990_out0 };
assign v$P$CD_10454_out0 = v$P$AD_727_out0;
assign v$P$CD_10460_out0 = v$P$AD_689_out0;
assign v$P$CD_10468_out0 = v$P$AD_702_out0;
assign v$P$CD_10473_out0 = v$P$AD_708_out0;
assign v$P$CD_10477_out0 = v$P$AD_722_out0;
assign v$P$CD_10478_out0 = v$P$AD_688_out0;
assign v$P$CD_10486_out0 = v$P$AD_705_out0;
assign v$P$CD_10577_out0 = v$P$AD_850_out0;
assign v$P$CD_10583_out0 = v$P$AD_812_out0;
assign v$P$CD_10591_out0 = v$P$AD_825_out0;
assign v$P$CD_10596_out0 = v$P$AD_831_out0;
assign v$P$CD_10600_out0 = v$P$AD_845_out0;
assign v$P$CD_10601_out0 = v$P$AD_811_out0;
assign v$P$CD_10609_out0 = v$P$AD_828_out0;
assign v$G4_11112_out0 = v$G5_4520_out0 || v$G$CD_915_out0;
assign v$G4_11113_out0 = v$G5_4521_out0 || v$G$CD_916_out0;
assign v$G4_11126_out0 = v$G5_4534_out0 || v$G$CD_929_out0;
assign v$G4_11128_out0 = v$G5_4536_out0 || v$G$CD_931_out0;
assign v$G4_11129_out0 = v$G5_4537_out0 || v$G$CD_932_out0;
assign v$G4_11132_out0 = v$G5_4540_out0 || v$G$CD_935_out0;
assign v$G4_11146_out0 = v$G5_4554_out0 || v$G$CD_949_out0;
assign v$G4_11151_out0 = v$G5_4559_out0 || v$G$CD_954_out0;
assign v$G4_11235_out0 = v$G5_4643_out0 || v$G$CD_1038_out0;
assign v$G4_11236_out0 = v$G5_4644_out0 || v$G$CD_1039_out0;
assign v$G4_11249_out0 = v$G5_4657_out0 || v$G$CD_1052_out0;
assign v$G4_11251_out0 = v$G5_4659_out0 || v$G$CD_1054_out0;
assign v$G4_11252_out0 = v$G5_4660_out0 || v$G$CD_1055_out0;
assign v$G4_11255_out0 = v$G5_4663_out0 || v$G$CD_1058_out0;
assign v$G4_11269_out0 = v$G5_4677_out0 || v$G$CD_1072_out0;
assign v$G4_11274_out0 = v$G5_4682_out0 || v$G$CD_1077_out0;
assign v$G8_11396_out0 = v$CINA_8465_out0 && v$P$AB_2002_out0;
assign v$G8_11397_out0 = v$CINA_8466_out0 && v$P$AB_2003_out0;
assign v$G8_11410_out0 = v$CINA_8479_out0 && v$P$AB_2016_out0;
assign v$G8_11412_out0 = v$CINA_8481_out0 && v$P$AB_2018_out0;
assign v$G8_11413_out0 = v$CINA_8482_out0 && v$P$AB_2019_out0;
assign v$G8_11416_out0 = v$CINA_8485_out0 && v$P$AB_2022_out0;
assign v$G8_11430_out0 = v$CINA_8499_out0 && v$P$AB_2036_out0;
assign v$G8_11435_out0 = v$CINA_8504_out0 && v$P$AB_2041_out0;
assign v$G8_11519_out0 = v$CINA_8588_out0 && v$P$AB_2125_out0;
assign v$G8_11520_out0 = v$CINA_8589_out0 && v$P$AB_2126_out0;
assign v$G8_11533_out0 = v$CINA_8602_out0 && v$P$AB_2139_out0;
assign v$G8_11535_out0 = v$CINA_8604_out0 && v$P$AB_2141_out0;
assign v$G8_11536_out0 = v$CINA_8605_out0 && v$P$AB_2142_out0;
assign v$G8_11539_out0 = v$CINA_8608_out0 && v$P$AB_2145_out0;
assign v$G8_11553_out0 = v$CINA_8622_out0 && v$P$AB_2159_out0;
assign v$G8_11558_out0 = v$CINA_8627_out0 && v$P$AB_2164_out0;
assign v$C1_11849_out0 = v$C1_16781_out0;
assign v$C1_11852_out0 = v$C1_16784_out0;
assign {v$A3A_11951_out1,v$A3A_11951_out0 } = v$A2_18266_out0 + v$B2_3113_out0 + v$C1_16781_out0;
assign {v$A3A_11954_out1,v$A3A_11954_out0 } = v$A2_18269_out0 + v$B2_3116_out0 + v$C1_16784_out0;
assign v$_16504_out0 = { v$SUM$3_7904_out0,v$_9488_out0 };
assign v$MUX1_2368_out0 = v$LEFT$SHIT_3060_out0 ? v$_4264_out0 : v$_8999_out0;
assign v$MUX1_2378_out0 = v$LEFT$SHIT_3070_out0 ? v$_4274_out0 : v$_9009_out0;
assign v$_4158_out0 = { v$SUM$8_15776_out0,v$_7621_out0 };
assign v$END2_5234_out0 = v$A3A_11951_out1;
assign v$END2_5237_out0 = v$A3A_11954_out1;
assign v$G1_5522_out0 = v$P$AB_2001_out0 && v$P$CD_10454_out0;
assign v$G1_5527_out0 = v$P$AB_2006_out0 && v$P$CD_10459_out0;
assign v$G1_5533_out0 = v$P$AB_2012_out0 && v$P$CD_10465_out0;
assign v$G1_5536_out0 = v$P$AB_2015_out0 && v$P$CD_10468_out0;
assign v$G1_5541_out0 = v$P$AB_2020_out0 && v$P$CD_10473_out0;
assign v$G1_5554_out0 = v$P$AB_2033_out0 && v$P$CD_10486_out0;
assign v$G1_5645_out0 = v$P$AB_2124_out0 && v$P$CD_10577_out0;
assign v$G1_5650_out0 = v$P$AB_2129_out0 && v$P$CD_10582_out0;
assign v$G1_5656_out0 = v$P$AB_2135_out0 && v$P$CD_10588_out0;
assign v$G1_5659_out0 = v$P$AB_2138_out0 && v$P$CD_10591_out0;
assign v$G1_5664_out0 = v$P$AB_2143_out0 && v$P$CD_10596_out0;
assign v$G1_5677_out0 = v$P$AB_2156_out0 && v$P$CD_10609_out0;
assign v$MUX25_8404_out0 = v$G2_11902_out0 ? v$C2_15178_out0 : v$MUX1_2865_out0;
assign v$MUX25_8405_out0 = v$G2_11903_out0 ? v$C2_15179_out0 : v$MUX1_2866_out0;
assign v$_8906_out0 = { v$C0_9374_out0,v$C1_11849_out0 };
assign v$_8909_out0 = { v$C0_9377_out0,v$C1_11852_out0 };
assign v$G7_9636_out0 = v$G8_11396_out0 && v$P$CD_10455_out0;
assign v$G7_9637_out0 = v$G8_11397_out0 && v$P$CD_10456_out0;
assign v$G7_9650_out0 = v$G8_11410_out0 && v$P$CD_10469_out0;
assign v$G7_9652_out0 = v$G8_11412_out0 && v$P$CD_10471_out0;
assign v$G7_9653_out0 = v$G8_11413_out0 && v$P$CD_10472_out0;
assign v$G7_9656_out0 = v$G8_11416_out0 && v$P$CD_10475_out0;
assign v$G7_9670_out0 = v$G8_11430_out0 && v$P$CD_10489_out0;
assign v$G7_9675_out0 = v$G8_11435_out0 && v$P$CD_10494_out0;
assign v$G7_9759_out0 = v$G8_11519_out0 && v$P$CD_10578_out0;
assign v$G7_9760_out0 = v$G8_11520_out0 && v$P$CD_10579_out0;
assign v$G7_9773_out0 = v$G8_11533_out0 && v$P$CD_10592_out0;
assign v$G7_9775_out0 = v$G8_11535_out0 && v$P$CD_10594_out0;
assign v$G7_9776_out0 = v$G8_11536_out0 && v$P$CD_10595_out0;
assign v$G7_9779_out0 = v$G8_11539_out0 && v$P$CD_10598_out0;
assign v$G7_9793_out0 = v$G8_11553_out0 && v$P$CD_10612_out0;
assign v$G7_9798_out0 = v$G8_11558_out0 && v$P$CD_10617_out0;
assign v$_16340_out0 = { v$SUM$2_9082_out0,v$_16504_out0 };
assign v$G$AD_17087_out0 = v$G4_11112_out0;
assign v$G$AD_17088_out0 = v$G4_11113_out0;
assign v$G$AD_17101_out0 = v$G4_11126_out0;
assign v$G$AD_17103_out0 = v$G4_11128_out0;
assign v$G$AD_17104_out0 = v$G4_11129_out0;
assign v$G$AD_17107_out0 = v$G4_11132_out0;
assign v$G$AD_17121_out0 = v$G4_11146_out0;
assign v$G$AD_17126_out0 = v$G4_11151_out0;
assign v$G$AD_17210_out0 = v$G4_11235_out0;
assign v$G$AD_17211_out0 = v$G4_11236_out0;
assign v$G$AD_17224_out0 = v$G4_11249_out0;
assign v$G$AD_17226_out0 = v$G4_11251_out0;
assign v$G$AD_17227_out0 = v$G4_11252_out0;
assign v$G$AD_17230_out0 = v$G4_11255_out0;
assign v$G$AD_17244_out0 = v$G4_11269_out0;
assign v$G$AD_17249_out0 = v$G4_11274_out0;
assign v$G6_434_out0 = v$G4_11112_out0 || v$G7_9636_out0;
assign v$G6_435_out0 = v$G4_11113_out0 || v$G7_9637_out0;
assign v$G6_448_out0 = v$G4_11126_out0 || v$G7_9650_out0;
assign v$G6_450_out0 = v$G4_11128_out0 || v$G7_9652_out0;
assign v$G6_451_out0 = v$G4_11129_out0 || v$G7_9653_out0;
assign v$G6_454_out0 = v$G4_11132_out0 || v$G7_9656_out0;
assign v$G6_468_out0 = v$G4_11146_out0 || v$G7_9670_out0;
assign v$G6_473_out0 = v$G4_11151_out0 || v$G7_9675_out0;
assign v$G6_557_out0 = v$G4_11235_out0 || v$G7_9759_out0;
assign v$G6_558_out0 = v$G4_11236_out0 || v$G7_9760_out0;
assign v$G6_571_out0 = v$G4_11249_out0 || v$G7_9773_out0;
assign v$G6_573_out0 = v$G4_11251_out0 || v$G7_9775_out0;
assign v$G6_574_out0 = v$G4_11252_out0 || v$G7_9776_out0;
assign v$G6_577_out0 = v$G4_11255_out0 || v$G7_9779_out0;
assign v$G6_591_out0 = v$G4_11269_out0 || v$G7_9793_out0;
assign v$G6_596_out0 = v$G4_11274_out0 || v$G7_9798_out0;
assign v$P$AD_687_out0 = v$G1_5522_out0;
assign v$P$AD_692_out0 = v$G1_5527_out0;
assign v$P$AD_698_out0 = v$G1_5533_out0;
assign v$P$AD_701_out0 = v$G1_5536_out0;
assign v$P$AD_706_out0 = v$G1_5541_out0;
assign v$P$AD_719_out0 = v$G1_5554_out0;
assign v$P$AD_810_out0 = v$G1_5645_out0;
assign v$P$AD_815_out0 = v$G1_5650_out0;
assign v$P$AD_821_out0 = v$G1_5656_out0;
assign v$P$AD_824_out0 = v$G1_5659_out0;
assign v$P$AD_829_out0 = v$G1_5664_out0;
assign v$P$AD_842_out0 = v$G1_5677_out0;
assign v$G$CD_914_out0 = v$G$AD_17126_out0;
assign v$G$CD_920_out0 = v$G$AD_17088_out0;
assign v$G$CD_928_out0 = v$G$AD_17101_out0;
assign v$G$CD_933_out0 = v$G$AD_17107_out0;
assign v$G$CD_937_out0 = v$G$AD_17121_out0;
assign v$G$CD_938_out0 = v$G$AD_17087_out0;
assign v$G$CD_946_out0 = v$G$AD_17104_out0;
assign v$G$CD_1037_out0 = v$G$AD_17249_out0;
assign v$G$CD_1043_out0 = v$G$AD_17211_out0;
assign v$G$CD_1051_out0 = v$G$AD_17224_out0;
assign v$G$CD_1056_out0 = v$G$AD_17230_out0;
assign v$G$CD_1060_out0 = v$G$AD_17244_out0;
assign v$G$CD_1061_out0 = v$G$AD_17210_out0;
assign v$G$CD_1069_out0 = v$G$AD_17227_out0;
assign v$MUX2_2478_out0 = v$EN_7876_out0 ? v$MUX1_2368_out0 : v$IN_11784_out0;
assign v$MUX2_2480_out0 = v$EN_7878_out0 ? v$MUX1_2378_out0 : v$IN_11786_out0;
assign v$G$AB_9136_out0 = v$G$AD_17088_out0;
assign v$G$AB_9141_out0 = v$G$AD_17103_out0;
assign v$G$AB_9147_out0 = v$G$AD_17103_out0;
assign v$G$AB_9150_out0 = v$G$AD_17121_out0;
assign v$G$AB_9155_out0 = v$G$AD_17087_out0;
assign v$G$AB_9168_out0 = v$G$AD_17103_out0;
assign v$G$AB_9259_out0 = v$G$AD_17211_out0;
assign v$G$AB_9264_out0 = v$G$AD_17226_out0;
assign v$G$AB_9270_out0 = v$G$AD_17226_out0;
assign v$G$AB_9273_out0 = v$G$AD_17244_out0;
assign v$G$AB_9278_out0 = v$G$AD_17210_out0;
assign v$G$AB_9291_out0 = v$G$AD_17226_out0;
assign v$OUT_9476_out0 = v$MUX25_8404_out0;
assign v$OUT_9477_out0 = v$MUX25_8405_out0;
assign v$_13316_out0 = { v$SUM$1_10360_out0,v$_16340_out0 };
assign v$_16351_out0 = { v$SUM$7_7743_out0,v$_4158_out0 };
assign v$P$AB_2007_out0 = v$P$AD_719_out0;
assign v$P$AB_2011_out0 = v$P$AD_719_out0;
assign v$P$AB_2030_out0 = v$P$AD_719_out0;
assign v$P$AB_2038_out0 = v$P$AD_706_out0;
assign v$P$AB_2040_out0 = v$P$AD_719_out0;
assign v$P$AB_2130_out0 = v$P$AD_842_out0;
assign v$P$AB_2134_out0 = v$P$AD_842_out0;
assign v$P$AB_2153_out0 = v$P$AD_842_out0;
assign v$P$AB_2161_out0 = v$P$AD_829_out0;
assign v$P$AB_2163_out0 = v$P$AD_842_out0;
assign v$_2533_out0 = { v$SEL8_12749_out0,v$_13316_out0 };
assign {v$A1_2662_out1,v$A1_2662_out0 } = v$LARGER$EXP_10274_out0 + v$SMALLER$EXP_2941_out0 + v$OUT_9476_out0;
assign {v$A1_2663_out1,v$A1_2663_out0 } = v$LARGER$EXP_10275_out0 + v$SMALLER$EXP_2942_out0 + v$OUT_9477_out0;
assign v$G5_4519_out0 = v$G$AB_9136_out0 && v$P$CD_10454_out0;
assign v$G5_4524_out0 = v$G$AB_9141_out0 && v$P$CD_10459_out0;
assign v$G5_4530_out0 = v$G$AB_9147_out0 && v$P$CD_10465_out0;
assign v$G5_4533_out0 = v$G$AB_9150_out0 && v$P$CD_10468_out0;
assign v$G5_4538_out0 = v$G$AB_9155_out0 && v$P$CD_10473_out0;
assign v$G5_4551_out0 = v$G$AB_9168_out0 && v$P$CD_10486_out0;
assign v$G5_4642_out0 = v$G$AB_9259_out0 && v$P$CD_10577_out0;
assign v$G5_4647_out0 = v$G$AB_9264_out0 && v$P$CD_10582_out0;
assign v$G5_4653_out0 = v$G$AB_9270_out0 && v$P$CD_10588_out0;
assign v$G5_4656_out0 = v$G$AB_9273_out0 && v$P$CD_10591_out0;
assign v$G5_4661_out0 = v$G$AB_9278_out0 && v$P$CD_10596_out0;
assign v$G5_4674_out0 = v$G$AB_9291_out0 && v$P$CD_10609_out0;
assign v$COUTD_6694_out0 = v$G6_434_out0;
assign v$COUTD_6695_out0 = v$G6_435_out0;
assign v$COUTD_6708_out0 = v$G6_448_out0;
assign v$COUTD_6710_out0 = v$G6_450_out0;
assign v$COUTD_6711_out0 = v$G6_451_out0;
assign v$COUTD_6714_out0 = v$G6_454_out0;
assign v$COUTD_6728_out0 = v$G6_468_out0;
assign v$COUTD_6733_out0 = v$G6_473_out0;
assign v$COUTD_6817_out0 = v$G6_557_out0;
assign v$COUTD_6818_out0 = v$G6_558_out0;
assign v$COUTD_6831_out0 = v$G6_571_out0;
assign v$COUTD_6833_out0 = v$G6_573_out0;
assign v$COUTD_6834_out0 = v$G6_574_out0;
assign v$COUTD_6837_out0 = v$G6_577_out0;
assign v$COUTD_6851_out0 = v$G6_591_out0;
assign v$COUTD_6856_out0 = v$G6_596_out0;
assign v$P$CD_10457_out0 = v$P$AD_706_out0;
assign v$P$CD_10483_out0 = v$P$AD_687_out0;
assign v$P$CD_10491_out0 = v$P$AD_701_out0;
assign v$P$CD_10580_out0 = v$P$AD_829_out0;
assign v$P$CD_10606_out0 = v$P$AD_810_out0;
assign v$P$CD_10614_out0 = v$P$AD_824_out0;
assign v$END11_12090_out0 = v$P$AD_698_out0;
assign v$END11_12093_out0 = v$P$AD_821_out0;
assign v$OUT_14920_out0 = v$MUX2_2478_out0;
assign v$OUT_14930_out0 = v$MUX2_2480_out0;
assign v$_17404_out0 = { v$SUM$6_12912_out0,v$_16351_out0 };
assign v$END13_18067_out0 = v$P$AD_692_out0;
assign v$END13_18070_out0 = v$P$AD_815_out0;
assign v$END1_1291_out0 = v$COUTD_6733_out0;
assign v$END1_1294_out0 = v$COUTD_6856_out0;
assign v$C2_2686_out0 = v$COUTD_6710_out0;
assign v$C2_2689_out0 = v$COUTD_6833_out0;
assign v$END_3319_out0 = v$COUTD_6711_out0;
assign v$END_3322_out0 = v$COUTD_6834_out0;
assign v$END3_3445_out0 = v$COUTD_6708_out0;
assign v$END3_3448_out0 = v$COUTD_6831_out0;
assign v$IN_5164_out0 = v$OUT_14920_out0;
assign v$IN_5174_out0 = v$OUT_14930_out0;
assign v$G1_5528_out0 = v$P$AB_2007_out0 && v$P$CD_10460_out0;
assign v$G1_5532_out0 = v$P$AB_2011_out0 && v$P$CD_10464_out0;
assign v$G1_5551_out0 = v$P$AB_2030_out0 && v$P$CD_10483_out0;
assign v$G1_5559_out0 = v$P$AB_2038_out0 && v$P$CD_10491_out0;
assign v$G1_5561_out0 = v$P$AB_2040_out0 && v$P$CD_10493_out0;
assign v$G1_5651_out0 = v$P$AB_2130_out0 && v$P$CD_10583_out0;
assign v$G1_5655_out0 = v$P$AB_2134_out0 && v$P$CD_10587_out0;
assign v$G1_5674_out0 = v$P$AB_2153_out0 && v$P$CD_10606_out0;
assign v$G1_5682_out0 = v$P$AB_2161_out0 && v$P$CD_10614_out0;
assign v$G1_5684_out0 = v$P$AB_2163_out0 && v$P$CD_10616_out0;
assign v$END2_7751_out0 = v$COUTD_6714_out0;
assign v$END2_7754_out0 = v$COUTD_6837_out0;
assign v$OUT_8212_out0 = v$_2533_out0;
assign v$_8260_out0 = { v$SUM$5_7817_out0,v$_17404_out0 };
assign v$CINA_8464_out0 = v$COUTD_6695_out0;
assign v$CINA_8469_out0 = v$COUTD_6710_out0;
assign v$CINA_8475_out0 = v$COUTD_6710_out0;
assign v$CINA_8478_out0 = v$COUTD_6728_out0;
assign v$CINA_8483_out0 = v$COUTD_6694_out0;
assign v$CINA_8496_out0 = v$COUTD_6710_out0;
assign v$CINA_8587_out0 = v$COUTD_6818_out0;
assign v$CINA_8592_out0 = v$COUTD_6833_out0;
assign v$CINA_8598_out0 = v$COUTD_6833_out0;
assign v$CINA_8601_out0 = v$COUTD_6851_out0;
assign v$CINA_8606_out0 = v$COUTD_6817_out0;
assign v$CINA_8619_out0 = v$COUTD_6833_out0;
assign v$END45_9057_out0 = v$COUTD_6728_out0;
assign v$END45_9060_out0 = v$COUTD_6851_out0;
assign {v$A2_10044_out1,v$A2_10044_out0 } = v$A1_2662_out0 + v$C1_5955_out0 + v$C2_16281_out0;
assign {v$A2_10045_out1,v$A2_10045_out0 } = v$A1_2663_out0 + v$C1_5956_out0 + v$C2_16282_out0;
assign v$G4_11111_out0 = v$G5_4519_out0 || v$G$CD_914_out0;
assign v$G4_11116_out0 = v$G5_4524_out0 || v$G$CD_919_out0;
assign v$G4_11122_out0 = v$G5_4530_out0 || v$G$CD_925_out0;
assign v$G4_11125_out0 = v$G5_4533_out0 || v$G$CD_928_out0;
assign v$G4_11130_out0 = v$G5_4538_out0 || v$G$CD_933_out0;
assign v$G4_11143_out0 = v$G5_4551_out0 || v$G$CD_946_out0;
assign v$G4_11234_out0 = v$G5_4642_out0 || v$G$CD_1037_out0;
assign v$G4_11239_out0 = v$G5_4647_out0 || v$G$CD_1042_out0;
assign v$G4_11245_out0 = v$G5_4653_out0 || v$G$CD_1048_out0;
assign v$G4_11248_out0 = v$G5_4656_out0 || v$G$CD_1051_out0;
assign v$G4_11253_out0 = v$G5_4661_out0 || v$G$CD_1056_out0;
assign v$G4_11266_out0 = v$G5_4674_out0 || v$G$CD_1069_out0;
assign v$NOT$USED$CARRY_18775_out0 = v$A1_2662_out1;
assign v$NOT$USED$CARRY_18776_out0 = v$A1_2663_out1;
assign v$P$AD_693_out0 = v$G1_5528_out0;
assign v$P$AD_697_out0 = v$G1_5532_out0;
assign v$P$AD_716_out0 = v$G1_5551_out0;
assign v$P$AD_724_out0 = v$G1_5559_out0;
assign v$P$AD_726_out0 = v$G1_5561_out0;
assign v$P$AD_816_out0 = v$G1_5651_out0;
assign v$P$AD_820_out0 = v$G1_5655_out0;
assign v$P$AD_839_out0 = v$G1_5674_out0;
assign v$P$AD_847_out0 = v$G1_5682_out0;
assign v$P$AD_849_out0 = v$G1_5684_out0;
assign v$MULTIPLIER$OUT_9344_out0 = v$OUT_8212_out0;
assign v$G8_11395_out0 = v$CINA_8464_out0 && v$P$AB_2001_out0;
assign v$G8_11400_out0 = v$CINA_8469_out0 && v$P$AB_2006_out0;
assign v$G8_11406_out0 = v$CINA_8475_out0 && v$P$AB_2012_out0;
assign v$G8_11409_out0 = v$CINA_8478_out0 && v$P$AB_2015_out0;
assign v$G8_11414_out0 = v$CINA_8483_out0 && v$P$AB_2020_out0;
assign v$G8_11427_out0 = v$CINA_8496_out0 && v$P$AB_2033_out0;
assign v$G8_11518_out0 = v$CINA_8587_out0 && v$P$AB_2124_out0;
assign v$G8_11523_out0 = v$CINA_8592_out0 && v$P$AB_2129_out0;
assign v$G8_11529_out0 = v$CINA_8598_out0 && v$P$AB_2135_out0;
assign v$G8_11532_out0 = v$CINA_8601_out0 && v$P$AB_2138_out0;
assign v$G8_11537_out0 = v$CINA_8606_out0 && v$P$AB_2143_out0;
assign v$G8_11550_out0 = v$CINA_8619_out0 && v$P$AB_2156_out0;
assign {v$A4A_13154_out1,v$A4A_13154_out0 } = v$A3_14607_out0 + v$B3_9471_out0 + v$C2_2686_out0;
assign {v$A4A_13157_out1,v$A4A_13157_out0 } = v$A3_14610_out0 + v$B3_9474_out0 + v$C2_2689_out0;
assign v$IN_15606_out0 = v$IN_5164_out0;
assign v$IN_15608_out0 = v$IN_5174_out0;
assign v$NOT$USED_15950_out0 = v$A2_10044_out1;
assign v$NOT$USED_15951_out0 = v$A2_10045_out1;
assign v$_16096_out0 = { v$SUM$4_15246_out0,v$_8260_out0 };
assign v$G$AD_17086_out0 = v$G4_11111_out0;
assign v$G$AD_17091_out0 = v$G4_11116_out0;
assign v$G$AD_17097_out0 = v$G4_11122_out0;
assign v$G$AD_17100_out0 = v$G4_11125_out0;
assign v$G$AD_17105_out0 = v$G4_11130_out0;
assign v$G$AD_17118_out0 = v$G4_11143_out0;
assign v$G$AD_17209_out0 = v$G4_11234_out0;
assign v$G$AD_17214_out0 = v$G4_11239_out0;
assign v$G$AD_17220_out0 = v$G4_11245_out0;
assign v$G$AD_17223_out0 = v$G4_11248_out0;
assign v$G$AD_17228_out0 = v$G4_11253_out0;
assign v$G$AD_17241_out0 = v$G4_11266_out0;
assign v$C2_18179_out0 = v$C2_2686_out0;
assign v$C2_18182_out0 = v$C2_2689_out0;
assign v$G$CD_917_out0 = v$G$AD_17105_out0;
assign v$G$CD_943_out0 = v$G$AD_17086_out0;
assign v$G$CD_951_out0 = v$G$AD_17100_out0;
assign v$G$CD_1040_out0 = v$G$AD_17228_out0;
assign v$G$CD_1066_out0 = v$G$AD_17209_out0;
assign v$G$CD_1074_out0 = v$G$AD_17223_out0;
assign v$END10_1151_out0 = v$G$AD_17097_out0;
assign v$END10_1154_out0 = v$G$AD_17220_out0;
assign v$P$AB_2004_out0 = v$P$AD_716_out0;
assign v$P$AB_2013_out0 = v$P$AD_716_out0;
assign v$P$AB_2014_out0 = v$P$AD_693_out0;
assign v$P$AB_2025_out0 = v$P$AD_716_out0;
assign v$P$AB_2027_out0 = v$P$AD_716_out0;
assign v$P$AB_2034_out0 = v$P$AD_716_out0;
assign v$P$AB_2035_out0 = v$P$AD_693_out0;
assign v$P$AB_2127_out0 = v$P$AD_839_out0;
assign v$P$AB_2136_out0 = v$P$AD_839_out0;
assign v$P$AB_2137_out0 = v$P$AD_816_out0;
assign v$P$AB_2148_out0 = v$P$AD_839_out0;
assign v$P$AB_2150_out0 = v$P$AD_839_out0;
assign v$P$AB_2157_out0 = v$P$AD_839_out0;
assign v$P$AB_2158_out0 = v$P$AD_816_out0;
assign v$END15_7382_out0 = v$P$AD_697_out0;
assign v$END15_7385_out0 = v$P$AD_820_out0;
assign v$END17_7637_out0 = v$P$AD_726_out0;
assign v$END17_7640_out0 = v$P$AD_849_out0;
assign v$END3_7932_out0 = v$A4A_13154_out1;
assign v$END3_7935_out0 = v$A4A_13157_out1;
assign v$SEL1_8712_out0 = v$IN_15606_out0[23:4];
assign v$SEL1_8722_out0 = v$IN_15608_out0[23:4];
assign v$G$AB_9142_out0 = v$G$AD_17118_out0;
assign v$G$AB_9146_out0 = v$G$AD_17118_out0;
assign v$G$AB_9165_out0 = v$G$AD_17118_out0;
assign v$G$AB_9173_out0 = v$G$AD_17105_out0;
assign v$G$AB_9175_out0 = v$G$AD_17118_out0;
assign v$G$AB_9265_out0 = v$G$AD_17241_out0;
assign v$G$AB_9269_out0 = v$G$AD_17241_out0;
assign v$G$AB_9288_out0 = v$G$AD_17241_out0;
assign v$G$AB_9296_out0 = v$G$AD_17228_out0;
assign v$G$AB_9298_out0 = v$G$AD_17241_out0;
assign v$G7_9635_out0 = v$G8_11395_out0 && v$P$CD_10454_out0;
assign v$G7_9640_out0 = v$G8_11400_out0 && v$P$CD_10459_out0;
assign v$G7_9646_out0 = v$G8_11406_out0 && v$P$CD_10465_out0;
assign v$G7_9649_out0 = v$G8_11409_out0 && v$P$CD_10468_out0;
assign v$G7_9654_out0 = v$G8_11414_out0 && v$P$CD_10473_out0;
assign v$G7_9667_out0 = v$G8_11427_out0 && v$P$CD_10486_out0;
assign v$G7_9758_out0 = v$G8_11518_out0 && v$P$CD_10577_out0;
assign v$G7_9763_out0 = v$G8_11523_out0 && v$P$CD_10582_out0;
assign v$G7_9769_out0 = v$G8_11529_out0 && v$P$CD_10588_out0;
assign v$G7_9772_out0 = v$G8_11532_out0 && v$P$CD_10591_out0;
assign v$G7_9777_out0 = v$G8_11537_out0 && v$P$CD_10596_out0;
assign v$G7_9790_out0 = v$G8_11550_out0 && v$P$CD_10609_out0;
assign v$P$CD_10480_out0 = v$P$AD_724_out0;
assign v$P$CD_10603_out0 = v$P$AD_847_out0;
assign v$END12_10780_out0 = v$G$AD_17091_out0;
assign v$END12_10783_out0 = v$G$AD_17214_out0;
assign v$IN_11073_out0 = v$MULTIPLIER$OUT_9344_out0;
assign v$IN_11074_out0 = v$MULTIPLIER$OUT_9344_out0;
assign v$END19_11655_out0 = v$P$AD_693_out0;
assign v$END19_11658_out0 = v$P$AD_816_out0;
assign v$_12992_out0 = { v$SUM$3_7904_out0,v$_16096_out0 };
assign v$SEL1_15403_out0 = v$IN_15606_out0[19:0];
assign v$SEL1_15413_out0 = v$IN_15608_out0[19:0];
assign v$_18664_out0 = { v$A3A_11951_out0,v$A4A_13154_out0 };
assign v$_18667_out0 = { v$A3A_11954_out0,v$A4A_13157_out0 };
assign v$G6_433_out0 = v$G4_11111_out0 || v$G7_9635_out0;
assign v$G6_438_out0 = v$G4_11116_out0 || v$G7_9640_out0;
assign v$G6_444_out0 = v$G4_11122_out0 || v$G7_9646_out0;
assign v$G6_447_out0 = v$G4_11125_out0 || v$G7_9649_out0;
assign v$G6_452_out0 = v$G4_11130_out0 || v$G7_9654_out0;
assign v$G6_465_out0 = v$G4_11143_out0 || v$G7_9667_out0;
assign v$G6_556_out0 = v$G4_11234_out0 || v$G7_9758_out0;
assign v$G6_561_out0 = v$G4_11239_out0 || v$G7_9763_out0;
assign v$G6_567_out0 = v$G4_11245_out0 || v$G7_9769_out0;
assign v$G6_570_out0 = v$G4_11248_out0 || v$G7_9772_out0;
assign v$G6_575_out0 = v$G4_11253_out0 || v$G7_9777_out0;
assign v$G6_588_out0 = v$G4_11266_out0 || v$G7_9790_out0;
assign v$_4262_out0 = { v$C2_120_out0,v$SEL1_15403_out0 };
assign v$_4272_out0 = { v$C2_130_out0,v$SEL1_15413_out0 };
assign v$G5_4525_out0 = v$G$AB_9142_out0 && v$P$CD_10460_out0;
assign v$G5_4529_out0 = v$G$AB_9146_out0 && v$P$CD_10464_out0;
assign v$G5_4548_out0 = v$G$AB_9165_out0 && v$P$CD_10483_out0;
assign v$G5_4556_out0 = v$G$AB_9173_out0 && v$P$CD_10491_out0;
assign v$G5_4558_out0 = v$G$AB_9175_out0 && v$P$CD_10493_out0;
assign v$G5_4648_out0 = v$G$AB_9265_out0 && v$P$CD_10583_out0;
assign v$G5_4652_out0 = v$G$AB_9269_out0 && v$P$CD_10587_out0;
assign v$G5_4671_out0 = v$G$AB_9288_out0 && v$P$CD_10606_out0;
assign v$G5_4679_out0 = v$G$AB_9296_out0 && v$P$CD_10614_out0;
assign v$G5_4681_out0 = v$G$AB_9298_out0 && v$P$CD_10616_out0;
assign v$G1_5525_out0 = v$P$AB_2004_out0 && v$P$CD_10457_out0;
assign v$G1_5534_out0 = v$P$AB_2013_out0 && v$P$CD_10466_out0;
assign v$G1_5535_out0 = v$P$AB_2014_out0 && v$P$CD_10467_out0;
assign v$G1_5546_out0 = v$P$AB_2025_out0 && v$P$CD_10478_out0;
assign v$G1_5548_out0 = v$P$AB_2027_out0 && v$P$CD_10480_out0;
assign v$G1_5555_out0 = v$P$AB_2034_out0 && v$P$CD_10487_out0;
assign v$G1_5556_out0 = v$P$AB_2035_out0 && v$P$CD_10488_out0;
assign v$G1_5648_out0 = v$P$AB_2127_out0 && v$P$CD_10580_out0;
assign v$G1_5657_out0 = v$P$AB_2136_out0 && v$P$CD_10589_out0;
assign v$G1_5658_out0 = v$P$AB_2137_out0 && v$P$CD_10590_out0;
assign v$G1_5669_out0 = v$P$AB_2148_out0 && v$P$CD_10601_out0;
assign v$G1_5671_out0 = v$P$AB_2150_out0 && v$P$CD_10603_out0;
assign v$G1_5678_out0 = v$P$AB_2157_out0 && v$P$CD_10610_out0;
assign v$G1_5679_out0 = v$P$AB_2158_out0 && v$P$CD_10611_out0;
assign v$_8997_out0 = { v$SEL1_8712_out0,v$C1_5978_out0 };
assign v$_9007_out0 = { v$SEL1_8722_out0,v$C1_5988_out0 };
assign v$_10355_out0 = { v$_13437_out0,v$_18664_out0 };
assign v$_10358_out0 = { v$_13440_out0,v$_18667_out0 };
assign v$IN_11644_out0 = v$IN_11073_out0;
assign v$IN_11645_out0 = v$IN_11074_out0;
assign v$_15860_out0 = { v$SUM$2_9082_out0,v$_12992_out0 };
assign v$P$AD_690_out0 = v$G1_5525_out0;
assign v$P$AD_699_out0 = v$G1_5534_out0;
assign v$P$AD_700_out0 = v$G1_5535_out0;
assign v$P$AD_711_out0 = v$G1_5546_out0;
assign v$P$AD_713_out0 = v$G1_5548_out0;
assign v$P$AD_720_out0 = v$G1_5555_out0;
assign v$P$AD_721_out0 = v$G1_5556_out0;
assign v$P$AD_813_out0 = v$G1_5648_out0;
assign v$P$AD_822_out0 = v$G1_5657_out0;
assign v$P$AD_823_out0 = v$G1_5658_out0;
assign v$P$AD_834_out0 = v$G1_5669_out0;
assign v$P$AD_836_out0 = v$G1_5671_out0;
assign v$P$AD_843_out0 = v$G1_5678_out0;
assign v$P$AD_844_out0 = v$G1_5679_out0;
assign v$_1828_out0 = { v$SUM$1_10360_out0,v$_15860_out0 };
assign v$MUX1_2366_out0 = v$LEFT$SHIT_3058_out0 ? v$_4262_out0 : v$_8997_out0;
assign v$MUX1_2376_out0 = v$LEFT$SHIT_3068_out0 ? v$_4272_out0 : v$_9007_out0;
assign v$COUTD_6693_out0 = v$G6_433_out0;
assign v$COUTD_6698_out0 = v$G6_438_out0;
assign v$COUTD_6704_out0 = v$G6_444_out0;
assign v$COUTD_6707_out0 = v$G6_447_out0;
assign v$COUTD_6712_out0 = v$G6_452_out0;
assign v$COUTD_6725_out0 = v$G6_465_out0;
assign v$COUTD_6816_out0 = v$G6_556_out0;
assign v$COUTD_6821_out0 = v$G6_561_out0;
assign v$COUTD_6827_out0 = v$G6_567_out0;
assign v$COUTD_6830_out0 = v$G6_570_out0;
assign v$COUTD_6835_out0 = v$G6_575_out0;
assign v$COUTD_6848_out0 = v$G6_588_out0;
assign v$IN_8296_out0 = v$IN_11644_out0;
assign v$IN_8297_out0 = v$IN_11645_out0;
assign v$G4_11117_out0 = v$G5_4525_out0 || v$G$CD_920_out0;
assign v$G4_11121_out0 = v$G5_4529_out0 || v$G$CD_924_out0;
assign v$G4_11140_out0 = v$G5_4548_out0 || v$G$CD_943_out0;
assign v$G4_11148_out0 = v$G5_4556_out0 || v$G$CD_951_out0;
assign v$G4_11150_out0 = v$G5_4558_out0 || v$G$CD_953_out0;
assign v$G4_11240_out0 = v$G5_4648_out0 || v$G$CD_1043_out0;
assign v$G4_11244_out0 = v$G5_4652_out0 || v$G$CD_1047_out0;
assign v$G4_11263_out0 = v$G5_4671_out0 || v$G$CD_1066_out0;
assign v$G4_11271_out0 = v$G5_4679_out0 || v$G$CD_1074_out0;
assign v$G4_11273_out0 = v$G5_4681_out0 || v$G$CD_1076_out0;
assign v$IN_13566_out0 = v$IN_11644_out0;
assign v$IN_13570_out0 = v$IN_11645_out0;
assign v$IN_18264_out0 = v$IN_11644_out0;
assign v$IN_18265_out0 = v$IN_11645_out0;
assign v$C4_1259_out0 = v$COUTD_6698_out0;
assign v$C4_1262_out0 = v$COUTD_6821_out0;
assign v$_1606_out0 = { v$SUM$0_12330_out0,v$_1828_out0 };
assign v$P$AB_2017_out0 = v$P$AD_690_out0;
assign v$P$AB_2024_out0 = v$P$AD_690_out0;
assign v$P$AB_2028_out0 = v$P$AD_711_out0;
assign v$P$AB_2031_out0 = v$P$AD_711_out0;
assign v$P$AB_2039_out0 = v$P$AD_690_out0;
assign v$P$AB_2140_out0 = v$P$AD_813_out0;
assign v$P$AB_2147_out0 = v$P$AD_813_out0;
assign v$P$AB_2151_out0 = v$P$AD_834_out0;
assign v$P$AB_2154_out0 = v$P$AD_834_out0;
assign v$P$AB_2162_out0 = v$P$AD_813_out0;
assign v$END27_2210_out0 = v$P$AD_720_out0;
assign v$END27_2213_out0 = v$P$AD_843_out0;
assign v$IN_4192_out0 = v$IN_8296_out0;
assign v$IN_4193_out0 = v$IN_8297_out0;
assign v$END21_4340_out0 = v$P$AD_700_out0;
assign v$END21_4343_out0 = v$P$AD_823_out0;
assign v$IN_5187_out0 = v$IN_18264_out0;
assign v$IN_5193_out0 = v$IN_18265_out0;
assign v$END40_5775_out0 = v$COUTD_6712_out0;
assign v$END40_5778_out0 = v$COUTD_6835_out0;
assign v$END29_5885_out0 = v$P$AD_711_out0;
assign v$END29_5888_out0 = v$P$AD_834_out0;
assign v$SEL3_7366_out0 = v$IN_13566_out0[47:32];
assign v$SEL3_7370_out0 = v$IN_13570_out0[47:32];
assign v$CINA_8470_out0 = v$COUTD_6725_out0;
assign v$CINA_8474_out0 = v$COUTD_6725_out0;
assign v$CINA_8493_out0 = v$COUTD_6725_out0;
assign v$CINA_8501_out0 = v$COUTD_6712_out0;
assign v$CINA_8503_out0 = v$COUTD_6725_out0;
assign v$CINA_8593_out0 = v$COUTD_6848_out0;
assign v$CINA_8597_out0 = v$COUTD_6848_out0;
assign v$CINA_8616_out0 = v$COUTD_6848_out0;
assign v$CINA_8624_out0 = v$COUTD_6835_out0;
assign v$CINA_8626_out0 = v$COUTD_6848_out0;
assign v$END4_9367_out0 = v$COUTD_6693_out0;
assign v$END4_9370_out0 = v$COUTD_6816_out0;
assign v$END52_11973_out0 = v$P$AD_713_out0;
assign v$END52_11976_out0 = v$P$AD_836_out0;
assign v$SEL2_13852_out0 = v$IN_13566_out0[31:16];
assign v$SEL2_13856_out0 = v$IN_13570_out0[31:16];
assign v$END60_15132_out0 = v$COUTD_6707_out0;
assign v$END60_15135_out0 = v$COUTD_6830_out0;
assign v$MUX2_15237_out0 = v$EN_4754_out0 ? v$MUX1_2366_out0 : v$IN_15606_out0;
assign v$MUX2_15239_out0 = v$EN_4756_out0 ? v$MUX1_2376_out0 : v$IN_15608_out0;
assign v$C3_15726_out0 = v$COUTD_6704_out0;
assign v$C3_15729_out0 = v$COUTD_6827_out0;
assign v$C5_15915_out0 = v$COUTD_6725_out0;
assign v$C5_15918_out0 = v$COUTD_6848_out0;
assign v$SEL1_16688_out0 = v$IN_13566_out0[15:0];
assign v$SEL1_16692_out0 = v$IN_13570_out0[15:0];
assign v$END23_16717_out0 = v$P$AD_721_out0;
assign v$END23_16720_out0 = v$P$AD_844_out0;
assign v$END25_17070_out0 = v$P$AD_699_out0;
assign v$END25_17073_out0 = v$P$AD_822_out0;
assign v$G$AD_17092_out0 = v$G4_11117_out0;
assign v$G$AD_17096_out0 = v$G4_11121_out0;
assign v$G$AD_17115_out0 = v$G4_11140_out0;
assign v$G$AD_17123_out0 = v$G4_11148_out0;
assign v$G$AD_17125_out0 = v$G4_11150_out0;
assign v$G$AD_17215_out0 = v$G4_11240_out0;
assign v$G$AD_17219_out0 = v$G4_11244_out0;
assign v$G$AD_17238_out0 = v$G4_11263_out0;
assign v$G$AD_17246_out0 = v$G4_11271_out0;
assign v$G$AD_17248_out0 = v$G4_11273_out0;
assign v$END16_216_out0 = v$G$AD_17125_out0;
assign v$END16_219_out0 = v$G$AD_17248_out0;
assign v$END14_274_out0 = v$G$AD_17096_out0;
assign v$END14_277_out0 = v$G$AD_17219_out0;
assign v$G$CD_940_out0 = v$G$AD_17123_out0;
assign v$G$CD_1063_out0 = v$G$AD_17246_out0;
assign {v$A7A_1657_out1,v$A7A_1657_out0 } = v$A5_6665_out0 + v$B5_18374_out0 + v$C4_1259_out0;
assign {v$A7A_1660_out1,v$A7A_1660_out0 } = v$A5_6668_out0 + v$B5_18377_out0 + v$C4_1262_out0;
assign v$C4_1876_out0 = v$C4_1259_out0;
assign v$C4_1879_out0 = v$C4_1262_out0;
assign {v$A6A_3121_out1,v$A6A_3121_out0 } = v$A6_308_out0 + v$B6_13298_out0 + v$C5_15915_out0;
assign {v$A6A_3124_out1,v$A6A_3124_out0 } = v$A6_311_out0 + v$B6_13301_out0 + v$C5_15918_out0;
assign v$IN_3868_out0 = v$IN_5187_out0;
assign v$IN_3871_out0 = v$IN_5193_out0;
assign v$SEL15_4888_out0 = v$IN_4192_out0[33:33];
assign v$SEL15_4889_out0 = v$IN_4193_out0[33:33];
assign v$G1_5538_out0 = v$P$AB_2017_out0 && v$P$CD_10470_out0;
assign v$G1_5545_out0 = v$P$AB_2024_out0 && v$P$CD_10477_out0;
assign v$G1_5549_out0 = v$P$AB_2028_out0 && v$P$CD_10481_out0;
assign v$G1_5552_out0 = v$P$AB_2031_out0 && v$P$CD_10484_out0;
assign v$G1_5560_out0 = v$P$AB_2039_out0 && v$P$CD_10492_out0;
assign v$G1_5661_out0 = v$P$AB_2140_out0 && v$P$CD_10593_out0;
assign v$G1_5668_out0 = v$P$AB_2147_out0 && v$P$CD_10600_out0;
assign v$G1_5672_out0 = v$P$AB_2151_out0 && v$P$CD_10604_out0;
assign v$G1_5675_out0 = v$P$AB_2154_out0 && v$P$CD_10607_out0;
assign v$G1_5683_out0 = v$P$AB_2162_out0 && v$P$CD_10615_out0;
assign v$SEL13_6926_out0 = v$IN_4192_out0[35:35];
assign v$SEL13_6927_out0 = v$IN_4193_out0[35:35];
assign v$SEL1_7090_out0 = v$IN_4192_out0[47:47];
assign v$SEL1_7091_out0 = v$IN_4193_out0[47:47];
assign v$SEL11_7227_out0 = v$IN_4192_out0[37:37];
assign v$SEL11_7228_out0 = v$IN_4193_out0[37:37];
assign v$SEL4_7323_out0 = v$IN_4192_out0[44:44];
assign v$SEL4_7324_out0 = v$IN_4193_out0[44:44];
assign v$SEL22_7399_out0 = v$IN_4192_out0[26:26];
assign v$SEL22_7400_out0 = v$IN_4193_out0[26:26];
assign v$SEL23_7619_out0 = v$IN_4192_out0[25:25];
assign v$SEL23_7620_out0 = v$IN_4193_out0[25:25];
assign v$SEL20_8176_out0 = v$IN_4192_out0[28:28];
assign v$SEL20_8177_out0 = v$IN_4193_out0[28:28];
assign v$G$AB_9139_out0 = v$G$AD_17115_out0;
assign v$G$AB_9148_out0 = v$G$AD_17115_out0;
assign v$G$AB_9149_out0 = v$G$AD_17092_out0;
assign v$G$AB_9160_out0 = v$G$AD_17115_out0;
assign v$G$AB_9162_out0 = v$G$AD_17115_out0;
assign v$G$AB_9169_out0 = v$G$AD_17115_out0;
assign v$G$AB_9170_out0 = v$G$AD_17092_out0;
assign v$G$AB_9262_out0 = v$G$AD_17238_out0;
assign v$G$AB_9271_out0 = v$G$AD_17238_out0;
assign v$G$AB_9272_out0 = v$G$AD_17215_out0;
assign v$G$AB_9283_out0 = v$G$AD_17238_out0;
assign v$G$AB_9285_out0 = v$G$AD_17238_out0;
assign v$G$AB_9292_out0 = v$G$AD_17238_out0;
assign v$G$AB_9293_out0 = v$G$AD_17215_out0;
assign v$SEL10_9508_out0 = v$IN_4192_out0[40:40];
assign v$SEL10_9509_out0 = v$IN_4193_out0[40:40];
assign v$SEL9_10265_out0 = v$IN_4192_out0[38:38];
assign v$SEL9_10266_out0 = v$IN_4193_out0[38:38];
assign v$SEL21_11050_out0 = v$IN_4192_out0[27:27];
assign v$SEL21_11051_out0 = v$IN_4193_out0[27:27];
assign v$SEL18_11381_out0 = v$IN_4192_out0[30:30];
assign v$SEL18_11382_out0 = v$IN_4193_out0[30:30];
assign v$G8_11401_out0 = v$CINA_8470_out0 && v$P$AB_2007_out0;
assign v$G8_11405_out0 = v$CINA_8474_out0 && v$P$AB_2011_out0;
assign v$G8_11424_out0 = v$CINA_8493_out0 && v$P$AB_2030_out0;
assign v$G8_11432_out0 = v$CINA_8501_out0 && v$P$AB_2038_out0;
assign v$G8_11434_out0 = v$CINA_8503_out0 && v$P$AB_2040_out0;
assign v$G8_11524_out0 = v$CINA_8593_out0 && v$P$AB_2130_out0;
assign v$G8_11528_out0 = v$CINA_8597_out0 && v$P$AB_2134_out0;
assign v$G8_11547_out0 = v$CINA_8616_out0 && v$P$AB_2153_out0;
assign v$G8_11555_out0 = v$CINA_8624_out0 && v$P$AB_2161_out0;
assign v$G8_11557_out0 = v$CINA_8626_out0 && v$P$AB_2163_out0;
assign v$C5_11686_out0 = v$C5_15915_out0;
assign v$C5_11689_out0 = v$C5_15918_out0;
assign v$SEL3_11731_out0 = v$IN_4192_out0[45:45];
assign v$SEL3_11732_out0 = v$IN_4193_out0[45:45];
assign v$END18_11946_out0 = v$G$AD_17092_out0;
assign v$END18_11949_out0 = v$G$AD_17215_out0;
assign v$SEL6_12474_out0 = v$IN_4192_out0[42:42];
assign v$SEL6_12475_out0 = v$IN_4193_out0[42:42];
assign v$SEL19_12817_out0 = v$IN_4192_out0[29:29];
assign v$SEL19_12818_out0 = v$IN_4193_out0[29:29];
assign v$SEL2_13323_out0 = v$IN_4192_out0[46:46];
assign v$SEL2_13324_out0 = v$IN_4193_out0[46:46];
assign v$IN_13567_out0 = v$SEL1_16688_out0;
assign v$IN_13568_out0 = v$SEL2_13852_out0;
assign v$IN_13569_out0 = v$SEL3_7366_out0;
assign v$IN_13571_out0 = v$SEL1_16692_out0;
assign v$IN_13572_out0 = v$SEL2_13856_out0;
assign v$IN_13573_out0 = v$SEL3_7370_out0;
assign v$SEL12_13846_out0 = v$IN_4192_out0[36:36];
assign v$SEL12_13847_out0 = v$IN_4193_out0[36:36];
assign v$SEL7_14334_out0 = v$IN_4192_out0[41:41];
assign v$SEL7_14335_out0 = v$IN_4193_out0[41:41];
assign v$OUT_14918_out0 = v$MUX2_15237_out0;
assign v$OUT_14928_out0 = v$MUX2_15239_out0;
assign v$SEL5_15453_out0 = v$IN_4192_out0[43:43];
assign v$SEL5_15454_out0 = v$IN_4193_out0[43:43];
assign v$C3_15817_out0 = v$C3_15726_out0;
assign v$C3_15820_out0 = v$C3_15729_out0;
assign v$SEL17_16071_out0 = v$IN_4192_out0[31:31];
assign v$SEL17_16072_out0 = v$IN_4193_out0[31:31];
assign {v$A5A_16099_out1,v$A5A_16099_out0 } = v$A4_17498_out0 + v$B4_14663_out0 + v$C3_15726_out0;
assign {v$A5A_16102_out1,v$A5A_16102_out0 } = v$A4_17501_out0 + v$B4_14666_out0 + v$C3_15729_out0;
assign v$SEL14_16349_out0 = v$IN_4192_out0[34:34];
assign v$SEL14_16350_out0 = v$IN_4193_out0[34:34];
assign v$SEL16_16896_out0 = v$IN_4192_out0[32:32];
assign v$SEL16_16897_out0 = v$IN_4193_out0[32:32];
assign v$SEL24_16924_out0 = v$IN_4192_out0[24:24];
assign v$SEL24_16925_out0 = v$IN_4193_out0[24:24];
assign v$SEL8_17685_out0 = v$IN_4192_out0[39:39];
assign v$SEL8_17686_out0 = v$IN_4193_out0[39:39];
assign v$_82_out0 = { v$A5A_16099_out0,v$A7A_1657_out0 };
assign v$_85_out0 = { v$A5A_16102_out0,v$A7A_1660_out0 };
assign v$P$AD_703_out0 = v$G1_5538_out0;
assign v$P$AD_710_out0 = v$G1_5545_out0;
assign v$P$AD_714_out0 = v$G1_5549_out0;
assign v$P$AD_717_out0 = v$G1_5552_out0;
assign v$P$AD_725_out0 = v$G1_5560_out0;
assign v$P$AD_826_out0 = v$G1_5661_out0;
assign v$P$AD_833_out0 = v$G1_5668_out0;
assign v$P$AD_837_out0 = v$G1_5672_out0;
assign v$P$AD_840_out0 = v$G1_5675_out0;
assign v$P$AD_848_out0 = v$G1_5683_out0;
assign v$_2453_out0 = { v$C4_1876_out0,v$C5_11686_out0 };
assign v$_2456_out0 = { v$C4_1879_out0,v$C5_11689_out0 };
assign v$SEL4_3370_out0 = v$IN_13567_out0[15:12];
assign v$SEL4_3371_out0 = v$IN_13568_out0[15:12];
assign v$SEL4_3372_out0 = v$IN_13569_out0[15:12];
assign v$SEL4_3373_out0 = v$IN_13571_out0[15:12];
assign v$SEL4_3374_out0 = v$IN_13572_out0[15:12];
assign v$SEL4_3375_out0 = v$IN_13573_out0[15:12];
assign v$END5_4143_out0 = v$A7A_1657_out1;
assign v$END5_4146_out0 = v$A7A_1660_out1;
assign v$G5_4522_out0 = v$G$AB_9139_out0 && v$P$CD_10457_out0;
assign v$G5_4531_out0 = v$G$AB_9148_out0 && v$P$CD_10466_out0;
assign v$G5_4532_out0 = v$G$AB_9149_out0 && v$P$CD_10467_out0;
assign v$G5_4543_out0 = v$G$AB_9160_out0 && v$P$CD_10478_out0;
assign v$G5_4545_out0 = v$G$AB_9162_out0 && v$P$CD_10480_out0;
assign v$G5_4552_out0 = v$G$AB_9169_out0 && v$P$CD_10487_out0;
assign v$G5_4553_out0 = v$G$AB_9170_out0 && v$P$CD_10488_out0;
assign v$G5_4645_out0 = v$G$AB_9262_out0 && v$P$CD_10580_out0;
assign v$G5_4654_out0 = v$G$AB_9271_out0 && v$P$CD_10589_out0;
assign v$G5_4655_out0 = v$G$AB_9272_out0 && v$P$CD_10590_out0;
assign v$G5_4666_out0 = v$G$AB_9283_out0 && v$P$CD_10601_out0;
assign v$G5_4668_out0 = v$G$AB_9285_out0 && v$P$CD_10603_out0;
assign v$G5_4675_out0 = v$G$AB_9292_out0 && v$P$CD_10610_out0;
assign v$G5_4676_out0 = v$G$AB_9293_out0 && v$P$CD_10611_out0;
assign v$IN_5163_out0 = v$OUT_14918_out0;
assign v$IN_5173_out0 = v$OUT_14928_out0;
assign v$END4_5246_out0 = v$A5A_16099_out1;
assign v$END4_5249_out0 = v$A5A_16102_out1;
assign v$SEL3_7367_out0 = v$IN_13567_out0[11:8];
assign v$SEL3_7368_out0 = v$IN_13568_out0[11:8];
assign v$SEL3_7369_out0 = v$IN_13569_out0[11:8];
assign v$SEL3_7371_out0 = v$IN_13571_out0[11:8];
assign v$SEL3_7372_out0 = v$IN_13572_out0[11:8];
assign v$SEL3_7373_out0 = v$IN_13573_out0[11:8];
assign v$SEL1_8735_out0 = v$IN_3868_out0[47:1];
assign v$SEL1_8741_out0 = v$IN_3871_out0[47:1];
assign v$G7_9641_out0 = v$G8_11401_out0 && v$P$CD_10460_out0;
assign v$G7_9645_out0 = v$G8_11405_out0 && v$P$CD_10464_out0;
assign v$G7_9664_out0 = v$G8_11424_out0 && v$P$CD_10483_out0;
assign v$G7_9672_out0 = v$G8_11432_out0 && v$P$CD_10491_out0;
assign v$G7_9674_out0 = v$G8_11434_out0 && v$P$CD_10493_out0;
assign v$G7_9764_out0 = v$G8_11524_out0 && v$P$CD_10583_out0;
assign v$G7_9768_out0 = v$G8_11528_out0 && v$P$CD_10587_out0;
assign v$G7_9787_out0 = v$G8_11547_out0 && v$P$CD_10606_out0;
assign v$G7_9795_out0 = v$G8_11555_out0 && v$P$CD_10614_out0;
assign v$G7_9797_out0 = v$G8_11557_out0 && v$P$CD_10616_out0;
assign v$SEL2_13853_out0 = v$IN_13567_out0[7:4];
assign v$SEL2_13854_out0 = v$IN_13568_out0[7:4];
assign v$SEL2_13855_out0 = v$IN_13569_out0[7:4];
assign v$SEL2_13857_out0 = v$IN_13571_out0[7:4];
assign v$SEL2_13858_out0 = v$IN_13572_out0[7:4];
assign v$SEL2_13859_out0 = v$IN_13573_out0[7:4];
assign v$_14998_out0 = { v$C2_18179_out0,v$C3_15817_out0 };
assign v$_15001_out0 = { v$C2_18182_out0,v$C3_15820_out0 };
assign v$END6_15249_out0 = v$A6A_3121_out1;
assign v$END6_15252_out0 = v$A6A_3124_out1;
assign v$SEL1_15426_out0 = v$IN_3868_out0[46:0];
assign v$SEL1_15432_out0 = v$IN_3871_out0[46:0];
assign v$SEL1_16689_out0 = v$IN_13567_out0[3:0];
assign v$SEL1_16690_out0 = v$IN_13568_out0[3:0];
assign v$SEL1_16691_out0 = v$IN_13569_out0[3:0];
assign v$SEL1_16693_out0 = v$IN_13571_out0[3:0];
assign v$SEL1_16694_out0 = v$IN_13572_out0[3:0];
assign v$SEL1_16695_out0 = v$IN_13573_out0[3:0];
assign v$MUX24_18058_out0 = v$EQ24_2538_out0 ? v$SEL24_16924_out0 : v$C1_15722_out0;
assign v$MUX24_18059_out0 = v$EQ24_2539_out0 ? v$SEL24_16925_out0 : v$C1_15723_out0;
assign v$END33_264_out0 = v$P$AD_717_out0;
assign v$END33_267_out0 = v$P$AD_840_out0;
assign v$G6_439_out0 = v$G4_11117_out0 || v$G7_9641_out0;
assign v$G6_443_out0 = v$G4_11121_out0 || v$G7_9645_out0;
assign v$G6_462_out0 = v$G4_11140_out0 || v$G7_9664_out0;
assign v$G6_470_out0 = v$G4_11148_out0 || v$G7_9672_out0;
assign v$G6_472_out0 = v$G4_11150_out0 || v$G7_9674_out0;
assign v$G6_562_out0 = v$G4_11240_out0 || v$G7_9764_out0;
assign v$G6_566_out0 = v$G4_11244_out0 || v$G7_9768_out0;
assign v$G6_585_out0 = v$G4_11263_out0 || v$G7_9787_out0;
assign v$G6_593_out0 = v$G4_11271_out0 || v$G7_9795_out0;
assign v$G6_595_out0 = v$G4_11273_out0 || v$G7_9797_out0;
assign v$P$AB_2010_out0 = v$P$AD_710_out0;
assign v$P$AB_2029_out0 = v$P$AD_710_out0;
assign v$P$AB_2133_out0 = v$P$AD_833_out0;
assign v$P$AB_2152_out0 = v$P$AD_833_out0;
assign v$END47_2679_out0 = v$P$AD_710_out0;
assign v$END47_2682_out0 = v$P$AD_833_out0;
assign v$_4285_out0 = { v$C2_143_out0,v$SEL1_15426_out0 };
assign v$_4291_out0 = { v$C2_149_out0,v$SEL1_15432_out0 };
assign v$IN_5024_out0 = v$IN_5163_out0;
assign v$IN_5027_out0 = v$IN_5173_out0;
assign v$_7253_out0 = { v$_8906_out0,v$_14998_out0 };
assign v$_7256_out0 = { v$_8909_out0,v$_15001_out0 };
assign v$_9020_out0 = { v$SEL1_8735_out0,v$C1_6001_out0 };
assign v$_9026_out0 = { v$SEL1_8741_out0,v$C1_6007_out0 };
assign v$G4_11114_out0 = v$G5_4522_out0 || v$G$CD_917_out0;
assign v$G4_11123_out0 = v$G5_4531_out0 || v$G$CD_926_out0;
assign v$G4_11124_out0 = v$G5_4532_out0 || v$G$CD_927_out0;
assign v$G4_11135_out0 = v$G5_4543_out0 || v$G$CD_938_out0;
assign v$G4_11137_out0 = v$G5_4545_out0 || v$G$CD_940_out0;
assign v$G4_11144_out0 = v$G5_4552_out0 || v$G$CD_947_out0;
assign v$G4_11145_out0 = v$G5_4553_out0 || v$G$CD_948_out0;
assign v$G4_11237_out0 = v$G5_4645_out0 || v$G$CD_1040_out0;
assign v$G4_11246_out0 = v$G5_4654_out0 || v$G$CD_1049_out0;
assign v$G4_11247_out0 = v$G5_4655_out0 || v$G$CD_1050_out0;
assign v$G4_11258_out0 = v$G5_4666_out0 || v$G$CD_1061_out0;
assign v$G4_11260_out0 = v$G5_4668_out0 || v$G$CD_1063_out0;
assign v$G4_11267_out0 = v$G5_4675_out0 || v$G$CD_1070_out0;
assign v$G4_11268_out0 = v$G5_4676_out0 || v$G$CD_1071_out0;
assign v$IN_15075_out0 = v$SEL3_7367_out0;
assign v$IN_15076_out0 = v$SEL1_16689_out0;
assign v$IN_15077_out0 = v$SEL2_13853_out0;
assign v$IN_15078_out0 = v$SEL4_3370_out0;
assign v$IN_15079_out0 = v$SEL3_7368_out0;
assign v$IN_15080_out0 = v$SEL1_16690_out0;
assign v$IN_15081_out0 = v$SEL2_13854_out0;
assign v$IN_15082_out0 = v$SEL4_3371_out0;
assign v$IN_15083_out0 = v$SEL3_7369_out0;
assign v$IN_15084_out0 = v$SEL1_16691_out0;
assign v$IN_15085_out0 = v$SEL2_13855_out0;
assign v$IN_15086_out0 = v$SEL4_3372_out0;
assign v$IN_15087_out0 = v$SEL3_7371_out0;
assign v$IN_15088_out0 = v$SEL1_16693_out0;
assign v$IN_15089_out0 = v$SEL2_13857_out0;
assign v$IN_15090_out0 = v$SEL4_3373_out0;
assign v$IN_15091_out0 = v$SEL3_7372_out0;
assign v$IN_15092_out0 = v$SEL1_16694_out0;
assign v$IN_15093_out0 = v$SEL2_13858_out0;
assign v$IN_15094_out0 = v$SEL4_3374_out0;
assign v$IN_15095_out0 = v$SEL3_7373_out0;
assign v$IN_15096_out0 = v$SEL1_16695_out0;
assign v$IN_15097_out0 = v$SEL2_13859_out0;
assign v$IN_15098_out0 = v$SEL4_3375_out0;
assign v$END44_15665_out0 = v$P$AD_725_out0;
assign v$END44_15668_out0 = v$P$AD_848_out0;
assign v$MUX23_16225_out0 = v$EQ23_3196_out0 ? v$SEL23_7619_out0 : v$MUX24_18058_out0;
assign v$MUX23_16226_out0 = v$EQ23_3197_out0 ? v$SEL23_7620_out0 : v$MUX24_18059_out0;
assign v$END42_18311_out0 = v$P$AD_703_out0;
assign v$END42_18314_out0 = v$P$AD_826_out0;
assign v$END31_18520_out0 = v$P$AD_714_out0;
assign v$END31_18523_out0 = v$P$AD_837_out0;
assign v$SEL3_2312_out0 = v$IN_15075_out0[2:2];
assign v$SEL3_2313_out0 = v$IN_15076_out0[2:2];
assign v$SEL3_2314_out0 = v$IN_15077_out0[2:2];
assign v$SEL3_2315_out0 = v$IN_15078_out0[2:2];
assign v$SEL3_2316_out0 = v$IN_15079_out0[2:2];
assign v$SEL3_2317_out0 = v$IN_15080_out0[2:2];
assign v$SEL3_2318_out0 = v$IN_15081_out0[2:2];
assign v$SEL3_2319_out0 = v$IN_15082_out0[2:2];
assign v$SEL3_2320_out0 = v$IN_15083_out0[2:2];
assign v$SEL3_2321_out0 = v$IN_15084_out0[2:2];
assign v$SEL3_2322_out0 = v$IN_15085_out0[2:2];
assign v$SEL3_2323_out0 = v$IN_15086_out0[2:2];
assign v$SEL3_2324_out0 = v$IN_15087_out0[2:2];
assign v$SEL3_2325_out0 = v$IN_15088_out0[2:2];
assign v$SEL3_2326_out0 = v$IN_15089_out0[2:2];
assign v$SEL3_2327_out0 = v$IN_15090_out0[2:2];
assign v$SEL3_2328_out0 = v$IN_15091_out0[2:2];
assign v$SEL3_2329_out0 = v$IN_15092_out0[2:2];
assign v$SEL3_2330_out0 = v$IN_15093_out0[2:2];
assign v$SEL3_2331_out0 = v$IN_15094_out0[2:2];
assign v$SEL3_2332_out0 = v$IN_15095_out0[2:2];
assign v$SEL3_2333_out0 = v$IN_15096_out0[2:2];
assign v$SEL3_2334_out0 = v$IN_15097_out0[2:2];
assign v$SEL3_2335_out0 = v$IN_15098_out0[2:2];
assign v$MUX1_2389_out0 = v$LEFT$SHIT_3081_out0 ? v$_4285_out0 : v$_9020_out0;
assign v$MUX1_2395_out0 = v$LEFT$SHIT_3087_out0 ? v$_4291_out0 : v$_9026_out0;
assign v$G1_5531_out0 = v$P$AB_2010_out0 && v$P$CD_10463_out0;
assign v$G1_5550_out0 = v$P$AB_2029_out0 && v$P$CD_10482_out0;
assign v$G1_5654_out0 = v$P$AB_2133_out0 && v$P$CD_10586_out0;
assign v$G1_5673_out0 = v$P$AB_2152_out0 && v$P$CD_10605_out0;
assign v$SEL4_6097_out0 = v$IN_15075_out0[3:3];
assign v$SEL4_6098_out0 = v$IN_15076_out0[3:3];
assign v$SEL4_6099_out0 = v$IN_15077_out0[3:3];
assign v$SEL4_6100_out0 = v$IN_15078_out0[3:3];
assign v$SEL4_6101_out0 = v$IN_15079_out0[3:3];
assign v$SEL4_6102_out0 = v$IN_15080_out0[3:3];
assign v$SEL4_6103_out0 = v$IN_15081_out0[3:3];
assign v$SEL4_6104_out0 = v$IN_15082_out0[3:3];
assign v$SEL4_6105_out0 = v$IN_15083_out0[3:3];
assign v$SEL4_6106_out0 = v$IN_15084_out0[3:3];
assign v$SEL4_6107_out0 = v$IN_15085_out0[3:3];
assign v$SEL4_6108_out0 = v$IN_15086_out0[3:3];
assign v$SEL4_6109_out0 = v$IN_15087_out0[3:3];
assign v$SEL4_6110_out0 = v$IN_15088_out0[3:3];
assign v$SEL4_6111_out0 = v$IN_15089_out0[3:3];
assign v$SEL4_6112_out0 = v$IN_15090_out0[3:3];
assign v$SEL4_6113_out0 = v$IN_15091_out0[3:3];
assign v$SEL4_6114_out0 = v$IN_15092_out0[3:3];
assign v$SEL4_6115_out0 = v$IN_15093_out0[3:3];
assign v$SEL4_6116_out0 = v$IN_15094_out0[3:3];
assign v$SEL4_6117_out0 = v$IN_15095_out0[3:3];
assign v$SEL4_6118_out0 = v$IN_15096_out0[3:3];
assign v$SEL4_6119_out0 = v$IN_15097_out0[3:3];
assign v$SEL4_6120_out0 = v$IN_15098_out0[3:3];
assign v$COUTD_6699_out0 = v$G6_439_out0;
assign v$COUTD_6703_out0 = v$G6_443_out0;
assign v$COUTD_6722_out0 = v$G6_462_out0;
assign v$COUTD_6730_out0 = v$G6_470_out0;
assign v$COUTD_6732_out0 = v$G6_472_out0;
assign v$COUTD_6822_out0 = v$G6_562_out0;
assign v$COUTD_6826_out0 = v$G6_566_out0;
assign v$COUTD_6845_out0 = v$G6_585_out0;
assign v$COUTD_6853_out0 = v$G6_593_out0;
assign v$COUTD_6855_out0 = v$G6_595_out0;
assign v$SEL2_7688_out0 = v$IN_15075_out0[1:1];
assign v$SEL2_7689_out0 = v$IN_15076_out0[1:1];
assign v$SEL2_7690_out0 = v$IN_15077_out0[1:1];
assign v$SEL2_7691_out0 = v$IN_15078_out0[1:1];
assign v$SEL2_7692_out0 = v$IN_15079_out0[1:1];
assign v$SEL2_7693_out0 = v$IN_15080_out0[1:1];
assign v$SEL2_7694_out0 = v$IN_15081_out0[1:1];
assign v$SEL2_7695_out0 = v$IN_15082_out0[1:1];
assign v$SEL2_7696_out0 = v$IN_15083_out0[1:1];
assign v$SEL2_7697_out0 = v$IN_15084_out0[1:1];
assign v$SEL2_7698_out0 = v$IN_15085_out0[1:1];
assign v$SEL2_7699_out0 = v$IN_15086_out0[1:1];
assign v$SEL2_7700_out0 = v$IN_15087_out0[1:1];
assign v$SEL2_7701_out0 = v$IN_15088_out0[1:1];
assign v$SEL2_7702_out0 = v$IN_15089_out0[1:1];
assign v$SEL2_7703_out0 = v$IN_15090_out0[1:1];
assign v$SEL2_7704_out0 = v$IN_15091_out0[1:1];
assign v$SEL2_7705_out0 = v$IN_15092_out0[1:1];
assign v$SEL2_7706_out0 = v$IN_15093_out0[1:1];
assign v$SEL2_7707_out0 = v$IN_15094_out0[1:1];
assign v$SEL2_7708_out0 = v$IN_15095_out0[1:1];
assign v$SEL2_7709_out0 = v$IN_15096_out0[1:1];
assign v$SEL2_7710_out0 = v$IN_15097_out0[1:1];
assign v$SEL2_7711_out0 = v$IN_15098_out0[1:1];
assign v$SEL1_8711_out0 = v$IN_5024_out0[23:8];
assign v$SEL1_8721_out0 = v$IN_5027_out0[23:8];
assign v$SEL1_13477_out0 = v$IN_15075_out0[0:0];
assign v$SEL1_13478_out0 = v$IN_15076_out0[0:0];
assign v$SEL1_13479_out0 = v$IN_15077_out0[0:0];
assign v$SEL1_13480_out0 = v$IN_15078_out0[0:0];
assign v$SEL1_13481_out0 = v$IN_15079_out0[0:0];
assign v$SEL1_13482_out0 = v$IN_15080_out0[0:0];
assign v$SEL1_13483_out0 = v$IN_15081_out0[0:0];
assign v$SEL1_13484_out0 = v$IN_15082_out0[0:0];
assign v$SEL1_13485_out0 = v$IN_15083_out0[0:0];
assign v$SEL1_13486_out0 = v$IN_15084_out0[0:0];
assign v$SEL1_13487_out0 = v$IN_15085_out0[0:0];
assign v$SEL1_13488_out0 = v$IN_15086_out0[0:0];
assign v$SEL1_13489_out0 = v$IN_15087_out0[0:0];
assign v$SEL1_13490_out0 = v$IN_15088_out0[0:0];
assign v$SEL1_13491_out0 = v$IN_15089_out0[0:0];
assign v$SEL1_13492_out0 = v$IN_15090_out0[0:0];
assign v$SEL1_13493_out0 = v$IN_15091_out0[0:0];
assign v$SEL1_13494_out0 = v$IN_15092_out0[0:0];
assign v$SEL1_13495_out0 = v$IN_15093_out0[0:0];
assign v$SEL1_13496_out0 = v$IN_15094_out0[0:0];
assign v$SEL1_13497_out0 = v$IN_15095_out0[0:0];
assign v$SEL1_13498_out0 = v$IN_15096_out0[0:0];
assign v$SEL1_13499_out0 = v$IN_15097_out0[0:0];
assign v$SEL1_13500_out0 = v$IN_15098_out0[0:0];
assign v$SEL1_15402_out0 = v$IN_5024_out0[15:0];
assign v$SEL1_15412_out0 = v$IN_5027_out0[15:0];
assign v$MUX22_16466_out0 = v$EQ22_2838_out0 ? v$SEL22_7399_out0 : v$MUX23_16225_out0;
assign v$MUX22_16467_out0 = v$EQ22_2839_out0 ? v$SEL22_7400_out0 : v$MUX23_16226_out0;
assign v$G$AD_17089_out0 = v$G4_11114_out0;
assign v$G$AD_17098_out0 = v$G4_11123_out0;
assign v$G$AD_17099_out0 = v$G4_11124_out0;
assign v$G$AD_17110_out0 = v$G4_11135_out0;
assign v$G$AD_17112_out0 = v$G4_11137_out0;
assign v$G$AD_17119_out0 = v$G4_11144_out0;
assign v$G$AD_17120_out0 = v$G4_11145_out0;
assign v$G$AD_17212_out0 = v$G4_11237_out0;
assign v$G$AD_17221_out0 = v$G4_11246_out0;
assign v$G$AD_17222_out0 = v$G4_11247_out0;
assign v$G$AD_17233_out0 = v$G4_11258_out0;
assign v$G$AD_17235_out0 = v$G4_11260_out0;
assign v$G$AD_17242_out0 = v$G4_11267_out0;
assign v$G$AD_17243_out0 = v$G4_11268_out0;
assign v$END53_317_out0 = v$G$AD_17112_out0;
assign v$END53_320_out0 = v$G$AD_17235_out0;
assign v$P$AD_696_out0 = v$G1_5531_out0;
assign v$P$AD_715_out0 = v$G1_5550_out0;
assign v$P$AD_819_out0 = v$G1_5654_out0;
assign v$P$AD_838_out0 = v$G1_5673_out0;
assign v$G10_1398_out0 = !(v$SEL1_13477_out0 || v$SEL2_7688_out0);
assign v$G10_1399_out0 = !(v$SEL1_13478_out0 || v$SEL2_7689_out0);
assign v$G10_1400_out0 = !(v$SEL1_13479_out0 || v$SEL2_7690_out0);
assign v$G10_1401_out0 = !(v$SEL1_13480_out0 || v$SEL2_7691_out0);
assign v$G10_1402_out0 = !(v$SEL1_13481_out0 || v$SEL2_7692_out0);
assign v$G10_1403_out0 = !(v$SEL1_13482_out0 || v$SEL2_7693_out0);
assign v$G10_1404_out0 = !(v$SEL1_13483_out0 || v$SEL2_7694_out0);
assign v$G10_1405_out0 = !(v$SEL1_13484_out0 || v$SEL2_7695_out0);
assign v$G10_1406_out0 = !(v$SEL1_13485_out0 || v$SEL2_7696_out0);
assign v$G10_1407_out0 = !(v$SEL1_13486_out0 || v$SEL2_7697_out0);
assign v$G10_1408_out0 = !(v$SEL1_13487_out0 || v$SEL2_7698_out0);
assign v$G10_1409_out0 = !(v$SEL1_13488_out0 || v$SEL2_7699_out0);
assign v$G10_1410_out0 = !(v$SEL1_13489_out0 || v$SEL2_7700_out0);
assign v$G10_1411_out0 = !(v$SEL1_13490_out0 || v$SEL2_7701_out0);
assign v$G10_1412_out0 = !(v$SEL1_13491_out0 || v$SEL2_7702_out0);
assign v$G10_1413_out0 = !(v$SEL1_13492_out0 || v$SEL2_7703_out0);
assign v$G10_1414_out0 = !(v$SEL1_13493_out0 || v$SEL2_7704_out0);
assign v$G10_1415_out0 = !(v$SEL1_13494_out0 || v$SEL2_7705_out0);
assign v$G10_1416_out0 = !(v$SEL1_13495_out0 || v$SEL2_7706_out0);
assign v$G10_1417_out0 = !(v$SEL1_13496_out0 || v$SEL2_7707_out0);
assign v$G10_1418_out0 = !(v$SEL1_13497_out0 || v$SEL2_7708_out0);
assign v$G10_1419_out0 = !(v$SEL1_13498_out0 || v$SEL2_7709_out0);
assign v$G10_1420_out0 = !(v$SEL1_13499_out0 || v$SEL2_7710_out0);
assign v$G10_1421_out0 = !(v$SEL1_13500_out0 || v$SEL2_7711_out0);
assign v$G6_3573_out0 = ! v$SEL2_7688_out0;
assign v$G6_3574_out0 = ! v$SEL2_7689_out0;
assign v$G6_3575_out0 = ! v$SEL2_7690_out0;
assign v$G6_3576_out0 = ! v$SEL2_7691_out0;
assign v$G6_3577_out0 = ! v$SEL2_7692_out0;
assign v$G6_3578_out0 = ! v$SEL2_7693_out0;
assign v$G6_3579_out0 = ! v$SEL2_7694_out0;
assign v$G6_3580_out0 = ! v$SEL2_7695_out0;
assign v$G6_3581_out0 = ! v$SEL2_7696_out0;
assign v$G6_3582_out0 = ! v$SEL2_7697_out0;
assign v$G6_3583_out0 = ! v$SEL2_7698_out0;
assign v$G6_3584_out0 = ! v$SEL2_7699_out0;
assign v$G6_3585_out0 = ! v$SEL2_7700_out0;
assign v$G6_3586_out0 = ! v$SEL2_7701_out0;
assign v$G6_3587_out0 = ! v$SEL2_7702_out0;
assign v$G6_3588_out0 = ! v$SEL2_7703_out0;
assign v$G6_3589_out0 = ! v$SEL2_7704_out0;
assign v$G6_3590_out0 = ! v$SEL2_7705_out0;
assign v$G6_3591_out0 = ! v$SEL2_7706_out0;
assign v$G6_3592_out0 = ! v$SEL2_7707_out0;
assign v$G6_3593_out0 = ! v$SEL2_7708_out0;
assign v$G6_3594_out0 = ! v$SEL2_7709_out0;
assign v$G6_3595_out0 = ! v$SEL2_7710_out0;
assign v$G6_3596_out0 = ! v$SEL2_7711_out0;
assign v$_4261_out0 = { v$C2_119_out0,v$SEL1_15402_out0 };
assign v$_4271_out0 = { v$C2_129_out0,v$SEL1_15412_out0 };
assign v$MUX21_4904_out0 = v$EQ21_3326_out0 ? v$SEL21_11050_out0 : v$MUX22_16466_out0;
assign v$MUX21_4905_out0 = v$EQ21_3327_out0 ? v$SEL21_11051_out0 : v$MUX22_16467_out0;
assign v$G5_5849_out0 = ! v$SEL4_6097_out0;
assign v$G5_5850_out0 = ! v$SEL4_6098_out0;
assign v$G5_5851_out0 = ! v$SEL4_6099_out0;
assign v$G5_5852_out0 = ! v$SEL4_6100_out0;
assign v$G5_5853_out0 = ! v$SEL4_6101_out0;
assign v$G5_5854_out0 = ! v$SEL4_6102_out0;
assign v$G5_5855_out0 = ! v$SEL4_6103_out0;
assign v$G5_5856_out0 = ! v$SEL4_6104_out0;
assign v$G5_5857_out0 = ! v$SEL4_6105_out0;
assign v$G5_5858_out0 = ! v$SEL4_6106_out0;
assign v$G5_5859_out0 = ! v$SEL4_6107_out0;
assign v$G5_5860_out0 = ! v$SEL4_6108_out0;
assign v$G5_5861_out0 = ! v$SEL4_6109_out0;
assign v$G5_5862_out0 = ! v$SEL4_6110_out0;
assign v$G5_5863_out0 = ! v$SEL4_6111_out0;
assign v$G5_5864_out0 = ! v$SEL4_6112_out0;
assign v$G5_5865_out0 = ! v$SEL4_6113_out0;
assign v$G5_5866_out0 = ! v$SEL4_6114_out0;
assign v$G5_5867_out0 = ! v$SEL4_6115_out0;
assign v$G5_5868_out0 = ! v$SEL4_6116_out0;
assign v$G5_5869_out0 = ! v$SEL4_6117_out0;
assign v$G5_5870_out0 = ! v$SEL4_6118_out0;
assign v$G5_5871_out0 = ! v$SEL4_6119_out0;
assign v$G5_5872_out0 = ! v$SEL4_6120_out0;
assign v$END26_6435_out0 = v$G$AD_17119_out0;
assign v$END26_6438_out0 = v$G$AD_17242_out0;
assign v$C8_7430_out0 = v$COUTD_6699_out0;
assign v$C8_7433_out0 = v$COUTD_6822_out0;
assign v$CINA_8467_out0 = v$COUTD_6722_out0;
assign v$CINA_8476_out0 = v$COUTD_6722_out0;
assign v$CINA_8477_out0 = v$COUTD_6699_out0;
assign v$CINA_8488_out0 = v$COUTD_6722_out0;
assign v$CINA_8490_out0 = v$COUTD_6722_out0;
assign v$CINA_8497_out0 = v$COUTD_6722_out0;
assign v$CINA_8498_out0 = v$COUTD_6699_out0;
assign v$CINA_8590_out0 = v$COUTD_6845_out0;
assign v$CINA_8599_out0 = v$COUTD_6845_out0;
assign v$CINA_8600_out0 = v$COUTD_6822_out0;
assign v$CINA_8611_out0 = v$COUTD_6845_out0;
assign v$CINA_8613_out0 = v$COUTD_6845_out0;
assign v$CINA_8620_out0 = v$COUTD_6845_out0;
assign v$CINA_8621_out0 = v$COUTD_6822_out0;
assign v$G11_8860_out0 = !(v$SEL3_2312_out0 || v$SEL4_6097_out0);
assign v$G11_8861_out0 = !(v$SEL3_2313_out0 || v$SEL4_6098_out0);
assign v$G11_8862_out0 = !(v$SEL3_2314_out0 || v$SEL4_6099_out0);
assign v$G11_8863_out0 = !(v$SEL3_2315_out0 || v$SEL4_6100_out0);
assign v$G11_8864_out0 = !(v$SEL3_2316_out0 || v$SEL4_6101_out0);
assign v$G11_8865_out0 = !(v$SEL3_2317_out0 || v$SEL4_6102_out0);
assign v$G11_8866_out0 = !(v$SEL3_2318_out0 || v$SEL4_6103_out0);
assign v$G11_8867_out0 = !(v$SEL3_2319_out0 || v$SEL4_6104_out0);
assign v$G11_8868_out0 = !(v$SEL3_2320_out0 || v$SEL4_6105_out0);
assign v$G11_8869_out0 = !(v$SEL3_2321_out0 || v$SEL4_6106_out0);
assign v$G11_8870_out0 = !(v$SEL3_2322_out0 || v$SEL4_6107_out0);
assign v$G11_8871_out0 = !(v$SEL3_2323_out0 || v$SEL4_6108_out0);
assign v$G11_8872_out0 = !(v$SEL3_2324_out0 || v$SEL4_6109_out0);
assign v$G11_8873_out0 = !(v$SEL3_2325_out0 || v$SEL4_6110_out0);
assign v$G11_8874_out0 = !(v$SEL3_2326_out0 || v$SEL4_6111_out0);
assign v$G11_8875_out0 = !(v$SEL3_2327_out0 || v$SEL4_6112_out0);
assign v$G11_8876_out0 = !(v$SEL3_2328_out0 || v$SEL4_6113_out0);
assign v$G11_8877_out0 = !(v$SEL3_2329_out0 || v$SEL4_6114_out0);
assign v$G11_8878_out0 = !(v$SEL3_2330_out0 || v$SEL4_6115_out0);
assign v$G11_8879_out0 = !(v$SEL3_2331_out0 || v$SEL4_6116_out0);
assign v$G11_8880_out0 = !(v$SEL3_2332_out0 || v$SEL4_6117_out0);
assign v$G11_8881_out0 = !(v$SEL3_2333_out0 || v$SEL4_6118_out0);
assign v$G11_8882_out0 = !(v$SEL3_2334_out0 || v$SEL4_6119_out0);
assign v$G11_8883_out0 = !(v$SEL3_2335_out0 || v$SEL4_6120_out0);
assign v$_8996_out0 = { v$SEL1_8711_out0,v$C1_5977_out0 };
assign v$_9006_out0 = { v$SEL1_8721_out0,v$C1_5987_out0 };
assign v$G$AB_9152_out0 = v$G$AD_17089_out0;
assign v$G$AB_9159_out0 = v$G$AD_17089_out0;
assign v$G$AB_9163_out0 = v$G$AD_17110_out0;
assign v$G$AB_9166_out0 = v$G$AD_17110_out0;
assign v$G$AB_9174_out0 = v$G$AD_17089_out0;
assign v$G$AB_9275_out0 = v$G$AD_17212_out0;
assign v$G$AB_9282_out0 = v$G$AD_17212_out0;
assign v$G$AB_9286_out0 = v$G$AD_17233_out0;
assign v$G$AB_9289_out0 = v$G$AD_17233_out0;
assign v$G$AB_9297_out0 = v$G$AD_17212_out0;
assign v$C6_9586_out0 = v$COUTD_6703_out0;
assign v$C6_9589_out0 = v$COUTD_6826_out0;
assign v$C7_10969_out0 = v$COUTD_6732_out0;
assign v$C7_10972_out0 = v$COUTD_6855_out0;
assign v$G8_12008_out0 = ! v$SEL3_2312_out0;
assign v$G8_12009_out0 = ! v$SEL3_2313_out0;
assign v$G8_12010_out0 = ! v$SEL3_2314_out0;
assign v$G8_12011_out0 = ! v$SEL3_2315_out0;
assign v$G8_12012_out0 = ! v$SEL3_2316_out0;
assign v$G8_12013_out0 = ! v$SEL3_2317_out0;
assign v$G8_12014_out0 = ! v$SEL3_2318_out0;
assign v$G8_12015_out0 = ! v$SEL3_2319_out0;
assign v$G8_12016_out0 = ! v$SEL3_2320_out0;
assign v$G8_12017_out0 = ! v$SEL3_2321_out0;
assign v$G8_12018_out0 = ! v$SEL3_2322_out0;
assign v$G8_12019_out0 = ! v$SEL3_2323_out0;
assign v$G8_12020_out0 = ! v$SEL3_2324_out0;
assign v$G8_12021_out0 = ! v$SEL3_2325_out0;
assign v$G8_12022_out0 = ! v$SEL3_2326_out0;
assign v$G8_12023_out0 = ! v$SEL3_2327_out0;
assign v$G8_12024_out0 = ! v$SEL3_2328_out0;
assign v$G8_12025_out0 = ! v$SEL3_2329_out0;
assign v$G8_12026_out0 = ! v$SEL3_2330_out0;
assign v$G8_12027_out0 = ! v$SEL3_2331_out0;
assign v$G8_12028_out0 = ! v$SEL3_2332_out0;
assign v$G8_12029_out0 = ! v$SEL3_2333_out0;
assign v$G8_12030_out0 = ! v$SEL3_2334_out0;
assign v$G8_12031_out0 = ! v$SEL3_2335_out0;
assign v$END20_13264_out0 = v$G$AD_17099_out0;
assign v$END20_13267_out0 = v$G$AD_17222_out0;
assign v$END28_13669_out0 = v$G$AD_17110_out0;
assign v$END28_13672_out0 = v$G$AD_17233_out0;
assign v$C11_14796_out0 = v$COUTD_6722_out0;
assign v$C11_14799_out0 = v$COUTD_6845_out0;
assign v$END22_15484_out0 = v$G$AD_17120_out0;
assign v$END22_15487_out0 = v$G$AD_17243_out0;
assign v$END24_16403_out0 = v$G$AD_17098_out0;
assign v$END24_16406_out0 = v$G$AD_17221_out0;
assign v$END61_17956_out0 = v$COUTD_6730_out0;
assign v$END61_17959_out0 = v$COUTD_6853_out0;
assign {v$A8A_1505_out1,v$A8A_1505_out0 } = v$A7_15307_out0 + v$B7_17040_out0 + v$C6_9586_out0;
assign {v$A8A_1508_out1,v$A8A_1508_out0 } = v$A7_15310_out0 + v$B7_17043_out0 + v$C6_9589_out0;
assign v$MUX1_2365_out0 = v$LEFT$SHIT_3057_out0 ? v$_4261_out0 : v$_8996_out0;
assign v$MUX1_2375_out0 = v$LEFT$SHIT_3067_out0 ? v$_4271_out0 : v$_9006_out0;
assign {v$A17A_2487_out1,v$A17A_2487_out0 } = v$A12_3138_out0 + v$B12_1950_out0 + v$C11_14796_out0;
assign {v$A17A_2490_out1,v$A17A_2490_out0 } = v$A12_3141_out0 + v$B12_1953_out0 + v$C11_14799_out0;
assign v$G5_4535_out0 = v$G$AB_9152_out0 && v$P$CD_10470_out0;
assign v$G5_4542_out0 = v$G$AB_9159_out0 && v$P$CD_10477_out0;
assign v$G5_4546_out0 = v$G$AB_9163_out0 && v$P$CD_10481_out0;
assign v$G5_4549_out0 = v$G$AB_9166_out0 && v$P$CD_10484_out0;
assign v$G5_4557_out0 = v$G$AB_9174_out0 && v$P$CD_10492_out0;
assign v$G5_4658_out0 = v$G$AB_9275_out0 && v$P$CD_10593_out0;
assign v$G5_4665_out0 = v$G$AB_9282_out0 && v$P$CD_10600_out0;
assign v$G5_4669_out0 = v$G$AB_9286_out0 && v$P$CD_10604_out0;
assign v$G5_4672_out0 = v$G$AB_9289_out0 && v$P$CD_10607_out0;
assign v$G5_4680_out0 = v$G$AB_9297_out0 && v$P$CD_10615_out0;
assign v$C6_7055_out0 = v$C6_9586_out0;
assign v$C6_7058_out0 = v$C6_9589_out0;
assign v$C11_9510_out0 = v$C11_14796_out0;
assign v$C11_9513_out0 = v$C11_14799_out0;
assign {v$A9A_10411_out1,v$A9A_10411_out0 } = v$A8_18090_out0 + v$B8_13138_out0 + v$C7_10969_out0;
assign {v$A9A_10414_out1,v$A9A_10414_out0 } = v$A8_18093_out0 + v$B8_13141_out0 + v$C7_10972_out0;
assign v$MUX20_11366_out0 = v$EQ20_9948_out0 ? v$SEL20_8176_out0 : v$MUX21_4904_out0;
assign v$MUX20_11367_out0 = v$EQ20_9949_out0 ? v$SEL20_8177_out0 : v$MUX21_4905_out0;
assign v$G8_11398_out0 = v$CINA_8467_out0 && v$P$AB_2004_out0;
assign v$G8_11407_out0 = v$CINA_8476_out0 && v$P$AB_2013_out0;
assign v$G8_11408_out0 = v$CINA_8477_out0 && v$P$AB_2014_out0;
assign v$G8_11419_out0 = v$CINA_8488_out0 && v$P$AB_2025_out0;
assign v$G8_11421_out0 = v$CINA_8490_out0 && v$P$AB_2027_out0;
assign v$G8_11428_out0 = v$CINA_8497_out0 && v$P$AB_2034_out0;
assign v$G8_11429_out0 = v$CINA_8498_out0 && v$P$AB_2035_out0;
assign v$G8_11521_out0 = v$CINA_8590_out0 && v$P$AB_2127_out0;
assign v$G8_11530_out0 = v$CINA_8599_out0 && v$P$AB_2136_out0;
assign v$G8_11531_out0 = v$CINA_8600_out0 && v$P$AB_2137_out0;
assign v$G8_11542_out0 = v$CINA_8611_out0 && v$P$AB_2148_out0;
assign v$G8_11544_out0 = v$CINA_8613_out0 && v$P$AB_2150_out0;
assign v$G8_11551_out0 = v$CINA_8620_out0 && v$P$AB_2157_out0;
assign v$G8_11552_out0 = v$CINA_8621_out0 && v$P$AB_2158_out0;
assign v$END51_11676_out0 = v$P$AD_696_out0;
assign v$END51_11679_out0 = v$P$AD_819_out0;
assign v$G3_12680_out0 = v$G10_1398_out0 && v$G11_8860_out0;
assign v$G3_12681_out0 = v$G10_1399_out0 && v$G11_8861_out0;
assign v$G3_12682_out0 = v$G10_1400_out0 && v$G11_8862_out0;
assign v$G3_12683_out0 = v$G10_1401_out0 && v$G11_8863_out0;
assign v$G3_12684_out0 = v$G10_1402_out0 && v$G11_8864_out0;
assign v$G3_12685_out0 = v$G10_1403_out0 && v$G11_8865_out0;
assign v$G3_12686_out0 = v$G10_1404_out0 && v$G11_8866_out0;
assign v$G3_12687_out0 = v$G10_1405_out0 && v$G11_8867_out0;
assign v$G3_12688_out0 = v$G10_1406_out0 && v$G11_8868_out0;
assign v$G3_12689_out0 = v$G10_1407_out0 && v$G11_8869_out0;
assign v$G3_12690_out0 = v$G10_1408_out0 && v$G11_8870_out0;
assign v$G3_12691_out0 = v$G10_1409_out0 && v$G11_8871_out0;
assign v$G3_12692_out0 = v$G10_1410_out0 && v$G11_8872_out0;
assign v$G3_12693_out0 = v$G10_1411_out0 && v$G11_8873_out0;
assign v$G3_12694_out0 = v$G10_1412_out0 && v$G11_8874_out0;
assign v$G3_12695_out0 = v$G10_1413_out0 && v$G11_8875_out0;
assign v$G3_12696_out0 = v$G10_1414_out0 && v$G11_8876_out0;
assign v$G3_12697_out0 = v$G10_1415_out0 && v$G11_8877_out0;
assign v$G3_12698_out0 = v$G10_1416_out0 && v$G11_8878_out0;
assign v$G3_12699_out0 = v$G10_1417_out0 && v$G11_8879_out0;
assign v$G3_12700_out0 = v$G10_1418_out0 && v$G11_8880_out0;
assign v$G3_12701_out0 = v$G10_1419_out0 && v$G11_8881_out0;
assign v$G3_12702_out0 = v$G10_1420_out0 && v$G11_8882_out0;
assign v$G3_12703_out0 = v$G10_1421_out0 && v$G11_8883_out0;
assign {v$A10A_16002_out1,v$A10A_16002_out0 } = v$A9_3435_out0 + v$B9_4065_out0 + v$C8_7430_out0;
assign {v$A10A_16005_out1,v$A10A_16005_out0 } = v$A9_3438_out0 + v$B9_4068_out0 + v$C8_7433_out0;
assign v$C7_16430_out0 = v$C7_10969_out0;
assign v$C7_16433_out0 = v$C7_10972_out0;
assign v$G9_17606_out0 = v$G8_12008_out0 && v$G5_5849_out0;
assign v$G9_17607_out0 = v$G8_12009_out0 && v$G5_5850_out0;
assign v$G9_17608_out0 = v$G8_12010_out0 && v$G5_5851_out0;
assign v$G9_17609_out0 = v$G8_12011_out0 && v$G5_5852_out0;
assign v$G9_17610_out0 = v$G8_12012_out0 && v$G5_5853_out0;
assign v$G9_17611_out0 = v$G8_12013_out0 && v$G5_5854_out0;
assign v$G9_17612_out0 = v$G8_12014_out0 && v$G5_5855_out0;
assign v$G9_17613_out0 = v$G8_12015_out0 && v$G5_5856_out0;
assign v$G9_17614_out0 = v$G8_12016_out0 && v$G5_5857_out0;
assign v$G9_17615_out0 = v$G8_12017_out0 && v$G5_5858_out0;
assign v$G9_17616_out0 = v$G8_12018_out0 && v$G5_5859_out0;
assign v$G9_17617_out0 = v$G8_12019_out0 && v$G5_5860_out0;
assign v$G9_17618_out0 = v$G8_12020_out0 && v$G5_5861_out0;
assign v$G9_17619_out0 = v$G8_12021_out0 && v$G5_5862_out0;
assign v$G9_17620_out0 = v$G8_12022_out0 && v$G5_5863_out0;
assign v$G9_17621_out0 = v$G8_12023_out0 && v$G5_5864_out0;
assign v$G9_17622_out0 = v$G8_12024_out0 && v$G5_5865_out0;
assign v$G9_17623_out0 = v$G8_12025_out0 && v$G5_5866_out0;
assign v$G9_17624_out0 = v$G8_12026_out0 && v$G5_5867_out0;
assign v$G9_17625_out0 = v$G8_12027_out0 && v$G5_5868_out0;
assign v$G9_17626_out0 = v$G8_12028_out0 && v$G5_5869_out0;
assign v$G9_17627_out0 = v$G8_12029_out0 && v$G5_5870_out0;
assign v$G9_17628_out0 = v$G8_12030_out0 && v$G5_5871_out0;
assign v$G9_17629_out0 = v$G8_12031_out0 && v$G5_5872_out0;
assign v$G7_18149_out0 = v$G6_3573_out0 || v$SEL3_2312_out0;
assign v$G7_18150_out0 = v$G6_3574_out0 || v$SEL3_2313_out0;
assign v$G7_18151_out0 = v$G6_3575_out0 || v$SEL3_2314_out0;
assign v$G7_18152_out0 = v$G6_3576_out0 || v$SEL3_2315_out0;
assign v$G7_18153_out0 = v$G6_3577_out0 || v$SEL3_2316_out0;
assign v$G7_18154_out0 = v$G6_3578_out0 || v$SEL3_2317_out0;
assign v$G7_18155_out0 = v$G6_3579_out0 || v$SEL3_2318_out0;
assign v$G7_18156_out0 = v$G6_3580_out0 || v$SEL3_2319_out0;
assign v$G7_18157_out0 = v$G6_3581_out0 || v$SEL3_2320_out0;
assign v$G7_18158_out0 = v$G6_3582_out0 || v$SEL3_2321_out0;
assign v$G7_18159_out0 = v$G6_3583_out0 || v$SEL3_2322_out0;
assign v$G7_18160_out0 = v$G6_3584_out0 || v$SEL3_2323_out0;
assign v$G7_18161_out0 = v$G6_3585_out0 || v$SEL3_2324_out0;
assign v$G7_18162_out0 = v$G6_3586_out0 || v$SEL3_2325_out0;
assign v$G7_18163_out0 = v$G6_3587_out0 || v$SEL3_2326_out0;
assign v$G7_18164_out0 = v$G6_3588_out0 || v$SEL3_2327_out0;
assign v$G7_18165_out0 = v$G6_3589_out0 || v$SEL3_2328_out0;
assign v$G7_18166_out0 = v$G6_3590_out0 || v$SEL3_2329_out0;
assign v$G7_18167_out0 = v$G6_3591_out0 || v$SEL3_2330_out0;
assign v$G7_18168_out0 = v$G6_3592_out0 || v$SEL3_2331_out0;
assign v$G7_18169_out0 = v$G6_3593_out0 || v$SEL3_2332_out0;
assign v$G7_18170_out0 = v$G6_3594_out0 || v$SEL3_2333_out0;
assign v$G7_18171_out0 = v$G6_3595_out0 || v$SEL3_2334_out0;
assign v$G7_18172_out0 = v$G6_3596_out0 || v$SEL3_2335_out0;
assign v$END49_18450_out0 = v$P$AD_715_out0;
assign v$END49_18453_out0 = v$P$AD_838_out0;
assign v$C8_18497_out0 = v$C8_7430_out0;
assign v$C8_18500_out0 = v$C8_7433_out0;
assign v$MUX2_2498_out0 = v$EN_1337_out0 ? v$MUX1_2365_out0 : v$IN_5024_out0;
assign v$MUX2_2501_out0 = v$EN_1340_out0 ? v$MUX1_2375_out0 : v$IN_5027_out0;
assign v$END7_3359_out0 = v$A8A_1505_out1;
assign v$END7_3362_out0 = v$A8A_1508_out1;
assign v$_3636_out0 = { v$A6A_3121_out0,v$A8A_1505_out0 };
assign v$_3639_out0 = { v$A6A_3124_out0,v$A8A_1508_out0 };
assign v$END8_3901_out0 = v$A9A_10411_out1;
assign v$END8_3904_out0 = v$A9A_10414_out1;
assign v$END9_4233_out0 = v$A10A_16002_out1;
assign v$END9_4236_out0 = v$A10A_16005_out1;
assign v$MUX19_6376_out0 = v$EQ19_5444_out0 ? v$SEL19_12817_out0 : v$MUX20_11366_out0;
assign v$MUX19_6377_out0 = v$EQ19_5445_out0 ? v$SEL19_12818_out0 : v$MUX20_11367_out0;
assign v$ENDw_9551_out0 = v$A17A_2487_out1;
assign v$ENDw_9554_out0 = v$A17A_2490_out1;
assign v$G7_9638_out0 = v$G8_11398_out0 && v$P$CD_10457_out0;
assign v$G7_9647_out0 = v$G8_11407_out0 && v$P$CD_10466_out0;
assign v$G7_9648_out0 = v$G8_11408_out0 && v$P$CD_10467_out0;
assign v$G7_9659_out0 = v$G8_11419_out0 && v$P$CD_10478_out0;
assign v$G7_9661_out0 = v$G8_11421_out0 && v$P$CD_10480_out0;
assign v$G7_9668_out0 = v$G8_11428_out0 && v$P$CD_10487_out0;
assign v$G7_9669_out0 = v$G8_11429_out0 && v$P$CD_10488_out0;
assign v$G7_9761_out0 = v$G8_11521_out0 && v$P$CD_10580_out0;
assign v$G7_9770_out0 = v$G8_11530_out0 && v$P$CD_10589_out0;
assign v$G7_9771_out0 = v$G8_11531_out0 && v$P$CD_10590_out0;
assign v$G7_9782_out0 = v$G8_11542_out0 && v$P$CD_10601_out0;
assign v$G7_9784_out0 = v$G8_11544_out0 && v$P$CD_10603_out0;
assign v$G7_9791_out0 = v$G8_11551_out0 && v$P$CD_10610_out0;
assign v$G7_9792_out0 = v$G8_11552_out0 && v$P$CD_10611_out0;
assign v$G4_11127_out0 = v$G5_4535_out0 || v$G$CD_930_out0;
assign v$G4_11134_out0 = v$G5_4542_out0 || v$G$CD_937_out0;
assign v$G4_11138_out0 = v$G5_4546_out0 || v$G$CD_941_out0;
assign v$G4_11141_out0 = v$G5_4549_out0 || v$G$CD_944_out0;
assign v$G4_11149_out0 = v$G5_4557_out0 || v$G$CD_952_out0;
assign v$G4_11250_out0 = v$G5_4658_out0 || v$G$CD_1053_out0;
assign v$G4_11257_out0 = v$G5_4665_out0 || v$G$CD_1060_out0;
assign v$G4_11261_out0 = v$G5_4669_out0 || v$G$CD_1064_out0;
assign v$G4_11264_out0 = v$G5_4672_out0 || v$G$CD_1067_out0;
assign v$G4_11272_out0 = v$G5_4680_out0 || v$G$CD_1075_out0;
assign v$Z_12571_out0 = v$G3_12680_out0;
assign v$Z_12572_out0 = v$G3_12681_out0;
assign v$Z_12573_out0 = v$G3_12682_out0;
assign v$Z_12574_out0 = v$G3_12683_out0;
assign v$Z_12575_out0 = v$G3_12684_out0;
assign v$Z_12576_out0 = v$G3_12685_out0;
assign v$Z_12577_out0 = v$G3_12686_out0;
assign v$Z_12578_out0 = v$G3_12687_out0;
assign v$Z_12579_out0 = v$G3_12688_out0;
assign v$Z_12580_out0 = v$G3_12689_out0;
assign v$Z_12581_out0 = v$G3_12690_out0;
assign v$Z_12582_out0 = v$G3_12691_out0;
assign v$Z_12583_out0 = v$G3_12692_out0;
assign v$Z_12584_out0 = v$G3_12693_out0;
assign v$Z_12585_out0 = v$G3_12694_out0;
assign v$Z_12586_out0 = v$G3_12695_out0;
assign v$Z_12587_out0 = v$G3_12696_out0;
assign v$Z_12588_out0 = v$G3_12697_out0;
assign v$Z_12589_out0 = v$G3_12698_out0;
assign v$Z_12590_out0 = v$G3_12699_out0;
assign v$Z_12591_out0 = v$G3_12700_out0;
assign v$Z_12592_out0 = v$G3_12701_out0;
assign v$Z_12593_out0 = v$G3_12702_out0;
assign v$Z_12594_out0 = v$G3_12703_out0;
assign v$_15013_out0 = { v$A9A_10411_out0,v$A10A_16002_out0 };
assign v$_15016_out0 = { v$A9A_10414_out0,v$A10A_16005_out0 };
assign v$_16310_out0 = { v$C6_7055_out0,v$C7_16430_out0 };
assign v$_16313_out0 = { v$C6_7058_out0,v$C7_16433_out0 };
assign v$G4_17541_out0 = v$G7_18149_out0 && v$G5_5849_out0;
assign v$G4_17542_out0 = v$G7_18150_out0 && v$G5_5850_out0;
assign v$G4_17543_out0 = v$G7_18151_out0 && v$G5_5851_out0;
assign v$G4_17544_out0 = v$G7_18152_out0 && v$G5_5852_out0;
assign v$G4_17545_out0 = v$G7_18153_out0 && v$G5_5853_out0;
assign v$G4_17546_out0 = v$G7_18154_out0 && v$G5_5854_out0;
assign v$G4_17547_out0 = v$G7_18155_out0 && v$G5_5855_out0;
assign v$G4_17548_out0 = v$G7_18156_out0 && v$G5_5856_out0;
assign v$G4_17549_out0 = v$G7_18157_out0 && v$G5_5857_out0;
assign v$G4_17550_out0 = v$G7_18158_out0 && v$G5_5858_out0;
assign v$G4_17551_out0 = v$G7_18159_out0 && v$G5_5859_out0;
assign v$G4_17552_out0 = v$G7_18160_out0 && v$G5_5860_out0;
assign v$G4_17553_out0 = v$G7_18161_out0 && v$G5_5861_out0;
assign v$G4_17554_out0 = v$G7_18162_out0 && v$G5_5862_out0;
assign v$G4_17555_out0 = v$G7_18163_out0 && v$G5_5863_out0;
assign v$G4_17556_out0 = v$G7_18164_out0 && v$G5_5864_out0;
assign v$G4_17557_out0 = v$G7_18165_out0 && v$G5_5865_out0;
assign v$G4_17558_out0 = v$G7_18166_out0 && v$G5_5866_out0;
assign v$G4_17559_out0 = v$G7_18167_out0 && v$G5_5867_out0;
assign v$G4_17560_out0 = v$G7_18168_out0 && v$G5_5868_out0;
assign v$G4_17561_out0 = v$G7_18169_out0 && v$G5_5869_out0;
assign v$G4_17562_out0 = v$G7_18170_out0 && v$G5_5870_out0;
assign v$G4_17563_out0 = v$G7_18171_out0 && v$G5_5871_out0;
assign v$G4_17564_out0 = v$G7_18172_out0 && v$G5_5872_out0;
assign v$G6_436_out0 = v$G4_11114_out0 || v$G7_9638_out0;
assign v$G6_445_out0 = v$G4_11123_out0 || v$G7_9647_out0;
assign v$G6_446_out0 = v$G4_11124_out0 || v$G7_9648_out0;
assign v$G6_457_out0 = v$G4_11135_out0 || v$G7_9659_out0;
assign v$G6_459_out0 = v$G4_11137_out0 || v$G7_9661_out0;
assign v$G6_466_out0 = v$G4_11144_out0 || v$G7_9668_out0;
assign v$G6_467_out0 = v$G4_11145_out0 || v$G7_9669_out0;
assign v$G6_559_out0 = v$G4_11237_out0 || v$G7_9761_out0;
assign v$G6_568_out0 = v$G4_11246_out0 || v$G7_9770_out0;
assign v$G6_569_out0 = v$G4_11247_out0 || v$G7_9771_out0;
assign v$G6_580_out0 = v$G4_11258_out0 || v$G7_9782_out0;
assign v$G6_582_out0 = v$G4_11260_out0 || v$G7_9784_out0;
assign v$G6_589_out0 = v$G4_11267_out0 || v$G7_9791_out0;
assign v$G6_590_out0 = v$G4_11268_out0 || v$G7_9792_out0;
assign v$MUX18_4860_out0 = v$EQ18_12808_out0 ? v$SEL18_11381_out0 : v$MUX19_6376_out0;
assign v$MUX18_4861_out0 = v$EQ18_12809_out0 ? v$SEL18_11382_out0 : v$MUX19_6377_out0;
assign v$_6284_out0 = { v$G4_17541_out0,v$G9_17606_out0 };
assign v$_6285_out0 = { v$G4_17542_out0,v$G9_17607_out0 };
assign v$_6286_out0 = { v$G4_17543_out0,v$G9_17608_out0 };
assign v$_6287_out0 = { v$G4_17544_out0,v$G9_17609_out0 };
assign v$_6288_out0 = { v$G4_17545_out0,v$G9_17610_out0 };
assign v$_6289_out0 = { v$G4_17546_out0,v$G9_17611_out0 };
assign v$_6290_out0 = { v$G4_17547_out0,v$G9_17612_out0 };
assign v$_6291_out0 = { v$G4_17548_out0,v$G9_17613_out0 };
assign v$_6292_out0 = { v$G4_17549_out0,v$G9_17614_out0 };
assign v$_6293_out0 = { v$G4_17550_out0,v$G9_17615_out0 };
assign v$_6294_out0 = { v$G4_17551_out0,v$G9_17616_out0 };
assign v$_6295_out0 = { v$G4_17552_out0,v$G9_17617_out0 };
assign v$_6296_out0 = { v$G4_17553_out0,v$G9_17618_out0 };
assign v$_6297_out0 = { v$G4_17554_out0,v$G9_17619_out0 };
assign v$_6298_out0 = { v$G4_17555_out0,v$G9_17620_out0 };
assign v$_6299_out0 = { v$G4_17556_out0,v$G9_17621_out0 };
assign v$_6300_out0 = { v$G4_17557_out0,v$G9_17622_out0 };
assign v$_6301_out0 = { v$G4_17558_out0,v$G9_17623_out0 };
assign v$_6302_out0 = { v$G4_17559_out0,v$G9_17624_out0 };
assign v$_6303_out0 = { v$G4_17560_out0,v$G9_17625_out0 };
assign v$_6304_out0 = { v$G4_17561_out0,v$G9_17626_out0 };
assign v$_6305_out0 = { v$G4_17562_out0,v$G9_17627_out0 };
assign v$_6306_out0 = { v$G4_17563_out0,v$G9_17628_out0 };
assign v$_6307_out0 = { v$G4_17564_out0,v$G9_17629_out0 };
assign v$Z2_6325_out0 = v$Z_12573_out0;
assign v$Z2_6326_out0 = v$Z_12577_out0;
assign v$Z2_6327_out0 = v$Z_12581_out0;
assign v$Z2_6329_out0 = v$Z_12585_out0;
assign v$Z2_6330_out0 = v$Z_12589_out0;
assign v$Z2_6331_out0 = v$Z_12593_out0;
assign v$_7404_out0 = { v$_2453_out0,v$_16310_out0 };
assign v$_7407_out0 = { v$_2456_out0,v$_16313_out0 };
assign v$Z4_7921_out0 = v$Z_12574_out0;
assign v$Z4_7922_out0 = v$Z_12578_out0;
assign v$Z4_7923_out0 = v$Z_12582_out0;
assign v$Z4_7924_out0 = v$Z_12586_out0;
assign v$Z4_7925_out0 = v$Z_12590_out0;
assign v$Z4_7926_out0 = v$Z_12594_out0;
assign v$OUT_14917_out0 = v$MUX2_2498_out0;
assign v$OUT_14927_out0 = v$MUX2_2501_out0;
assign v$Z1_16999_out0 = v$Z_12572_out0;
assign v$Z1_17000_out0 = v$Z_12576_out0;
assign v$Z1_17001_out0 = v$Z_12580_out0;
assign v$Z1_17003_out0 = v$Z_12584_out0;
assign v$Z1_17004_out0 = v$Z_12588_out0;
assign v$Z1_17005_out0 = v$Z_12592_out0;
assign v$G$AD_17102_out0 = v$G4_11127_out0;
assign v$G$AD_17109_out0 = v$G4_11134_out0;
assign v$G$AD_17113_out0 = v$G4_11138_out0;
assign v$G$AD_17116_out0 = v$G4_11141_out0;
assign v$G$AD_17124_out0 = v$G4_11149_out0;
assign v$G$AD_17225_out0 = v$G4_11250_out0;
assign v$G$AD_17232_out0 = v$G4_11257_out0;
assign v$G$AD_17236_out0 = v$G4_11261_out0;
assign v$G$AD_17239_out0 = v$G4_11264_out0;
assign v$G$AD_17247_out0 = v$G4_11272_out0;
assign v$Z3_17780_out0 = v$Z_12571_out0;
assign v$Z3_17781_out0 = v$Z_12575_out0;
assign v$Z3_17782_out0 = v$Z_12579_out0;
assign v$Z3_17784_out0 = v$Z_12583_out0;
assign v$Z3_17785_out0 = v$Z_12587_out0;
assign v$Z3_17786_out0 = v$Z_12591_out0;
assign v$_17964_out0 = { v$_82_out0,v$_3636_out0 };
assign v$_17967_out0 = { v$_85_out0,v$_3639_out0 };
assign v$END32_2470_out0 = v$G$AD_17116_out0;
assign v$END32_2473_out0 = v$G$AD_17239_out0;
assign v$IN_5165_out0 = v$OUT_14917_out0;
assign v$IN_5175_out0 = v$OUT_14927_out0;
assign v$G4_6055_out0 = ! v$Z4_7921_out0;
assign v$G4_6056_out0 = ! v$Z4_7922_out0;
assign v$G4_6057_out0 = ! v$Z4_7923_out0;
assign v$G4_6058_out0 = ! v$Z4_7924_out0;
assign v$G4_6059_out0 = ! v$Z4_7925_out0;
assign v$G4_6060_out0 = ! v$Z4_7926_out0;
assign v$G6_6174_out0 = ! v$Z2_6325_out0;
assign v$G6_6175_out0 = ! v$Z2_6326_out0;
assign v$G6_6176_out0 = ! v$Z2_6327_out0;
assign v$G6_6178_out0 = ! v$Z2_6329_out0;
assign v$G6_6179_out0 = ! v$Z2_6330_out0;
assign v$G6_6180_out0 = ! v$Z2_6331_out0;
assign v$Y_6501_out0 = v$_6284_out0;
assign v$Y_6502_out0 = v$_6285_out0;
assign v$Y_6503_out0 = v$_6286_out0;
assign v$Y_6504_out0 = v$_6287_out0;
assign v$Y_6505_out0 = v$_6288_out0;
assign v$Y_6506_out0 = v$_6289_out0;
assign v$Y_6507_out0 = v$_6290_out0;
assign v$Y_6508_out0 = v$_6291_out0;
assign v$Y_6509_out0 = v$_6292_out0;
assign v$Y_6510_out0 = v$_6293_out0;
assign v$Y_6511_out0 = v$_6294_out0;
assign v$Y_6512_out0 = v$_6295_out0;
assign v$Y_6513_out0 = v$_6296_out0;
assign v$Y_6514_out0 = v$_6297_out0;
assign v$Y_6515_out0 = v$_6298_out0;
assign v$Y_6516_out0 = v$_6299_out0;
assign v$Y_6517_out0 = v$_6300_out0;
assign v$Y_6518_out0 = v$_6301_out0;
assign v$Y_6519_out0 = v$_6302_out0;
assign v$Y_6520_out0 = v$_6303_out0;
assign v$Y_6521_out0 = v$_6304_out0;
assign v$Y_6522_out0 = v$_6305_out0;
assign v$Y_6523_out0 = v$_6306_out0;
assign v$Y_6524_out0 = v$_6307_out0;
assign v$COUTD_6696_out0 = v$G6_436_out0;
assign v$COUTD_6705_out0 = v$G6_445_out0;
assign v$COUTD_6706_out0 = v$G6_446_out0;
assign v$COUTD_6717_out0 = v$G6_457_out0;
assign v$COUTD_6719_out0 = v$G6_459_out0;
assign v$COUTD_6726_out0 = v$G6_466_out0;
assign v$COUTD_6727_out0 = v$G6_467_out0;
assign v$COUTD_6819_out0 = v$G6_559_out0;
assign v$COUTD_6828_out0 = v$G6_568_out0;
assign v$COUTD_6829_out0 = v$G6_569_out0;
assign v$COUTD_6840_out0 = v$G6_580_out0;
assign v$COUTD_6842_out0 = v$G6_582_out0;
assign v$COUTD_6849_out0 = v$G6_589_out0;
assign v$COUTD_6850_out0 = v$G6_590_out0;
assign v$_7790_out0 = { v$_7253_out0,v$_7404_out0 };
assign v$_7793_out0 = { v$_7256_out0,v$_7407_out0 };
assign v$G$AB_9145_out0 = v$G$AD_17109_out0;
assign v$G$AB_9164_out0 = v$G$AD_17109_out0;
assign v$G$AB_9268_out0 = v$G$AD_17232_out0;
assign v$G$AB_9287_out0 = v$G$AD_17232_out0;
assign v$END43_13192_out0 = v$G$AD_17124_out0;
assign v$END43_13195_out0 = v$G$AD_17247_out0;
assign v$END46_15045_out0 = v$G$AD_17109_out0;
assign v$END46_15048_out0 = v$G$AD_17232_out0;
assign v$G9_15203_out0 = v$Z1_16999_out0 && v$Z2_6325_out0;
assign v$G9_15204_out0 = v$Z1_17000_out0 && v$Z2_6326_out0;
assign v$G9_15205_out0 = v$Z1_17001_out0 && v$Z2_6327_out0;
assign v$G9_15207_out0 = v$Z1_17003_out0 && v$Z2_6329_out0;
assign v$G9_15208_out0 = v$Z1_17004_out0 && v$Z2_6330_out0;
assign v$G9_15209_out0 = v$Z1_17005_out0 && v$Z2_6331_out0;
assign v$END30_15713_out0 = v$G$AD_17113_out0;
assign v$END30_15716_out0 = v$G$AD_17236_out0;
assign v$MUX17_16538_out0 = v$EQ17_5881_out0 ? v$SEL17_16071_out0 : v$MUX18_4860_out0;
assign v$MUX17_16539_out0 = v$EQ17_5882_out0 ? v$SEL17_16072_out0 : v$MUX18_4861_out0;
assign v$END41_16665_out0 = v$G$AD_17102_out0;
assign v$END41_16668_out0 = v$G$AD_17225_out0;
assign v$G5_17509_out0 = ! v$Z3_17780_out0;
assign v$G5_17510_out0 = ! v$Z3_17781_out0;
assign v$G5_17511_out0 = ! v$Z3_17782_out0;
assign v$G5_17512_out0 = ! v$Z3_17784_out0;
assign v$G5_17513_out0 = ! v$Z3_17785_out0;
assign v$G5_17514_out0 = ! v$Z3_17786_out0;
assign v$_17748_out0 = { v$_10355_out0,v$_17964_out0 };
assign v$_17751_out0 = { v$_10358_out0,v$_17967_out0 };
assign v$C14_279_out0 = v$COUTD_6717_out0;
assign v$C14_282_out0 = v$COUTD_6840_out0;
assign v$C17_2520_out0 = v$COUTD_6696_out0;
assign v$C17_2523_out0 = v$COUTD_6819_out0;
assign v$IN_3860_out0 = v$IN_5165_out0;
assign v$IN_3863_out0 = v$IN_5175_out0;
assign v$_3979_out0 = { v$Y_6504_out0,v$C3_3304_out0 };
assign v$_3980_out0 = { v$Y_6508_out0,v$C3_3305_out0 };
assign v$_3981_out0 = { v$Y_6512_out0,v$C3_3306_out0 };
assign v$_3982_out0 = { v$Y_6516_out0,v$C3_3307_out0 };
assign v$_3983_out0 = { v$Y_6520_out0,v$C3_3308_out0 };
assign v$_3984_out0 = { v$Y_6524_out0,v$C3_3309_out0 };
assign v$G5_4528_out0 = v$G$AB_9145_out0 && v$P$CD_10463_out0;
assign v$G5_4547_out0 = v$G$AB_9164_out0 && v$P$CD_10482_out0;
assign v$G5_4651_out0 = v$G$AB_9268_out0 && v$P$CD_10586_out0;
assign v$G5_4670_out0 = v$G$AB_9287_out0 && v$P$CD_10605_out0;
assign v$C23_4843_out0 = v$COUTD_6719_out0;
assign v$C23_4846_out0 = v$COUTD_6842_out0;
assign v$_5094_out0 = { v$Y_6503_out0,v$C5_16913_out0 };
assign v$_5095_out0 = { v$Y_6507_out0,v$C5_16914_out0 };
assign v$_5096_out0 = { v$Y_6511_out0,v$C5_16915_out0 };
assign v$_5098_out0 = { v$Y_6515_out0,v$C5_16917_out0 };
assign v$_5099_out0 = { v$Y_6519_out0,v$C5_16918_out0 };
assign v$_5100_out0 = { v$Y_6523_out0,v$C5_16919_out0 };
assign v$C9_5937_out0 = v$COUTD_6706_out0;
assign v$C9_5940_out0 = v$COUTD_6829_out0;
assign v$CINA_8480_out0 = v$COUTD_6696_out0;
assign v$CINA_8487_out0 = v$COUTD_6696_out0;
assign v$CINA_8491_out0 = v$COUTD_6717_out0;
assign v$CINA_8494_out0 = v$COUTD_6717_out0;
assign v$CINA_8502_out0 = v$COUTD_6696_out0;
assign v$CINA_8603_out0 = v$COUTD_6819_out0;
assign v$CINA_8610_out0 = v$COUTD_6819_out0;
assign v$CINA_8614_out0 = v$COUTD_6840_out0;
assign v$CINA_8617_out0 = v$COUTD_6840_out0;
assign v$CINA_8625_out0 = v$COUTD_6819_out0;
assign v$_8785_out0 = { v$Y_6502_out0,v$C6_6539_out0 };
assign v$_8786_out0 = { v$Y_6506_out0,v$C6_6540_out0 };
assign v$_8787_out0 = { v$Y_6510_out0,v$C6_6541_out0 };
assign v$_8789_out0 = { v$Y_6514_out0,v$C6_6543_out0 };
assign v$_8790_out0 = { v$Y_6518_out0,v$C6_6544_out0 };
assign v$_8791_out0 = { v$Y_6522_out0,v$C6_6545_out0 };
assign v$_8899_out0 = { v$Y_6501_out0,v$C4_16512_out0 };
assign v$_8900_out0 = { v$Y_6505_out0,v$C4_16513_out0 };
assign v$_8901_out0 = { v$Y_6509_out0,v$C4_16514_out0 };
assign v$_8903_out0 = { v$Y_6513_out0,v$C4_16516_out0 };
assign v$_8904_out0 = { v$Y_6517_out0,v$C4_16517_out0 };
assign v$_8905_out0 = { v$Y_6521_out0,v$C4_16518_out0 };
assign v$G7_9854_out0 = v$G9_15203_out0 && v$Z3_17780_out0;
assign v$G7_9855_out0 = v$G9_15204_out0 && v$Z3_17781_out0;
assign v$G7_9856_out0 = v$G9_15205_out0 && v$Z3_17782_out0;
assign v$G7_9858_out0 = v$G9_15207_out0 && v$Z3_17784_out0;
assign v$G7_9859_out0 = v$G9_15208_out0 && v$Z3_17785_out0;
assign v$G7_9860_out0 = v$G9_15209_out0 && v$Z3_17786_out0;
assign v$C13_11776_out0 = v$COUTD_6726_out0;
assign v$C13_11779_out0 = v$COUTD_6849_out0;
assign v$C10_12732_out0 = v$COUTD_6727_out0;
assign v$C10_12735_out0 = v$COUTD_6850_out0;
assign v$C12_13520_out0 = v$COUTD_6705_out0;
assign v$C12_13523_out0 = v$COUTD_6828_out0;
assign v$MUX16_16764_out0 = v$EQ16_8288_out0 ? v$SEL16_16896_out0 : v$MUX17_16538_out0;
assign v$MUX16_16765_out0 = v$EQ16_8289_out0 ? v$SEL16_16897_out0 : v$MUX17_16539_out0;
assign v$C14_325_out0 = v$C14_279_out0;
assign v$C14_328_out0 = v$C14_282_out0;
assign v$C10_1940_out0 = v$C10_12732_out0;
assign v$C10_1943_out0 = v$C10_12735_out0;
assign v$MUX5_4058_out0 = v$G6_6174_out0 ? v$_5094_out0 : v$_8785_out0;
assign v$MUX5_4059_out0 = v$G6_6175_out0 ? v$_5095_out0 : v$_8786_out0;
assign v$MUX5_4060_out0 = v$G6_6176_out0 ? v$_5096_out0 : v$_8787_out0;
assign v$MUX5_4062_out0 = v$G6_6178_out0 ? v$_5098_out0 : v$_8789_out0;
assign v$MUX5_4063_out0 = v$G6_6179_out0 ? v$_5099_out0 : v$_8790_out0;
assign v$MUX5_4064_out0 = v$G6_6180_out0 ? v$_5100_out0 : v$_8791_out0;
assign {v$A12A_4445_out1,v$A12A_4445_out0 } = v$A11_9962_out0 + v$B11_9116_out0 + v$C10_12732_out0;
assign {v$A12A_4448_out1,v$A12A_4448_out0 } = v$A11_9965_out0 + v$B11_9119_out0 + v$C10_12735_out0;
assign v$C17_6066_out0 = v$C17_2520_out0;
assign v$C17_6069_out0 = v$C17_2523_out0;
assign v$LOWER$PART_6316_out0 = v$MUX16_16764_out0;
assign v$LOWER$PART_6317_out0 = v$MUX16_16765_out0;
assign {v$A13_7240_out1,v$A13_7240_out0 } = v$A15_17318_out0 + v$B15_10021_out0 + v$C14_279_out0;
assign {v$A13_7243_out1,v$A13_7243_out0 } = v$A15_17321_out0 + v$B15_10024_out0 + v$C14_282_out0;
assign v$SEL1_8713_out0 = v$IN_3860_out0[23:16];
assign v$SEL1_8723_out0 = v$IN_3863_out0[23:16];
assign v$C12_9394_out0 = v$C12_13520_out0;
assign v$C12_9397_out0 = v$C12_13523_out0;
assign {v$A18_10032_out1,v$A18_10032_out0 } = v$A13_13862_out0 + v$B13_8675_out0 + v$C12_13520_out0;
assign {v$A18_10035_out1,v$A18_10035_out0 } = v$A13_13865_out0 + v$B13_8678_out0 + v$C12_13523_out0;
assign v$G4_11120_out0 = v$G5_4528_out0 || v$G$CD_923_out0;
assign v$G4_11139_out0 = v$G5_4547_out0 || v$G$CD_942_out0;
assign v$G4_11243_out0 = v$G5_4651_out0 || v$G$CD_1046_out0;
assign v$G4_11262_out0 = v$G5_4670_out0 || v$G$CD_1065_out0;
assign v$G8_11411_out0 = v$CINA_8480_out0 && v$P$AB_2017_out0;
assign v$G8_11418_out0 = v$CINA_8487_out0 && v$P$AB_2024_out0;
assign v$G8_11422_out0 = v$CINA_8491_out0 && v$P$AB_2028_out0;
assign v$G8_11425_out0 = v$CINA_8494_out0 && v$P$AB_2031_out0;
assign v$G8_11433_out0 = v$CINA_8502_out0 && v$P$AB_2039_out0;
assign v$G8_11534_out0 = v$CINA_8603_out0 && v$P$AB_2140_out0;
assign v$G8_11541_out0 = v$CINA_8610_out0 && v$P$AB_2147_out0;
assign v$G8_11545_out0 = v$CINA_8614_out0 && v$P$AB_2151_out0;
assign v$G8_11548_out0 = v$CINA_8617_out0 && v$P$AB_2154_out0;
assign v$G8_11556_out0 = v$CINA_8625_out0 && v$P$AB_2162_out0;
assign v$C9_12155_out0 = v$C9_5937_out0;
assign v$C9_12158_out0 = v$C9_5940_out0;
assign {v$A15_13216_out1,v$A15_13216_out0 } = v$A18_17695_out0 + v$B18_10867_out0 + v$C17_2520_out0;
assign {v$A15_13219_out1,v$A15_13219_out0 } = v$A18_17698_out0 + v$B18_10870_out0 + v$C17_2523_out0;
assign {v$A16A_14559_out1,v$A16A_14559_out0 } = v$A10_1548_out0 + v$B10_9877_out0 + v$C9_5937_out0;
assign {v$A16A_14562_out1,v$A16A_14562_out0 } = v$A10_1551_out0 + v$B10_9880_out0 + v$C9_5940_out0;
assign v$SEL1_15404_out0 = v$IN_3860_out0[7:0];
assign v$SEL1_15414_out0 = v$IN_3863_out0[7:0];
assign v$G1_16143_out0 = v$G7_9854_out0 && v$Z4_7921_out0;
assign v$G1_16144_out0 = v$G7_9855_out0 && v$Z4_7922_out0;
assign v$G1_16145_out0 = v$G7_9856_out0 && v$Z4_7923_out0;
assign v$G1_16146_out0 = v$G7_9858_out0 && v$Z4_7924_out0;
assign v$G1_16147_out0 = v$G7_9859_out0 && v$Z4_7925_out0;
assign v$G1_16148_out0 = v$G7_9860_out0 && v$Z4_7926_out0;
assign v$C23_16149_out0 = v$C23_4843_out0;
assign v$C23_16152_out0 = v$C23_4846_out0;
assign {v$A20_16374_out1,v$A20_16374_out0 } = v$A14_676_out0 + v$B14_4002_out0 + v$C13_11776_out0;
assign {v$A20_16377_out1,v$A20_16377_out0 } = v$A14_679_out0 + v$B14_4005_out0 + v$C13_11779_out0;
assign v$C13_18589_out0 = v$C13_11776_out0;
assign v$C13_18592_out0 = v$C13_11779_out0;
assign v$MUX15_1319_out0 = v$EQ15_15967_out0 ? v$SEL15_4888_out0 : v$LOWER$PART_6316_out0;
assign v$MUX15_1320_out0 = v$EQ15_15968_out0 ? v$SEL15_4889_out0 : v$LOWER$PART_6317_out0;
assign v$ENDq_1458_out0 = v$A12A_4445_out1;
assign v$ENDq_1461_out0 = v$A12A_4448_out1;
assign v$Z_2556_out0 = v$G1_16143_out0;
assign v$Z_2557_out0 = v$G1_16144_out0;
assign v$Z_2558_out0 = v$G1_16145_out0;
assign v$Z_2560_out0 = v$G1_16146_out0;
assign v$Z_2561_out0 = v$G1_16147_out0;
assign v$Z_2562_out0 = v$G1_16148_out0;
assign v$MUX4_2874_out0 = v$G5_17509_out0 ? v$_8899_out0 : v$MUX5_4058_out0;
assign v$MUX4_2875_out0 = v$G5_17510_out0 ? v$_8900_out0 : v$MUX5_4059_out0;
assign v$MUX4_2876_out0 = v$G5_17511_out0 ? v$_8901_out0 : v$MUX5_4060_out0;
assign v$MUX4_2878_out0 = v$G5_17512_out0 ? v$_8903_out0 : v$MUX5_4062_out0;
assign v$MUX4_2879_out0 = v$G5_17513_out0 ? v$_8904_out0 : v$MUX5_4063_out0;
assign v$MUX4_2880_out0 = v$G5_17514_out0 ? v$_8905_out0 : v$MUX5_4064_out0;
assign v$_4263_out0 = { v$C2_121_out0,v$SEL1_15404_out0 };
assign v$_4273_out0 = { v$C2_131_out0,v$SEL1_15414_out0 };
assign v$_5896_out0 = { v$A17A_2487_out0,v$A18_10032_out0 };
assign v$_5899_out0 = { v$A17A_2490_out0,v$A18_10035_out0 };
assign v$CARRY_6332_out0 = v$C23_16149_out0;
assign v$CARRY_6335_out0 = v$C23_16152_out0;
assign v$ENDr_7522_out0 = v$A20_16374_out1;
assign v$ENDr_7525_out0 = v$A20_16377_out1;
assign v$_7552_out0 = { v$C8_18497_out0,v$C9_12155_out0 };
assign v$_7555_out0 = { v$C8_18500_out0,v$C9_12158_out0 };
assign v$ENDi_8682_out0 = v$A15_13216_out1;
assign v$ENDi_8685_out0 = v$A15_13219_out1;
assign v$_8998_out0 = { v$SEL1_8713_out0,v$C1_5979_out0 };
assign v$_9008_out0 = { v$SEL1_8723_out0,v$C1_5989_out0 };
assign v$END0_9352_out0 = v$A16A_14559_out1;
assign v$END0_9355_out0 = v$A16A_14562_out1;
assign v$G7_9651_out0 = v$G8_11411_out0 && v$P$CD_10470_out0;
assign v$G7_9658_out0 = v$G8_11418_out0 && v$P$CD_10477_out0;
assign v$G7_9662_out0 = v$G8_11422_out0 && v$P$CD_10481_out0;
assign v$G7_9665_out0 = v$G8_11425_out0 && v$P$CD_10484_out0;
assign v$G7_9673_out0 = v$G8_11433_out0 && v$P$CD_10492_out0;
assign v$G7_9774_out0 = v$G8_11534_out0 && v$P$CD_10593_out0;
assign v$G7_9781_out0 = v$G8_11541_out0 && v$P$CD_10600_out0;
assign v$G7_9785_out0 = v$G8_11545_out0 && v$P$CD_10604_out0;
assign v$G7_9788_out0 = v$G8_11548_out0 && v$P$CD_10607_out0;
assign v$G7_9796_out0 = v$G8_11556_out0 && v$P$CD_10615_out0;
assign v$_10237_out0 = { v$C12_9394_out0,v$C13_18589_out0 };
assign v$_10240_out0 = { v$C12_9397_out0,v$C13_18592_out0 };
assign v$ENDt_10258_out0 = v$A13_7240_out1;
assign v$ENDt_10261_out0 = v$A13_7243_out1;
assign v$_10958_out0 = { v$A16A_14559_out0,v$A12A_4445_out0 };
assign v$_10961_out0 = { v$A16A_14562_out0,v$A12A_4448_out0 };
assign v$_14836_out0 = { v$C10_1940_out0,v$C11_9510_out0 };
assign v$_14839_out0 = { v$C10_1943_out0,v$C11_9513_out0 };
assign v$G$AD_17095_out0 = v$G4_11120_out0;
assign v$G$AD_17114_out0 = v$G4_11139_out0;
assign v$G$AD_17218_out0 = v$G4_11243_out0;
assign v$G$AD_17237_out0 = v$G4_11262_out0;
assign v$_17456_out0 = { v$A20_16374_out0,v$A13_7240_out0 };
assign v$_17459_out0 = { v$A20_16377_out0,v$A13_7243_out0 };
assign v$ENDe_17892_out0 = v$A18_10032_out1;
assign v$ENDe_17895_out0 = v$A18_10035_out1;
assign v$G6_449_out0 = v$G4_11127_out0 || v$G7_9651_out0;
assign v$G6_456_out0 = v$G4_11134_out0 || v$G7_9658_out0;
assign v$G6_460_out0 = v$G4_11138_out0 || v$G7_9662_out0;
assign v$G6_463_out0 = v$G4_11141_out0 || v$G7_9665_out0;
assign v$G6_471_out0 = v$G4_11149_out0 || v$G7_9673_out0;
assign v$G6_572_out0 = v$G4_11250_out0 || v$G7_9774_out0;
assign v$G6_579_out0 = v$G4_11257_out0 || v$G7_9781_out0;
assign v$G6_583_out0 = v$G4_11261_out0 || v$G7_9785_out0;
assign v$G6_586_out0 = v$G4_11264_out0 || v$G7_9788_out0;
assign v$G6_594_out0 = v$G4_11272_out0 || v$G7_9796_out0;
assign v$_1557_out0 = { v$_15013_out0,v$_10958_out0 };
assign v$_1560_out0 = { v$_15016_out0,v$_10961_out0 };
assign v$MUX1_2367_out0 = v$LEFT$SHIT_3059_out0 ? v$_4263_out0 : v$_8998_out0;
assign v$MUX1_2377_out0 = v$LEFT$SHIT_3069_out0 ? v$_4273_out0 : v$_9008_out0;
assign v$TWOS$COMPLEMENT$ADDER$COUT_3431_out0 = v$CARRY_6332_out0;
assign v$TWOS$COMPLEMENT$ADDER$COUT_3432_out0 = v$CARRY_6335_out0;
assign v$MUX14_4921_out0 = v$EQ14_5403_out0 ? v$SEL14_16349_out0 : v$MUX15_1319_out0;
assign v$MUX14_4922_out0 = v$EQ14_5404_out0 ? v$SEL14_16350_out0 : v$MUX15_1320_out0;
assign v$Z2_6324_out0 = v$Z_2557_out0;
assign v$Z2_6328_out0 = v$Z_2561_out0;
assign v$END50_7413_out0 = v$G$AD_17095_out0;
assign v$END50_7416_out0 = v$G$AD_17218_out0;
assign v$END48_10365_out0 = v$G$AD_17114_out0;
assign v$END48_10368_out0 = v$G$AD_17237_out0;
assign v$_14293_out0 = { v$_5896_out0,v$_17456_out0 };
assign v$_14296_out0 = { v$_5899_out0,v$_17459_out0 };
assign v$Z1_16998_out0 = v$Z_2556_out0;
assign v$Z1_17002_out0 = v$Z_2560_out0;
assign v$MUX3_17472_out0 = v$G4_6055_out0 ? v$_3979_out0 : v$MUX4_2874_out0;
assign v$MUX3_17473_out0 = v$G4_6056_out0 ? v$_3980_out0 : v$MUX4_2875_out0;
assign v$MUX3_17474_out0 = v$G4_6057_out0 ? v$_3981_out0 : v$MUX4_2876_out0;
assign v$MUX3_17475_out0 = v$G4_6058_out0 ? v$_3982_out0 : v$MUX4_2878_out0;
assign v$MUX3_17476_out0 = v$G4_6059_out0 ? v$_3983_out0 : v$MUX4_2879_out0;
assign v$MUX3_17477_out0 = v$G4_6060_out0 ? v$_3984_out0 : v$MUX4_2880_out0;
assign v$Z3_17779_out0 = v$Z_2558_out0;
assign v$Z3_17783_out0 = v$Z_2562_out0;
assign v$_18303_out0 = { v$_7552_out0,v$_14836_out0 };
assign v$_18306_out0 = { v$_7555_out0,v$_14839_out0 };
assign v$_1173_out0 = { v$_1557_out0,v$_14293_out0 };
assign v$_1176_out0 = { v$_1560_out0,v$_14296_out0 };
assign v$G6_6173_out0 = ! v$Z2_6324_out0;
assign v$G6_6177_out0 = ! v$Z2_6328_out0;
assign v$COUTD_6709_out0 = v$G6_449_out0;
assign v$COUTD_6716_out0 = v$G6_456_out0;
assign v$COUTD_6720_out0 = v$G6_460_out0;
assign v$COUTD_6723_out0 = v$G6_463_out0;
assign v$COUTD_6731_out0 = v$G6_471_out0;
assign v$COUTD_6832_out0 = v$G6_572_out0;
assign v$COUTD_6839_out0 = v$G6_579_out0;
assign v$COUTD_6843_out0 = v$G6_583_out0;
assign v$COUTD_6846_out0 = v$G6_586_out0;
assign v$COUTD_6854_out0 = v$G6_594_out0;
assign v$OUT_8956_out0 = v$MUX3_17472_out0;
assign v$OUT_8957_out0 = v$MUX3_17473_out0;
assign v$OUT_8958_out0 = v$MUX3_17474_out0;
assign v$OUT_8960_out0 = v$MUX3_17475_out0;
assign v$OUT_8961_out0 = v$MUX3_17476_out0;
assign v$OUT_8962_out0 = v$MUX3_17477_out0;
assign v$MUX13_13684_out0 = v$EQ13_9517_out0 ? v$SEL13_6926_out0 : v$MUX14_4921_out0;
assign v$MUX13_13685_out0 = v$EQ13_9518_out0 ? v$SEL13_6927_out0 : v$MUX14_4922_out0;
assign v$G9_15202_out0 = v$Z1_16998_out0 && v$Z2_6324_out0;
assign v$G9_15206_out0 = v$Z1_17002_out0 && v$Z2_6328_out0;
assign v$G10_16091_out0 = ! v$Z3_17779_out0;
assign v$G10_16092_out0 = ! v$Z3_17783_out0;
assign v$MUX2_18576_out0 = v$EN_5213_out0 ? v$MUX1_2367_out0 : v$IN_3860_out0;
assign v$MUX2_18578_out0 = v$EN_5215_out0 ? v$MUX1_2377_out0 : v$IN_3863_out0;
assign v$C16_1268_out0 = v$COUTD_6723_out0;
assign v$C16_1271_out0 = v$COUTD_6846_out0;
assign v$_5093_out0 = { v$OUT_8957_out0,v$C5_16912_out0 };
assign v$_5097_out0 = { v$OUT_8961_out0,v$C5_16916_out0 };
assign v$C15_8143_out0 = v$COUTD_6720_out0;
assign v$C15_8146_out0 = v$COUTD_6843_out0;
assign v$C19_8160_out0 = v$COUTD_6731_out0;
assign v$C19_8163_out0 = v$COUTD_6854_out0;
assign v$CINA_8473_out0 = v$COUTD_6716_out0;
assign v$CINA_8492_out0 = v$COUTD_6716_out0;
assign v$CINA_8596_out0 = v$COUTD_6839_out0;
assign v$CINA_8615_out0 = v$COUTD_6839_out0;
assign v$_8784_out0 = { v$OUT_8956_out0,v$C6_6538_out0 };
assign v$_8788_out0 = { v$OUT_8960_out0,v$C6_6542_out0 };
assign v$_8898_out0 = { v$OUT_8958_out0,v$C4_16511_out0 };
assign v$_8902_out0 = { v$OUT_8962_out0,v$C4_16515_out0 };
assign v$G7_9853_out0 = v$G9_15202_out0 && v$Z3_17779_out0;
assign v$G7_9857_out0 = v$G9_15206_out0 && v$Z3_17783_out0;
assign v$OUT_14919_out0 = v$MUX2_18576_out0;
assign v$OUT_14929_out0 = v$MUX2_18578_out0;
assign v$C20_15489_out0 = v$COUTD_6716_out0;
assign v$C20_15492_out0 = v$COUTD_6839_out0;
assign v$C18_16289_out0 = v$COUTD_6709_out0;
assign v$C18_16292_out0 = v$COUTD_6832_out0;
assign v$MUX12_17815_out0 = v$EQ12_13840_out0 ? v$SEL12_13846_out0 : v$MUX13_13684_out0;
assign v$MUX12_17816_out0 = v$EQ12_13841_out0 ? v$SEL12_13847_out0 : v$MUX13_13685_out0;
assign v$_18233_out0 = { v$_17748_out0,v$_1173_out0 };
assign v$_18236_out0 = { v$_17751_out0,v$_1176_out0 };
assign v$Z_2555_out0 = v$G7_9853_out0;
assign v$Z_2559_out0 = v$G7_9857_out0;
assign v$MUX5_4057_out0 = v$G6_6173_out0 ? v$_5093_out0 : v$_8784_out0;
assign v$MUX5_4061_out0 = v$G6_6177_out0 ? v$_5097_out0 : v$_8788_out0;
assign v$OUT_4913_out0 = v$OUT_14919_out0;
assign v$OUT_4914_out0 = v$OUT_14929_out0;
assign v$G8_11404_out0 = v$CINA_8473_out0 && v$P$AB_2010_out0;
assign v$G8_11423_out0 = v$CINA_8492_out0 && v$P$AB_2029_out0;
assign v$G8_11527_out0 = v$CINA_8596_out0 && v$P$AB_2133_out0;
assign v$G8_11546_out0 = v$CINA_8615_out0 && v$P$AB_2152_out0;
assign v$C15_13131_out0 = v$C15_8143_out0;
assign v$C15_13134_out0 = v$C15_8146_out0;
assign v$C19_13833_out0 = v$C19_8160_out0;
assign v$C19_13836_out0 = v$C19_8163_out0;
assign v$C20_14978_out0 = v$C20_15489_out0;
assign v$C20_14981_out0 = v$C20_15492_out0;
assign v$C16_15157_out0 = v$C16_1268_out0;
assign v$C16_15160_out0 = v$C16_1271_out0;
assign {v$A14_15353_out1,v$A14_15353_out0 } = v$A16_13614_out0 + v$B16_16414_out0 + v$C15_8143_out0;
assign {v$A14_15356_out1,v$A14_15356_out0 } = v$A16_13617_out0 + v$B16_16417_out0 + v$C15_8146_out0;
assign {v$A19_15908_out1,v$A19_15908_out0 } = v$A19_1213_out0 + v$B19_16789_out0 + v$C18_16289_out0;
assign {v$A19_15911_out1,v$A19_15911_out0 } = v$A19_1216_out0 + v$B19_16792_out0 + v$C18_16292_out0;
assign {v$A24_16973_out1,v$A24_16973_out0 } = v$A21_2598_out0 + v$B21_18082_out0 + v$C20_15489_out0;
assign {v$A24_16976_out1,v$A24_16976_out0 } = v$A21_2601_out0 + v$B21_18085_out0 + v$C20_15492_out0;
assign {v$A22_17488_out1,v$A22_17488_out0 } = v$A20_4436_out0 + v$B20_3943_out0 + v$C19_8160_out0;
assign {v$A22_17491_out1,v$A22_17491_out0 } = v$A20_4439_out0 + v$B20_3946_out0 + v$C19_8163_out0;
assign {v$A11_17874_out1,v$A11_17874_out0 } = v$A17_16722_out0 + v$B17_15535_out0 + v$C16_1268_out0;
assign {v$A11_17877_out1,v$A11_17877_out0 } = v$A17_16725_out0 + v$B17_15538_out0 + v$C16_1271_out0;
assign v$MUX11_17935_out0 = v$EQ11_6145_out0 ? v$SEL11_7227_out0 : v$MUX12_17815_out0;
assign v$MUX11_17936_out0 = v$EQ11_6146_out0 ? v$SEL11_7228_out0 : v$MUX12_17816_out0;
assign v$C18_18005_out0 = v$C18_16289_out0;
assign v$C18_18008_out0 = v$C18_16292_out0;
assign v$_1199_out0 = { v$A15_13216_out0,v$A19_15908_out0 };
assign v$_1202_out0 = { v$A15_13219_out0,v$A19_15911_out0 };
assign v$_1793_out0 = { v$A22_17488_out0,v$A24_16973_out0 };
assign v$_1796_out0 = { v$A22_17491_out0,v$A24_16976_out0 };
assign v$_2840_out0 = { v$C14_325_out0,v$C15_13131_out0 };
assign v$_2843_out0 = { v$C14_328_out0,v$C15_13134_out0 };
assign v$MUX4_2873_out0 = v$G10_16091_out0 ? v$_8898_out0 : v$MUX5_4057_out0;
assign v$MUX4_2877_out0 = v$G10_16092_out0 ? v$_8902_out0 : v$MUX5_4061_out0;
assign v$MUX8_2947_out0 = v$EQ9_13777_out0 ? v$SEL9_10265_out0 : v$MUX11_17935_out0;
assign v$MUX8_2948_out0 = v$EQ9_13778_out0 ? v$SEL9_10266_out0 : v$MUX11_17936_out0;
assign v$ENDp_3189_out0 = v$A22_17488_out1;
assign v$ENDp_3192_out0 = v$A22_17491_out1;
assign v$ENDy_4114_out0 = v$A14_15353_out1;
assign v$ENDy_4117_out0 = v$A14_15356_out1;
assign v$SEL1_6028_out0 = v$OUT_4914_out0[22:0];
assign v$ENDu_7029_out0 = v$A11_17874_out1;
assign v$ENDu_7032_out0 = v$A11_17877_out1;
assign v$_7868_out0 = { v$C16_15157_out0,v$C17_6066_out0 };
assign v$_7871_out0 = { v$C16_15160_out0,v$C17_6069_out0 };
assign v$SEL2_8098_out0 = v$OUT_4913_out0[22:13];
assign v$_8329_out0 = { v$C18_18005_out0,v$C19_13833_out0 };
assign v$_8332_out0 = { v$C18_18008_out0,v$C19_13836_out0 };
assign v$G7_9644_out0 = v$G8_11404_out0 && v$P$CD_10463_out0;
assign v$G7_9663_out0 = v$G8_11423_out0 && v$P$CD_10482_out0;
assign v$G7_9767_out0 = v$G8_11527_out0 && v$P$CD_10586_out0;
assign v$G7_9786_out0 = v$G8_11546_out0 && v$P$CD_10605_out0;
assign v$_13293_out0 = { v$A14_15353_out0,v$A11_17874_out0 };
assign v$_13296_out0 = { v$A14_15356_out0,v$A11_17877_out0 };
assign v$Z_15810_out0 = v$Z_2555_out0;
assign v$Z_15811_out0 = v$Z_2559_out0;
assign v$ENDa_16564_out0 = v$A24_16973_out1;
assign v$ENDa_16567_out0 = v$A24_16976_out1;
assign v$ENDo_18692_out0 = v$A19_15908_out1;
assign v$ENDo_18695_out0 = v$A19_15911_out1;
assign v$G6_442_out0 = v$G4_11120_out0 || v$G7_9644_out0;
assign v$G6_461_out0 = v$G4_11139_out0 || v$G7_9663_out0;
assign v$G6_565_out0 = v$G4_11243_out0 || v$G7_9767_out0;
assign v$G6_584_out0 = v$G4_11262_out0 || v$G7_9786_out0;
assign v$_1242_out0 = { v$_10237_out0,v$_2840_out0 };
assign v$_1245_out0 = { v$_10240_out0,v$_2843_out0 };
assign v$OUT_8955_out0 = v$MUX4_2873_out0;
assign v$OUT_8959_out0 = v$MUX4_2877_out0;
assign v$_10349_out0 = { v$_7868_out0,v$_8329_out0 };
assign v$_10352_out0 = { v$_7871_out0,v$_8332_out0 };
assign v$MUX10_15674_out0 = v$EQ10_5894_out0 ? v$SEL8_17685_out0 : v$MUX8_2947_out0;
assign v$MUX10_15675_out0 = v$EQ10_5895_out0 ? v$SEL8_17686_out0 : v$MUX8_2948_out0;
assign v$_15846_out0 = { v$SEL2_8098_out0,v$A2_10044_out0 };
assign v$_15847_out0 = { v$SEL1_6028_out0,v$A2_10045_out0 };
assign v$_16256_out0 = { v$_13293_out0,v$_1199_out0 };
assign v$_16259_out0 = { v$_13296_out0,v$_1202_out0 };
assign v$COUTD_6702_out0 = v$G6_442_out0;
assign v$COUTD_6721_out0 = v$G6_461_out0;
assign v$COUTD_6825_out0 = v$G6_565_out0;
assign v$COUTD_6844_out0 = v$G6_584_out0;
assign v$MUX9_8245_out0 = v$EQ8_14416_out0 ? v$SEL10_9508_out0 : v$MUX10_15674_out0;
assign v$MUX9_8246_out0 = v$EQ8_14417_out0 ? v$SEL10_9509_out0 : v$MUX10_15675_out0;
assign v$AMOUNT$OF$SHIFT_9461_out0 = v$OUT_8955_out0;
assign v$AMOUNT$OF$SHIFT_9462_out0 = v$OUT_8959_out0;
assign v$MUX2_13630_out0 = v$Z_15808_out0 ? v$C4_8256_out0 : v$_15846_out0;
assign v$MUX2_13631_out0 = v$Z_15809_out0 ? v$C4_8257_out0 : v$_15847_out0;
assign v$_17353_out0 = { v$_18303_out0,v$_1242_out0 };
assign v$_17356_out0 = { v$_18306_out0,v$_1245_out0 };
assign v$MUX7_1229_out0 = v$EQ7_4087_out0 ? v$SEL7_14334_out0 : v$MUX9_8245_out0;
assign v$MUX7_1230_out0 = v$EQ7_4088_out0 ? v$SEL7_14335_out0 : v$MUX9_8246_out0;
assign v$SEL4_1847_out0 = v$AMOUNT$OF$SHIFT_9461_out0[3:3];
assign v$SEL4_1848_out0 = v$AMOUNT$OF$SHIFT_9462_out0[3:3];
assign v$_4867_out0 = { v$_7790_out0,v$_17353_out0 };
assign v$_4870_out0 = { v$_7793_out0,v$_17356_out0 };
assign v$SEL6_8932_out0 = v$AMOUNT$OF$SHIFT_9461_out0[5:5];
assign v$SEL6_8933_out0 = v$AMOUNT$OF$SHIFT_9462_out0[5:5];
assign v$C21_10767_out0 = v$COUTD_6721_out0;
assign v$C21_10770_out0 = v$COUTD_6844_out0;
assign v$C22_10981_out0 = v$COUTD_6702_out0;
assign v$C22_10984_out0 = v$COUTD_6825_out0;
assign v$SEL5_11669_out0 = v$AMOUNT$OF$SHIFT_9461_out0[4:4];
assign v$SEL5_11670_out0 = v$AMOUNT$OF$SHIFT_9462_out0[4:4];
assign v$SEL1_13357_out0 = v$AMOUNT$OF$SHIFT_9461_out0[0:0];
assign v$SEL1_13358_out0 = v$AMOUNT$OF$SHIFT_9462_out0[0:0];
assign v$SEL3_14008_out0 = v$AMOUNT$OF$SHIFT_9461_out0[2:2];
assign v$SEL3_14009_out0 = v$AMOUNT$OF$SHIFT_9462_out0[2:2];
assign v$_18416_out0 = { v$MUX2_13630_out0,v$SIGN_1366_out0 };
assign v$_18417_out0 = { v$MUX2_13631_out0,v$SIGN_1367_out0 };
assign v$SEL2_18504_out0 = v$AMOUNT$OF$SHIFT_9461_out0[1:1];
assign v$SEL2_18505_out0 = v$AMOUNT$OF$SHIFT_9462_out0[1:1];
assign v$EN_1343_out0 = v$SEL4_1847_out0;
assign v$EN_1344_out0 = v$SEL4_1848_out0;
assign v$EN_4758_out0 = v$SEL3_14008_out0;
assign v$EN_4759_out0 = v$SEL3_14009_out0;
assign v$EN_5217_out0 = v$SEL6_8932_out0;
assign v$EN_5218_out0 = v$SEL5_11669_out0;
assign v$EN_5219_out0 = v$SEL1_13357_out0;
assign v$EN_5220_out0 = v$SEL6_8933_out0;
assign v$EN_5221_out0 = v$SEL5_11670_out0;
assign v$EN_5222_out0 = v$SEL1_13358_out0;
assign v$C21_6369_out0 = v$C21_10767_out0;
assign v$C21_6372_out0 = v$C21_10770_out0;
assign v$EN_7880_out0 = v$SEL2_18504_out0;
assign v$EN_7881_out0 = v$SEL2_18505_out0;
assign v$C22_8410_out0 = v$C22_10981_out0;
assign v$C22_8413_out0 = v$C22_10984_out0;
assign {v$A23_9546_out1,v$A23_9546_out0 } = v$A23_5063_out0 + v$B23_1283_out0 + v$C22_10981_out0;
assign {v$A23_9549_out1,v$A23_9549_out0 } = v$A23_5066_out0 + v$B23_1286_out0 + v$C22_10984_out0;
assign v$OUT_12478_out0 = v$_18416_out0;
assign v$OUT_12479_out0 = v$_18417_out0;
assign v$MUX6_16287_out0 = v$EQ6_5427_out0 ? v$SEL6_12474_out0 : v$MUX7_1229_out0;
assign v$MUX6_16288_out0 = v$EQ6_5428_out0 ? v$SEL6_12475_out0 : v$MUX7_1230_out0;
assign {v$A21_18568_out1,v$A21_18568_out0 } = v$A22_4424_out0 + v$B22_10805_out0 + v$C21_10767_out0;
assign {v$A21_18571_out1,v$A21_18571_out0 } = v$A22_4427_out0 + v$B22_10808_out0 + v$C21_10770_out0;
assign v$_650_out0 = { v$C20_14978_out0,v$C21_6369_out0 };
assign v$_653_out0 = { v$C20_14981_out0,v$C21_6372_out0 };
assign v$_1576_out0 = { v$A21_18568_out0,v$A23_9546_out0 };
assign v$_1579_out0 = { v$A21_18571_out0,v$A23_9549_out0 };
assign v$ENDs_3213_out0 = v$A21_18568_out1;
assign v$ENDs_3216_out0 = v$A21_18571_out1;
assign v$MUX5_6930_out0 = v$EQ5_3317_out0 ? v$SEL5_15453_out0 : v$MUX6_16287_out0;
assign v$MUX5_6931_out0 = v$EQ5_3318_out0 ? v$SEL5_15454_out0 : v$MUX6_16288_out0;
assign v$MUX11_8669_out0 = v$G5_6198_out0 ? v$C9_18760_out0 : v$OUT_12478_out0;
assign v$MUX3_8965_out0 = v$G3_16009_out0 ? v$C1_15226_out0 : v$OUT_12479_out0;
assign v$ENDd_10832_out0 = v$A23_9546_out1;
assign v$ENDd_10835_out0 = v$A23_9549_out1;
assign v$_15708_out0 = { v$C22_8410_out0,v$C23_16149_out0 };
assign v$_15711_out0 = { v$C22_8413_out0,v$C23_16152_out0 };
assign v$MUX2_18582_out0 = v$EN_5219_out0 ? v$MUX1_2389_out0 : v$IN_3868_out0;
assign v$MUX2_18585_out0 = v$EN_5222_out0 ? v$MUX1_2395_out0 : v$IN_3871_out0;
assign v$MUX4_7801_out0 = v$EQ4_18601_out0 ? v$SEL4_7323_out0 : v$MUX5_6930_out0;
assign v$MUX4_7802_out0 = v$EQ4_18602_out0 ? v$SEL4_7324_out0 : v$MUX5_6931_out0;
assign v$SINGLE$PRECISION_7900_out0 = v$MUX3_8965_out0;
assign v$_9491_out0 = { v$_1793_out0,v$_1576_out0 };
assign v$_9494_out0 = { v$_1796_out0,v$_1579_out0 };
assign v$_13732_out0 = { v$_650_out0,v$_15708_out0 };
assign v$_13735_out0 = { v$_653_out0,v$_15711_out0 };
assign v$OUT_14941_out0 = v$MUX2_18582_out0;
assign v$OUT_14947_out0 = v$MUX2_18585_out0;
assign v$_17036_out0 = { v$C10_6384_out0,v$MUX11_8669_out0 };
assign v$_4092_out0 = { v$_10349_out0,v$_13732_out0 };
assign v$_4095_out0 = { v$_10352_out0,v$_13735_out0 };
assign v$IN_5185_out0 = v$OUT_14941_out0;
assign v$IN_5191_out0 = v$OUT_14947_out0;
assign v$_6658_out0 = { v$_16256_out0,v$_9491_out0 };
assign v$_6661_out0 = { v$_16259_out0,v$_9494_out0 };
assign v$MUX3_7602_out0 = v$EQ3_1818_out0 ? v$SEL3_11731_out0 : v$MUX4_7801_out0;
assign v$MUX3_7603_out0 = v$EQ3_1819_out0 ? v$SEL3_11732_out0 : v$MUX4_7802_out0;
assign v$HALF$PRECISION_10311_out0 = v$_17036_out0;
assign v$_3759_out0 = { v$_4867_out0,v$_4092_out0 };
assign v$_3762_out0 = { v$_4870_out0,v$_4095_out0 };
assign v$_9906_out0 = { v$_18233_out0,v$_6658_out0 };
assign v$_9909_out0 = { v$_18236_out0,v$_6661_out0 };
assign v$IN_11788_out0 = v$IN_5185_out0;
assign v$IN_11789_out0 = v$IN_5191_out0;
assign v$MUX2_13610_out0 = v$EQ2_14210_out0 ? v$SEL2_13323_out0 : v$MUX3_7602_out0;
assign v$MUX2_13611_out0 = v$EQ2_14211_out0 ? v$SEL2_13324_out0 : v$MUX3_7603_out0;
assign v$MUX12_16796_out0 = v$IS$32$BITS_2992_out0 ? v$SINGLE$PRECISION_7900_out0 : v$HALF$PRECISION_10311_out0;
assign v$MUX1_2867_out0 = v$EQ1_13416_out0 ? v$SEL1_7090_out0 : v$MUX2_13610_out0;
assign v$MUX1_2868_out0 = v$EQ1_13417_out0 ? v$SEL1_7091_out0 : v$MUX2_13611_out0;
assign v$OUT_3364_out0 = v$MUX12_16796_out0;
assign v$SEL1_8733_out0 = v$IN_11788_out0[47:2];
assign v$SEL1_8739_out0 = v$IN_11789_out0[47:2];
assign v$SUM_9362_out0 = v$_9906_out0;
assign v$SUM_9365_out0 = v$_9909_out0;
assign v$SUM1_12827_out0 = v$_3759_out0;
assign v$SUM1_12830_out0 = v$_3762_out0;
assign v$SEL1_15424_out0 = v$IN_11788_out0[45:0];
assign v$SEL1_15430_out0 = v$IN_11789_out0[45:0];
assign v$END_1870_out0 = v$SUM1_12827_out0;
assign v$END_1871_out0 = v$SUM1_12830_out0;
assign v$_4283_out0 = { v$C2_141_out0,v$SEL1_15424_out0 };
assign v$_4289_out0 = { v$C2_147_out0,v$SEL1_15430_out0 };
assign v$MUX5_6222_out0 = v$IS$A$LARGER_10444_out0 ? v$SUM_1905_out0 : v$SUM_9362_out0;
assign v$MUX5_6223_out0 = v$IS$A$LARGER_10445_out0 ? v$SUM_1906_out0 : v$SUM_9365_out0;
assign v$MUX25_8406_out0 = v$G2_11904_out0 ? v$C2_15180_out0 : v$MUX1_2867_out0;
assign v$MUX25_8407_out0 = v$G2_11905_out0 ? v$C2_15181_out0 : v$MUX1_2868_out0;
assign v$_9018_out0 = { v$SEL1_8733_out0,v$C1_5999_out0 };
assign v$_9024_out0 = { v$SEL1_8739_out0,v$C1_6005_out0 };
assign v$MUX1_2387_out0 = v$LEFT$SHIT_3079_out0 ? v$_4283_out0 : v$_9018_out0;
assign v$MUX1_2393_out0 = v$LEFT$SHIT_3085_out0 ? v$_4289_out0 : v$_9024_out0;
assign v$LZD$INPUT_8837_out0 = v$MUX5_6222_out0;
assign v$LZD$INPUT_8838_out0 = v$MUX5_6223_out0;
assign v$OUT_9478_out0 = v$MUX25_8406_out0;
assign v$OUT_9479_out0 = v$MUX25_8407_out0;
assign v$MUX2_2482_out0 = v$EN_7880_out0 ? v$MUX1_2387_out0 : v$IN_11788_out0;
assign v$MUX2_2483_out0 = v$EN_7881_out0 ? v$MUX1_2393_out0 : v$IN_11789_out0;
assign {v$A1_2664_out1,v$A1_2664_out0 } = v$LARGER$EXP_10276_out0 + v$SMALLER$EXP_2943_out0 + v$OUT_9478_out0;
assign {v$A1_2665_out1,v$A1_2665_out0 } = v$LARGER$EXP_10277_out0 + v$SMALLER$EXP_2944_out0 + v$OUT_9479_out0;
assign v$IN_13167_out0 = v$LZD$INPUT_8837_out0;
assign v$IN_13172_out0 = v$LZD$INPUT_8838_out0;
assign v$IN_17987_out0 = v$LZD$INPUT_8837_out0;
assign v$IN_17988_out0 = v$LZD$INPUT_8838_out0;
assign v$SEL1_351_out0 = v$IN_17987_out0[23:16];
assign v$SEL1_352_out0 = v$IN_17988_out0[23:16];
assign v$IN_5159_out0 = v$IN_13167_out0;
assign v$IN_5207_out0 = v$IN_13172_out0;
assign {v$A2_10046_out1,v$A2_10046_out0 } = v$A1_2664_out0 + v$C1_5957_out0 + v$C2_16283_out0;
assign {v$A2_10047_out1,v$A2_10047_out0 } = v$A1_2665_out0 + v$C1_5958_out0 + v$C2_16284_out0;
assign v$OUT_14939_out0 = v$MUX2_2482_out0;
assign v$OUT_14945_out0 = v$MUX2_2483_out0;
assign v$SEL2_17370_out0 = v$IN_17987_out0[15:8];
assign v$SEL2_17371_out0 = v$IN_17988_out0[15:8];
assign v$SEL1_17423_out0 = v$IN_17987_out0[7:0];
assign v$SEL1_17424_out0 = v$IN_17988_out0[7:0];
assign v$NOT$USED$CARRY_18777_out0 = v$A1_2664_out1;
assign v$NOT$USED$CARRY_18778_out0 = v$A1_2665_out1;
assign v$IN_3858_out0 = v$IN_5159_out0;
assign v$IN_3874_out0 = v$IN_5207_out0;
assign v$IN_5188_out0 = v$OUT_14939_out0;
assign v$IN_5194_out0 = v$OUT_14945_out0;
assign v$IN_14854_out0 = v$SEL1_351_out0;
assign v$IN_14855_out0 = v$SEL2_17370_out0;
assign v$IN_14856_out0 = v$SEL1_17423_out0;
assign v$IN_14859_out0 = v$SEL1_352_out0;
assign v$IN_14860_out0 = v$SEL2_17371_out0;
assign v$IN_14861_out0 = v$SEL1_17424_out0;
assign v$NOT$USED_15952_out0 = v$A2_10046_out1;
assign v$NOT$USED_15953_out0 = v$A2_10047_out1;
assign v$SEL2_3024_out0 = v$IN_14854_out0[7:4];
assign v$SEL2_3025_out0 = v$IN_14855_out0[7:4];
assign v$SEL2_3026_out0 = v$IN_14856_out0[7:4];
assign v$SEL2_3029_out0 = v$IN_14859_out0[7:4];
assign v$SEL2_3030_out0 = v$IN_14860_out0[7:4];
assign v$SEL2_3031_out0 = v$IN_14861_out0[7:4];
assign v$SEL1_8707_out0 = v$IN_3858_out0[23:1];
assign v$SEL1_8755_out0 = v$IN_3874_out0[23:1];
assign v$SEL1_15398_out0 = v$IN_3858_out0[22:0];
assign v$SEL1_15446_out0 = v$IN_3874_out0[22:0];
assign v$IN_15610_out0 = v$IN_5188_out0;
assign v$IN_15611_out0 = v$IN_5194_out0;
assign v$SEL1_16455_out0 = v$IN_14854_out0[3:0];
assign v$SEL1_16456_out0 = v$IN_14855_out0[3:0];
assign v$SEL1_16457_out0 = v$IN_14856_out0[3:0];
assign v$SEL1_16460_out0 = v$IN_14859_out0[3:0];
assign v$SEL1_16461_out0 = v$IN_14860_out0[3:0];
assign v$SEL1_16462_out0 = v$IN_14861_out0[3:0];
assign v$_4257_out0 = { v$C2_115_out0,v$SEL1_15398_out0 };
assign v$_4305_out0 = { v$C2_163_out0,v$SEL1_15446_out0 };
assign v$SEL1_8736_out0 = v$IN_15610_out0[47:4];
assign v$SEL1_8742_out0 = v$IN_15611_out0[47:4];
assign v$_8992_out0 = { v$SEL1_8707_out0,v$C1_5973_out0 };
assign v$_9040_out0 = { v$SEL1_8755_out0,v$C1_6021_out0 };
assign v$IN_15057_out0 = v$SEL1_16455_out0;
assign v$IN_15058_out0 = v$SEL2_3024_out0;
assign v$IN_15059_out0 = v$SEL1_16456_out0;
assign v$IN_15060_out0 = v$SEL2_3025_out0;
assign v$IN_15061_out0 = v$SEL1_16457_out0;
assign v$IN_15062_out0 = v$SEL2_3026_out0;
assign v$IN_15099_out0 = v$SEL1_16460_out0;
assign v$IN_15100_out0 = v$SEL2_3029_out0;
assign v$IN_15101_out0 = v$SEL1_16461_out0;
assign v$IN_15102_out0 = v$SEL2_3030_out0;
assign v$IN_15103_out0 = v$SEL1_16462_out0;
assign v$IN_15104_out0 = v$SEL2_3031_out0;
assign v$SEL1_15427_out0 = v$IN_15610_out0[43:0];
assign v$SEL1_15433_out0 = v$IN_15611_out0[43:0];
assign v$SEL3_2294_out0 = v$IN_15057_out0[2:2];
assign v$SEL3_2295_out0 = v$IN_15058_out0[2:2];
assign v$SEL3_2296_out0 = v$IN_15059_out0[2:2];
assign v$SEL3_2297_out0 = v$IN_15060_out0[2:2];
assign v$SEL3_2298_out0 = v$IN_15061_out0[2:2];
assign v$SEL3_2299_out0 = v$IN_15062_out0[2:2];
assign v$SEL3_2336_out0 = v$IN_15099_out0[2:2];
assign v$SEL3_2337_out0 = v$IN_15100_out0[2:2];
assign v$SEL3_2338_out0 = v$IN_15101_out0[2:2];
assign v$SEL3_2339_out0 = v$IN_15102_out0[2:2];
assign v$SEL3_2340_out0 = v$IN_15103_out0[2:2];
assign v$SEL3_2341_out0 = v$IN_15104_out0[2:2];
assign v$MUX1_2361_out0 = v$LEFT$SHIT_3053_out0 ? v$_4257_out0 : v$_8992_out0;
assign v$MUX1_2409_out0 = v$LEFT$SHIT_3101_out0 ? v$_4305_out0 : v$_9040_out0;
assign v$_4286_out0 = { v$C2_144_out0,v$SEL1_15427_out0 };
assign v$_4292_out0 = { v$C2_150_out0,v$SEL1_15433_out0 };
assign v$SEL4_6079_out0 = v$IN_15057_out0[3:3];
assign v$SEL4_6080_out0 = v$IN_15058_out0[3:3];
assign v$SEL4_6081_out0 = v$IN_15059_out0[3:3];
assign v$SEL4_6082_out0 = v$IN_15060_out0[3:3];
assign v$SEL4_6083_out0 = v$IN_15061_out0[3:3];
assign v$SEL4_6084_out0 = v$IN_15062_out0[3:3];
assign v$SEL4_6121_out0 = v$IN_15099_out0[3:3];
assign v$SEL4_6122_out0 = v$IN_15100_out0[3:3];
assign v$SEL4_6123_out0 = v$IN_15101_out0[3:3];
assign v$SEL4_6124_out0 = v$IN_15102_out0[3:3];
assign v$SEL4_6125_out0 = v$IN_15103_out0[3:3];
assign v$SEL4_6126_out0 = v$IN_15104_out0[3:3];
assign v$SEL2_7670_out0 = v$IN_15057_out0[1:1];
assign v$SEL2_7671_out0 = v$IN_15058_out0[1:1];
assign v$SEL2_7672_out0 = v$IN_15059_out0[1:1];
assign v$SEL2_7673_out0 = v$IN_15060_out0[1:1];
assign v$SEL2_7674_out0 = v$IN_15061_out0[1:1];
assign v$SEL2_7675_out0 = v$IN_15062_out0[1:1];
assign v$SEL2_7712_out0 = v$IN_15099_out0[1:1];
assign v$SEL2_7713_out0 = v$IN_15100_out0[1:1];
assign v$SEL2_7714_out0 = v$IN_15101_out0[1:1];
assign v$SEL2_7715_out0 = v$IN_15102_out0[1:1];
assign v$SEL2_7716_out0 = v$IN_15103_out0[1:1];
assign v$SEL2_7717_out0 = v$IN_15104_out0[1:1];
assign v$_9021_out0 = { v$SEL1_8736_out0,v$C1_6002_out0 };
assign v$_9027_out0 = { v$SEL1_8742_out0,v$C1_6008_out0 };
assign v$SEL1_13459_out0 = v$IN_15057_out0[0:0];
assign v$SEL1_13460_out0 = v$IN_15058_out0[0:0];
assign v$SEL1_13461_out0 = v$IN_15059_out0[0:0];
assign v$SEL1_13462_out0 = v$IN_15060_out0[0:0];
assign v$SEL1_13463_out0 = v$IN_15061_out0[0:0];
assign v$SEL1_13464_out0 = v$IN_15062_out0[0:0];
assign v$SEL1_13501_out0 = v$IN_15099_out0[0:0];
assign v$SEL1_13502_out0 = v$IN_15100_out0[0:0];
assign v$SEL1_13503_out0 = v$IN_15101_out0[0:0];
assign v$SEL1_13504_out0 = v$IN_15102_out0[0:0];
assign v$SEL1_13505_out0 = v$IN_15103_out0[0:0];
assign v$SEL1_13506_out0 = v$IN_15104_out0[0:0];
assign v$G10_1380_out0 = !(v$SEL1_13459_out0 || v$SEL2_7670_out0);
assign v$G10_1381_out0 = !(v$SEL1_13460_out0 || v$SEL2_7671_out0);
assign v$G10_1382_out0 = !(v$SEL1_13461_out0 || v$SEL2_7672_out0);
assign v$G10_1383_out0 = !(v$SEL1_13462_out0 || v$SEL2_7673_out0);
assign v$G10_1384_out0 = !(v$SEL1_13463_out0 || v$SEL2_7674_out0);
assign v$G10_1385_out0 = !(v$SEL1_13464_out0 || v$SEL2_7675_out0);
assign v$G10_1422_out0 = !(v$SEL1_13501_out0 || v$SEL2_7712_out0);
assign v$G10_1423_out0 = !(v$SEL1_13502_out0 || v$SEL2_7713_out0);
assign v$G10_1424_out0 = !(v$SEL1_13503_out0 || v$SEL2_7714_out0);
assign v$G10_1425_out0 = !(v$SEL1_13504_out0 || v$SEL2_7715_out0);
assign v$G10_1426_out0 = !(v$SEL1_13505_out0 || v$SEL2_7716_out0);
assign v$G10_1427_out0 = !(v$SEL1_13506_out0 || v$SEL2_7717_out0);
assign v$MUX1_2390_out0 = v$LEFT$SHIT_3082_out0 ? v$_4286_out0 : v$_9021_out0;
assign v$MUX1_2396_out0 = v$LEFT$SHIT_3088_out0 ? v$_4292_out0 : v$_9027_out0;
assign v$G6_3555_out0 = ! v$SEL2_7670_out0;
assign v$G6_3556_out0 = ! v$SEL2_7671_out0;
assign v$G6_3557_out0 = ! v$SEL2_7672_out0;
assign v$G6_3558_out0 = ! v$SEL2_7673_out0;
assign v$G6_3559_out0 = ! v$SEL2_7674_out0;
assign v$G6_3560_out0 = ! v$SEL2_7675_out0;
assign v$G6_3597_out0 = ! v$SEL2_7712_out0;
assign v$G6_3598_out0 = ! v$SEL2_7713_out0;
assign v$G6_3599_out0 = ! v$SEL2_7714_out0;
assign v$G6_3600_out0 = ! v$SEL2_7715_out0;
assign v$G6_3601_out0 = ! v$SEL2_7716_out0;
assign v$G6_3602_out0 = ! v$SEL2_7717_out0;
assign v$G5_5831_out0 = ! v$SEL4_6079_out0;
assign v$G5_5832_out0 = ! v$SEL4_6080_out0;
assign v$G5_5833_out0 = ! v$SEL4_6081_out0;
assign v$G5_5834_out0 = ! v$SEL4_6082_out0;
assign v$G5_5835_out0 = ! v$SEL4_6083_out0;
assign v$G5_5836_out0 = ! v$SEL4_6084_out0;
assign v$G5_5873_out0 = ! v$SEL4_6121_out0;
assign v$G5_5874_out0 = ! v$SEL4_6122_out0;
assign v$G5_5875_out0 = ! v$SEL4_6123_out0;
assign v$G5_5876_out0 = ! v$SEL4_6124_out0;
assign v$G5_5877_out0 = ! v$SEL4_6125_out0;
assign v$G5_5878_out0 = ! v$SEL4_6126_out0;
assign v$G11_8842_out0 = !(v$SEL3_2294_out0 || v$SEL4_6079_out0);
assign v$G11_8843_out0 = !(v$SEL3_2295_out0 || v$SEL4_6080_out0);
assign v$G11_8844_out0 = !(v$SEL3_2296_out0 || v$SEL4_6081_out0);
assign v$G11_8845_out0 = !(v$SEL3_2297_out0 || v$SEL4_6082_out0);
assign v$G11_8846_out0 = !(v$SEL3_2298_out0 || v$SEL4_6083_out0);
assign v$G11_8847_out0 = !(v$SEL3_2299_out0 || v$SEL4_6084_out0);
assign v$G11_8884_out0 = !(v$SEL3_2336_out0 || v$SEL4_6121_out0);
assign v$G11_8885_out0 = !(v$SEL3_2337_out0 || v$SEL4_6122_out0);
assign v$G11_8886_out0 = !(v$SEL3_2338_out0 || v$SEL4_6123_out0);
assign v$G11_8887_out0 = !(v$SEL3_2339_out0 || v$SEL4_6124_out0);
assign v$G11_8888_out0 = !(v$SEL3_2340_out0 || v$SEL4_6125_out0);
assign v$G11_8889_out0 = !(v$SEL3_2341_out0 || v$SEL4_6126_out0);
assign v$G8_11990_out0 = ! v$SEL3_2294_out0;
assign v$G8_11991_out0 = ! v$SEL3_2295_out0;
assign v$G8_11992_out0 = ! v$SEL3_2296_out0;
assign v$G8_11993_out0 = ! v$SEL3_2297_out0;
assign v$G8_11994_out0 = ! v$SEL3_2298_out0;
assign v$G8_11995_out0 = ! v$SEL3_2299_out0;
assign v$G8_12032_out0 = ! v$SEL3_2336_out0;
assign v$G8_12033_out0 = ! v$SEL3_2337_out0;
assign v$G8_12034_out0 = ! v$SEL3_2338_out0;
assign v$G8_12035_out0 = ! v$SEL3_2339_out0;
assign v$G8_12036_out0 = ! v$SEL3_2340_out0;
assign v$G8_12037_out0 = ! v$SEL3_2341_out0;
assign v$G3_12662_out0 = v$G10_1380_out0 && v$G11_8842_out0;
assign v$G3_12663_out0 = v$G10_1381_out0 && v$G11_8843_out0;
assign v$G3_12664_out0 = v$G10_1382_out0 && v$G11_8844_out0;
assign v$G3_12665_out0 = v$G10_1383_out0 && v$G11_8845_out0;
assign v$G3_12666_out0 = v$G10_1384_out0 && v$G11_8846_out0;
assign v$G3_12667_out0 = v$G10_1385_out0 && v$G11_8847_out0;
assign v$G3_12704_out0 = v$G10_1422_out0 && v$G11_8884_out0;
assign v$G3_12705_out0 = v$G10_1423_out0 && v$G11_8885_out0;
assign v$G3_12706_out0 = v$G10_1424_out0 && v$G11_8886_out0;
assign v$G3_12707_out0 = v$G10_1425_out0 && v$G11_8887_out0;
assign v$G3_12708_out0 = v$G10_1426_out0 && v$G11_8888_out0;
assign v$G3_12709_out0 = v$G10_1427_out0 && v$G11_8889_out0;
assign v$MUX2_15241_out0 = v$EN_4758_out0 ? v$MUX1_2390_out0 : v$IN_15610_out0;
assign v$MUX2_15242_out0 = v$EN_4759_out0 ? v$MUX1_2396_out0 : v$IN_15611_out0;
assign v$G9_17588_out0 = v$G8_11990_out0 && v$G5_5831_out0;
assign v$G9_17589_out0 = v$G8_11991_out0 && v$G5_5832_out0;
assign v$G9_17590_out0 = v$G8_11992_out0 && v$G5_5833_out0;
assign v$G9_17591_out0 = v$G8_11993_out0 && v$G5_5834_out0;
assign v$G9_17592_out0 = v$G8_11994_out0 && v$G5_5835_out0;
assign v$G9_17593_out0 = v$G8_11995_out0 && v$G5_5836_out0;
assign v$G9_17630_out0 = v$G8_12032_out0 && v$G5_5873_out0;
assign v$G9_17631_out0 = v$G8_12033_out0 && v$G5_5874_out0;
assign v$G9_17632_out0 = v$G8_12034_out0 && v$G5_5875_out0;
assign v$G9_17633_out0 = v$G8_12035_out0 && v$G5_5876_out0;
assign v$G9_17634_out0 = v$G8_12036_out0 && v$G5_5877_out0;
assign v$G9_17635_out0 = v$G8_12037_out0 && v$G5_5878_out0;
assign v$G7_18131_out0 = v$G6_3555_out0 || v$SEL3_2294_out0;
assign v$G7_18132_out0 = v$G6_3556_out0 || v$SEL3_2295_out0;
assign v$G7_18133_out0 = v$G6_3557_out0 || v$SEL3_2296_out0;
assign v$G7_18134_out0 = v$G6_3558_out0 || v$SEL3_2297_out0;
assign v$G7_18135_out0 = v$G6_3559_out0 || v$SEL3_2298_out0;
assign v$G7_18136_out0 = v$G6_3560_out0 || v$SEL3_2299_out0;
assign v$G7_18173_out0 = v$G6_3597_out0 || v$SEL3_2336_out0;
assign v$G7_18174_out0 = v$G6_3598_out0 || v$SEL3_2337_out0;
assign v$G7_18175_out0 = v$G6_3599_out0 || v$SEL3_2338_out0;
assign v$G7_18176_out0 = v$G6_3600_out0 || v$SEL3_2339_out0;
assign v$G7_18177_out0 = v$G6_3601_out0 || v$SEL3_2340_out0;
assign v$G7_18178_out0 = v$G6_3602_out0 || v$SEL3_2341_out0;
assign v$Z_12553_out0 = v$G3_12662_out0;
assign v$Z_12554_out0 = v$G3_12663_out0;
assign v$Z_12555_out0 = v$G3_12664_out0;
assign v$Z_12556_out0 = v$G3_12665_out0;
assign v$Z_12557_out0 = v$G3_12666_out0;
assign v$Z_12558_out0 = v$G3_12667_out0;
assign v$Z_12595_out0 = v$G3_12704_out0;
assign v$Z_12596_out0 = v$G3_12705_out0;
assign v$Z_12597_out0 = v$G3_12706_out0;
assign v$Z_12598_out0 = v$G3_12707_out0;
assign v$Z_12599_out0 = v$G3_12708_out0;
assign v$Z_12600_out0 = v$G3_12709_out0;
assign v$OUT_14942_out0 = v$MUX2_15241_out0;
assign v$OUT_14948_out0 = v$MUX2_15242_out0;
assign v$G4_17523_out0 = v$G7_18131_out0 && v$G5_5831_out0;
assign v$G4_17524_out0 = v$G7_18132_out0 && v$G5_5832_out0;
assign v$G4_17525_out0 = v$G7_18133_out0 && v$G5_5833_out0;
assign v$G4_17526_out0 = v$G7_18134_out0 && v$G5_5834_out0;
assign v$G4_17527_out0 = v$G7_18135_out0 && v$G5_5835_out0;
assign v$G4_17528_out0 = v$G7_18136_out0 && v$G5_5836_out0;
assign v$G4_17565_out0 = v$G7_18173_out0 && v$G5_5873_out0;
assign v$G4_17566_out0 = v$G7_18174_out0 && v$G5_5874_out0;
assign v$G4_17567_out0 = v$G7_18175_out0 && v$G5_5875_out0;
assign v$G4_17568_out0 = v$G7_18176_out0 && v$G5_5876_out0;
assign v$G4_17569_out0 = v$G7_18177_out0 && v$G5_5877_out0;
assign v$G4_17570_out0 = v$G7_18178_out0 && v$G5_5878_out0;
assign v$Z2_179_out0 = v$Z_12553_out0;
assign v$Z2_180_out0 = v$Z_12555_out0;
assign v$Z2_181_out0 = v$Z_12557_out0;
assign v$Z2_184_out0 = v$Z_12595_out0;
assign v$Z2_185_out0 = v$Z_12597_out0;
assign v$Z2_186_out0 = v$Z_12599_out0;
assign v$IN_5184_out0 = v$OUT_14942_out0;
assign v$IN_5190_out0 = v$OUT_14948_out0;
assign v$Z1_5764_out0 = v$Z_12554_out0;
assign v$Z1_5765_out0 = v$Z_12556_out0;
assign v$Z1_5766_out0 = v$Z_12558_out0;
assign v$Z1_5769_out0 = v$Z_12596_out0;
assign v$Z1_5770_out0 = v$Z_12598_out0;
assign v$Z1_5771_out0 = v$Z_12600_out0;
assign v$_6266_out0 = { v$G4_17523_out0,v$G9_17588_out0 };
assign v$_6267_out0 = { v$G4_17524_out0,v$G9_17589_out0 };
assign v$_6268_out0 = { v$G4_17525_out0,v$G9_17590_out0 };
assign v$_6269_out0 = { v$G4_17526_out0,v$G9_17591_out0 };
assign v$_6270_out0 = { v$G4_17527_out0,v$G9_17592_out0 };
assign v$_6271_out0 = { v$G4_17528_out0,v$G9_17593_out0 };
assign v$_6308_out0 = { v$G4_17565_out0,v$G9_17630_out0 };
assign v$_6309_out0 = { v$G4_17566_out0,v$G9_17631_out0 };
assign v$_6310_out0 = { v$G4_17567_out0,v$G9_17632_out0 };
assign v$_6311_out0 = { v$G4_17568_out0,v$G9_17633_out0 };
assign v$_6312_out0 = { v$G4_17569_out0,v$G9_17634_out0 };
assign v$_6313_out0 = { v$G4_17570_out0,v$G9_17635_out0 };
assign v$IN_5030_out0 = v$IN_5184_out0;
assign v$IN_5031_out0 = v$IN_5190_out0;
assign v$Y_6483_out0 = v$_6266_out0;
assign v$Y_6484_out0 = v$_6267_out0;
assign v$Y_6485_out0 = v$_6268_out0;
assign v$Y_6486_out0 = v$_6269_out0;
assign v$Y_6487_out0 = v$_6270_out0;
assign v$Y_6488_out0 = v$_6271_out0;
assign v$Y_6525_out0 = v$_6308_out0;
assign v$Y_6526_out0 = v$_6309_out0;
assign v$Y_6527_out0 = v$_6310_out0;
assign v$Y_6528_out0 = v$_6311_out0;
assign v$Y_6529_out0 = v$_6312_out0;
assign v$Y_6530_out0 = v$_6313_out0;
assign v$G1_14591_out0 = v$Z1_5764_out0 && v$Z2_179_out0;
assign v$G1_14592_out0 = v$Z1_5765_out0 && v$Z2_180_out0;
assign v$G1_14593_out0 = v$Z1_5766_out0 && v$Z2_181_out0;
assign v$G1_14596_out0 = v$Z1_5769_out0 && v$Z2_184_out0;
assign v$G1_14597_out0 = v$Z1_5770_out0 && v$Z2_185_out0;
assign v$G1_14598_out0 = v$Z1_5771_out0 && v$Z2_186_out0;
assign v$_5466_out0 = { v$Y_6484_out0,v$C1_17666_out0 };
assign v$_5467_out0 = { v$Y_6486_out0,v$C1_17667_out0 };
assign v$_5468_out0 = { v$Y_6488_out0,v$C1_17668_out0 };
assign v$_5471_out0 = { v$Y_6526_out0,v$C1_17671_out0 };
assign v$_5472_out0 = { v$Y_6528_out0,v$C1_17672_out0 };
assign v$_5473_out0 = { v$Y_6530_out0,v$C1_17673_out0 };
assign v$_8148_out0 = { v$Y_6483_out0,v$C2_7624_out0 };
assign v$_8149_out0 = { v$Y_6485_out0,v$C2_7625_out0 };
assign v$_8150_out0 = { v$Y_6487_out0,v$C2_7626_out0 };
assign v$_8153_out0 = { v$Y_6525_out0,v$C2_7629_out0 };
assign v$_8154_out0 = { v$Y_6527_out0,v$C2_7630_out0 };
assign v$_8155_out0 = { v$Y_6529_out0,v$C2_7631_out0 };
assign v$SEL1_8732_out0 = v$IN_5030_out0[47:8];
assign v$SEL1_8738_out0 = v$IN_5031_out0[47:8];
assign v$Z_10329_out0 = v$G1_14591_out0;
assign v$Z_10330_out0 = v$G1_14592_out0;
assign v$Z_10331_out0 = v$G1_14593_out0;
assign v$Z_10334_out0 = v$G1_14596_out0;
assign v$Z_10335_out0 = v$G1_14597_out0;
assign v$Z_10336_out0 = v$G1_14598_out0;
assign v$SEL1_15423_out0 = v$IN_5030_out0[39:0];
assign v$SEL1_15429_out0 = v$IN_5031_out0[39:0];
assign v$Z2_2256_out0 = v$Z_10330_out0;
assign v$Z2_2257_out0 = v$Z_10335_out0;
assign v$_4282_out0 = { v$C2_140_out0,v$SEL1_15423_out0 };
assign v$_4288_out0 = { v$C2_146_out0,v$SEL1_15429_out0 };
assign v$_9017_out0 = { v$SEL1_8732_out0,v$C1_5998_out0 };
assign v$_9023_out0 = { v$SEL1_8738_out0,v$C1_6004_out0 };
assign v$Z3_11986_out0 = v$Z_10329_out0;
assign v$Z3_11987_out0 = v$Z_10334_out0;
assign v$MUX1_14693_out0 = v$Z1_5764_out0 ? v$_8148_out0 : v$_5466_out0;
assign v$MUX1_14694_out0 = v$Z1_5765_out0 ? v$_8149_out0 : v$_5467_out0;
assign v$MUX1_14695_out0 = v$Z1_5766_out0 ? v$_8150_out0 : v$_5468_out0;
assign v$MUX1_14698_out0 = v$Z1_5769_out0 ? v$_8153_out0 : v$_5471_out0;
assign v$MUX1_14699_out0 = v$Z1_5770_out0 ? v$_8154_out0 : v$_5472_out0;
assign v$MUX1_14700_out0 = v$Z1_5771_out0 ? v$_8155_out0 : v$_5473_out0;
assign v$Z1_17723_out0 = v$Z_10331_out0;
assign v$Z1_17724_out0 = v$Z_10336_out0;
assign v$MUX1_2386_out0 = v$LEFT$SHIT_3078_out0 ? v$_4282_out0 : v$_9017_out0;
assign v$MUX1_2392_out0 = v$LEFT$SHIT_3084_out0 ? v$_4288_out0 : v$_9023_out0;
assign v$Y_7756_out0 = v$MUX1_14693_out0;
assign v$Y_7757_out0 = v$MUX1_14694_out0;
assign v$Y_7758_out0 = v$MUX1_14695_out0;
assign v$Y_7761_out0 = v$MUX1_14698_out0;
assign v$Y_7762_out0 = v$MUX1_14699_out0;
assign v$Y_7763_out0 = v$MUX1_14700_out0;
assign v$G2_15863_out0 = v$Z2_2256_out0 && v$Z3_11986_out0;
assign v$G2_15864_out0 = v$Z2_2257_out0 && v$Z3_11987_out0;
assign v$_1325_out0 = { v$Y_7758_out0,v$C1_7724_out0 };
assign v$_1326_out0 = { v$Y_7763_out0,v$C1_7725_out0 };
assign v$MUX2_2504_out0 = v$EN_1343_out0 ? v$MUX1_2386_out0 : v$IN_5030_out0;
assign v$MUX2_2505_out0 = v$EN_1344_out0 ? v$MUX1_2392_out0 : v$IN_5031_out0;
assign v$_2675_out0 = { v$Y_7757_out0,v$C2_13386_out0 };
assign v$_2676_out0 = { v$Y_7762_out0,v$C2_13387_out0 };
assign v$_3328_out0 = { v$Y_7756_out0,v$C4_16302_out0 };
assign v$_3329_out0 = { v$Y_7761_out0,v$C4_16303_out0 };
assign v$G1_17016_out0 = v$Z1_17723_out0 && v$G2_15863_out0;
assign v$G1_17017_out0 = v$Z1_17724_out0 && v$G2_15864_out0;
assign v$Z_13551_out0 = v$G1_17016_out0;
assign v$Z_13552_out0 = v$G1_17017_out0;
assign v$OUT_14938_out0 = v$MUX2_2504_out0;
assign v$OUT_14944_out0 = v$MUX2_2505_out0;
assign v$MUX1_15287_out0 = v$Z2_2256_out0 ? v$_1325_out0 : v$_2675_out0;
assign v$MUX1_15288_out0 = v$Z2_2257_out0 ? v$_1326_out0 : v$_2676_out0;
assign v$IN_5186_out0 = v$OUT_14938_out0;
assign v$IN_5192_out0 = v$OUT_14944_out0;
assign v$MUX2_13544_out0 = v$Z3_11986_out0 ? v$MUX1_15287_out0 : v$_3328_out0;
assign v$MUX2_13545_out0 = v$Z3_11987_out0 ? v$MUX1_15288_out0 : v$_3329_out0;
assign v$IS$SUM$0_15623_out0 = v$Z_13551_out0;
assign v$IS$SUM$0_15624_out0 = v$Z_13552_out0;
assign v$IN_3867_out0 = v$IN_5186_out0;
assign v$IN_3870_out0 = v$IN_5192_out0;
assign v$OUT_8923_out0 = v$MUX2_13544_out0;
assign v$OUT_8924_out0 = v$MUX2_13545_out0;
assign v$IS$SUM$0_15681_out0 = v$IS$SUM$0_15623_out0;
assign v$IS$SUM$0_15682_out0 = v$IS$SUM$0_15624_out0;
assign v$IS$SUM$0_897_out0 = v$IS$SUM$0_15681_out0;
assign v$IS$SUM$0_898_out0 = v$IS$SUM$0_15682_out0;
assign v$SEL1_8734_out0 = v$IN_3867_out0[47:16];
assign v$SEL1_8740_out0 = v$IN_3870_out0[47:16];
assign v$_10370_out0 = { v$OUT_8923_out0,v$C10_13540_out0 };
assign v$_10371_out0 = { v$OUT_8924_out0,v$C10_13541_out0 };
assign v$SEL1_15425_out0 = v$IN_3867_out0[31:0];
assign v$SEL1_15431_out0 = v$IN_3870_out0[31:0];
assign v$NORMALIZATION$SHIFT_3253_out0 = v$_10370_out0;
assign v$NORMALIZATION$SHIFT_3254_out0 = v$_10371_out0;
assign v$_4284_out0 = { v$C2_142_out0,v$SEL1_15425_out0 };
assign v$_4290_out0 = { v$C2_148_out0,v$SEL1_15431_out0 };
assign v$_9019_out0 = { v$SEL1_8734_out0,v$C1_6000_out0 };
assign v$_9025_out0 = { v$SEL1_8740_out0,v$C1_6006_out0 };
assign v$NORMALIZATION$SHIFT_1165_out0 = v$NORMALIZATION$SHIFT_3253_out0;
assign v$NORMALIZATION$SHIFT_1166_out0 = v$NORMALIZATION$SHIFT_3254_out0;
assign v$MUX1_2388_out0 = v$LEFT$SHIT_3080_out0 ? v$_4284_out0 : v$_9019_out0;
assign v$MUX1_2394_out0 = v$LEFT$SHIT_3086_out0 ? v$_4290_out0 : v$_9025_out0;
assign v$SHIFT$AMOUNT_7389_out0 = v$NORMALIZATION$SHIFT_3253_out0;
assign v$SHIFT$AMOUNT_7394_out0 = v$NORMALIZATION$SHIFT_3254_out0;
assign v$SEL3_1139_out0 = v$SHIFT$AMOUNT_7389_out0[2:2];
assign v$SEL3_1144_out0 = v$SHIFT$AMOUNT_7394_out0[2:2];
assign v$SEL1_2271_out0 = v$SHIFT$AMOUNT_7389_out0[0:0];
assign v$SEL1_2276_out0 = v$SHIFT$AMOUNT_7394_out0[0:0];
assign v$SEL4_4939_out0 = v$SHIFT$AMOUNT_7389_out0[3:3];
assign v$SEL4_4944_out0 = v$SHIFT$AMOUNT_7394_out0[3:3];
assign v$SEL7_6347_out0 = v$SHIFT$AMOUNT_7389_out0[5:5];
assign v$SEL7_6352_out0 = v$SHIFT$AMOUNT_7394_out0[5:5];
assign v$SEL5_12217_out0 = v$SHIFT$AMOUNT_7389_out0[4:4];
assign v$SEL5_12222_out0 = v$SHIFT$AMOUNT_7394_out0[4:4];
assign v$SEL6_13781_out0 = v$SHIFT$AMOUNT_7389_out0[6:6];
assign v$SEL6_13786_out0 = v$SHIFT$AMOUNT_7394_out0[6:6];
assign v$SEL8_16572_out0 = v$SHIFT$AMOUNT_7389_out0[7:7];
assign v$SEL8_16577_out0 = v$SHIFT$AMOUNT_7394_out0[7:7];
assign v$SEL2_18357_out0 = v$SHIFT$AMOUNT_7389_out0[1:1];
assign v$SEL2_18362_out0 = v$SHIFT$AMOUNT_7394_out0[1:1];
assign v$MUX2_18581_out0 = v$EN_5218_out0 ? v$MUX1_2388_out0 : v$IN_3867_out0;
assign v$MUX2_18584_out0 = v$EN_5221_out0 ? v$MUX1_2394_out0 : v$IN_3870_out0;
assign v$NORMALIZATION$SHIFT_18622_out0 = v$NORMALIZATION$SHIFT_1165_out0;
assign v$NORMALIZATION$SHIFT_18623_out0 = v$NORMALIZATION$SHIFT_1166_out0;
assign v$EN_1335_out0 = v$SEL5_12217_out0;
assign v$EN_1336_out0 = v$SEL4_4939_out0;
assign v$EN_1349_out0 = v$SEL5_12222_out0;
assign v$EN_1350_out0 = v$SEL4_4944_out0;
assign v$EN_4753_out0 = v$SEL3_1139_out0;
assign v$EN_4762_out0 = v$SEL3_1144_out0;
assign v$EN_5212_out0 = v$SEL1_2271_out0;
assign v$EN_5225_out0 = v$SEL1_2276_out0;
assign v$EN_7875_out0 = v$SEL2_18357_out0;
assign v$EN_7884_out0 = v$SEL2_18362_out0;
assign v$SEL14_9100_out0 = v$NORMALIZATION$SHIFT_18622_out0[4:0];
assign v$SEL14_9101_out0 = v$NORMALIZATION$SHIFT_18623_out0[4:0];
assign v$NORMALIZATION$SHIFT_10742_out0 = v$NORMALIZATION$SHIFT_18622_out0;
assign v$NORMALIZATION$SHIFT_10743_out0 = v$NORMALIZATION$SHIFT_18623_out0;
assign v$OUT_14940_out0 = v$MUX2_18581_out0;
assign v$OUT_14946_out0 = v$MUX2_18584_out0;
assign v$G1_16031_out0 = v$SEL7_6347_out0 || v$SEL6_13781_out0;
assign v$G1_16036_out0 = v$SEL7_6352_out0 || v$SEL6_13786_out0;
assign v$NORMALIZATION$SHIFT_4397_out0 = v$SEL14_9100_out0;
assign v$NORMALIZATION$SHIFT_4398_out0 = v$SEL14_9101_out0;
assign v$IN_5183_out0 = v$OUT_14940_out0;
assign v$IN_5189_out0 = v$OUT_14946_out0;
assign v$XOR1_14547_out0 = v$NORMALIZATION$SHIFT_10742_out0 ^ v$C1_1555_out0;
assign v$XOR1_14548_out0 = v$NORMALIZATION$SHIFT_10743_out0 ^ v$C1_1556_out0;
assign v$G2_17413_out0 = v$G1_16031_out0 || v$SEL8_16572_out0;
assign v$G2_17418_out0 = v$G1_16036_out0 || v$SEL8_16577_out0;
assign v$MUX2_18575_out0 = v$EN_5212_out0 ? v$MUX1_2361_out0 : v$IN_3858_out0;
assign v$MUX2_18588_out0 = v$EN_5225_out0 ? v$MUX1_2409_out0 : v$IN_3874_out0;
assign {v$A1_638_out1,v$A1_638_out0 } = v$EXPONENT_1358_out0 + v$XOR1_14547_out0 + v$C2_2975_out0;
assign {v$A1_639_out1,v$A1_639_out0 } = v$EXPONENT_1359_out0 + v$XOR1_14548_out0 + v$C2_2976_out0;
assign v$IN_3866_out0 = v$IN_5183_out0;
assign v$IN_3869_out0 = v$IN_5189_out0;
assign v$XOR1_10930_out0 = v$NORMALIZATION$SHIFT_4397_out0 ^ v$C1_15734_out0;
assign v$XOR1_10931_out0 = v$NORMALIZATION$SHIFT_4398_out0 ^ v$C1_15735_out0;
assign v$OUT_14913_out0 = v$MUX2_18575_out0;
assign v$OUT_14961_out0 = v$MUX2_18588_out0;
assign v$IN_5161_out0 = v$OUT_14913_out0;
assign v$IN_5209_out0 = v$OUT_14961_out0;
assign {v$A1_7730_out1,v$A1_7730_out0 } = v$EXPONENT_16395_out0 + v$XOR1_10930_out0 + v$C2_1456_out0;
assign {v$A1_7731_out1,v$A1_7731_out0 } = v$EXPONENT_16396_out0 + v$XOR1_10931_out0 + v$C2_1457_out0;
assign v$SEL1_8731_out0 = v$IN_3866_out0[47:32];
assign v$SEL1_8737_out0 = v$IN_3869_out0[47:32];
assign v$IGNORE_11704_out0 = v$A1_638_out1;
assign v$IGNORE_11705_out0 = v$A1_639_out1;
assign v$SEL1_15422_out0 = v$IN_3866_out0[15:0];
assign v$SEL1_15428_out0 = v$IN_3869_out0[15:0];
assign v$OUT_16097_out0 = v$A1_638_out0;
assign v$OUT_16098_out0 = v$A1_639_out0;
assign v$_4281_out0 = { v$C2_139_out0,v$SEL1_15422_out0 };
assign v$_4287_out0 = { v$C2_145_out0,v$SEL1_15428_out0 };
assign v$OUT_6193_out0 = v$A1_7730_out0;
assign v$OUT_6194_out0 = v$A1_7731_out0;
assign v$_9016_out0 = { v$SEL1_8731_out0,v$C1_5997_out0 };
assign v$_9022_out0 = { v$SEL1_8737_out0,v$C1_6003_out0 };
assign v$IN_11783_out0 = v$IN_5161_out0;
assign v$IN_11792_out0 = v$IN_5209_out0;
assign v$IGNORE_16561_out0 = v$A1_7730_out1;
assign v$IGNORE_16562_out0 = v$A1_7731_out1;
assign v$MUX1_2385_out0 = v$LEFT$SHIT_3077_out0 ? v$_4281_out0 : v$_9016_out0;
assign v$MUX1_2391_out0 = v$LEFT$SHIT_3083_out0 ? v$_4287_out0 : v$_9022_out0;
assign v$SEL1_8709_out0 = v$IN_11783_out0[23:2];
assign v$SEL1_8757_out0 = v$IN_11792_out0[23:2];
assign v$SEL1_15400_out0 = v$IN_11783_out0[21:0];
assign v$SEL1_15448_out0 = v$IN_11792_out0[21:0];
assign v$_4259_out0 = { v$C2_117_out0,v$SEL1_15400_out0 };
assign v$_4307_out0 = { v$C2_165_out0,v$SEL1_15448_out0 };
assign v$_8994_out0 = { v$SEL1_8709_out0,v$C1_5975_out0 };
assign v$_9042_out0 = { v$SEL1_8757_out0,v$C1_6023_out0 };
assign v$MUX2_18580_out0 = v$EN_5217_out0 ? v$MUX1_2385_out0 : v$IN_3866_out0;
assign v$MUX2_18583_out0 = v$EN_5220_out0 ? v$MUX1_2391_out0 : v$IN_3869_out0;
assign v$MUX1_2363_out0 = v$LEFT$SHIT_3055_out0 ? v$_4259_out0 : v$_8994_out0;
assign v$MUX1_2411_out0 = v$LEFT$SHIT_3103_out0 ? v$_4307_out0 : v$_9042_out0;
assign v$OUT_14937_out0 = v$MUX2_18580_out0;
assign v$OUT_14943_out0 = v$MUX2_18583_out0;
assign v$MUX2_2477_out0 = v$EN_7875_out0 ? v$MUX1_2363_out0 : v$IN_11783_out0;
assign v$MUX2_2486_out0 = v$EN_7884_out0 ? v$MUX1_2411_out0 : v$IN_11792_out0;
assign v$OUT_4915_out0 = v$OUT_14937_out0;
assign v$OUT_4916_out0 = v$OUT_14943_out0;
assign v$SEL2_8099_out0 = v$OUT_4915_out0[46:37];
assign v$SEL2_8100_out0 = v$OUT_4916_out0[46:24];
assign v$OUT_14915_out0 = v$MUX2_2477_out0;
assign v$OUT_14963_out0 = v$MUX2_2486_out0;
assign v$IN_5160_out0 = v$OUT_14915_out0;
assign v$IN_5208_out0 = v$OUT_14963_out0;
assign v$_15848_out0 = { v$SEL2_8099_out0,v$A2_10046_out0 };
assign v$_15849_out0 = { v$SEL2_8100_out0,v$A2_10047_out0 };
assign v$MUX2_13632_out0 = v$Z_15810_out0 ? v$C4_8258_out0 : v$_15848_out0;
assign v$MUX2_13633_out0 = v$Z_15811_out0 ? v$C4_8259_out0 : v$_15849_out0;
assign v$IN_15605_out0 = v$IN_5160_out0;
assign v$IN_15614_out0 = v$IN_5208_out0;
assign v$SEL1_8708_out0 = v$IN_15605_out0[23:4];
assign v$SEL1_8756_out0 = v$IN_15614_out0[23:4];
assign v$SEL1_15399_out0 = v$IN_15605_out0[19:0];
assign v$SEL1_15447_out0 = v$IN_15614_out0[19:0];
assign v$_18418_out0 = { v$MUX2_13632_out0,v$SIGN_1368_out0 };
assign v$_18419_out0 = { v$MUX2_13633_out0,v$SIGN_1369_out0 };
assign v$_4258_out0 = { v$C2_116_out0,v$SEL1_15399_out0 };
assign v$_4306_out0 = { v$C2_164_out0,v$SEL1_15447_out0 };
assign v$_8993_out0 = { v$SEL1_8708_out0,v$C1_5974_out0 };
assign v$_9041_out0 = { v$SEL1_8756_out0,v$C1_6022_out0 };
assign v$OUT_12480_out0 = v$_18418_out0;
assign v$OUT_12481_out0 = v$_18419_out0;
assign v$MUX1_2362_out0 = v$LEFT$SHIT_3054_out0 ? v$_4258_out0 : v$_8993_out0;
assign v$MUX1_2410_out0 = v$LEFT$SHIT_3102_out0 ? v$_4306_out0 : v$_9041_out0;
assign v$MUX11_8670_out0 = v$G5_6199_out0 ? v$C9_18761_out0 : v$OUT_12480_out0;
assign v$MUX3_8966_out0 = v$G3_16010_out0 ? v$C1_15227_out0 : v$OUT_12481_out0;
assign v$SINGLE$PRECISION_7901_out0 = v$MUX3_8966_out0;
assign v$MUX2_15236_out0 = v$EN_4753_out0 ? v$MUX1_2362_out0 : v$IN_15605_out0;
assign v$MUX2_15245_out0 = v$EN_4762_out0 ? v$MUX1_2410_out0 : v$IN_15614_out0;
assign v$_17037_out0 = { v$C10_6385_out0,v$MUX11_8670_out0 };
assign v$HALF$PRECISION_10312_out0 = v$_17037_out0;
assign v$OUT_14914_out0 = v$MUX2_15236_out0;
assign v$OUT_14962_out0 = v$MUX2_15245_out0;
assign v$IN_5158_out0 = v$OUT_14914_out0;
assign v$IN_5206_out0 = v$OUT_14962_out0;
assign v$MUX12_16797_out0 = v$IS$32$BITS_1282_out0 ? v$SINGLE$PRECISION_7901_out0 : v$HALF$PRECISION_10312_out0;
assign v$OUT_3365_out0 = v$MUX12_16797_out0;
assign v$IN_5023_out0 = v$IN_5158_out0;
assign v$IN_5037_out0 = v$IN_5206_out0;
assign v$SEL1_8706_out0 = v$IN_5023_out0[23:8];
assign v$SEL1_8754_out0 = v$IN_5037_out0[23:8];
assign v$SEL1_15397_out0 = v$IN_5023_out0[15:0];
assign v$SEL1_15445_out0 = v$IN_5037_out0[15:0];
assign v$_4256_out0 = { v$C2_114_out0,v$SEL1_15397_out0 };
assign v$_4304_out0 = { v$C2_162_out0,v$SEL1_15445_out0 };
assign v$_8991_out0 = { v$SEL1_8706_out0,v$C1_5972_out0 };
assign v$_9039_out0 = { v$SEL1_8754_out0,v$C1_6020_out0 };
assign v$MUX1_2360_out0 = v$LEFT$SHIT_3052_out0 ? v$_4256_out0 : v$_8991_out0;
assign v$MUX1_2408_out0 = v$LEFT$SHIT_3100_out0 ? v$_4304_out0 : v$_9039_out0;
assign v$MUX2_2497_out0 = v$EN_1336_out0 ? v$MUX1_2360_out0 : v$IN_5023_out0;
assign v$MUX2_2511_out0 = v$EN_1350_out0 ? v$MUX1_2408_out0 : v$IN_5037_out0;
assign v$OUT_14912_out0 = v$MUX2_2497_out0;
assign v$OUT_14960_out0 = v$MUX2_2511_out0;
assign v$IN_5157_out0 = v$OUT_14912_out0;
assign v$IN_5205_out0 = v$OUT_14960_out0;
assign v$IN_5022_out0 = v$IN_5157_out0;
assign v$IN_5036_out0 = v$IN_5205_out0;
assign v$SEL1_8705_out0 = v$IN_5022_out0[23:16];
assign v$SEL1_8753_out0 = v$IN_5036_out0[23:16];
assign v$SEL1_15396_out0 = v$IN_5022_out0[7:0];
assign v$SEL1_15444_out0 = v$IN_5036_out0[7:0];
assign v$_4255_out0 = { v$C2_113_out0,v$SEL1_15396_out0 };
assign v$_4303_out0 = { v$C2_161_out0,v$SEL1_15444_out0 };
assign v$_8990_out0 = { v$SEL1_8705_out0,v$C1_5971_out0 };
assign v$_9038_out0 = { v$SEL1_8753_out0,v$C1_6019_out0 };
assign v$MUX1_2359_out0 = v$LEFT$SHIT_3051_out0 ? v$_4255_out0 : v$_8990_out0;
assign v$MUX1_2407_out0 = v$LEFT$SHIT_3099_out0 ? v$_4303_out0 : v$_9038_out0;
assign v$MUX2_2496_out0 = v$EN_1335_out0 ? v$MUX1_2359_out0 : v$IN_5022_out0;
assign v$MUX2_2510_out0 = v$EN_1349_out0 ? v$MUX1_2407_out0 : v$IN_5036_out0;
assign v$OUT_14911_out0 = v$MUX2_2496_out0;
assign v$OUT_14959_out0 = v$MUX2_2510_out0;
assign v$MUX1_11632_out0 = v$G2_17413_out0 ? v$C1_4456_out0 : v$OUT_14911_out0;
assign v$MUX1_11637_out0 = v$G2_17418_out0 ? v$C1_4461_out0 : v$OUT_14959_out0;
assign v$OUT_10013_out0 = v$MUX1_11632_out0;
assign v$OUT_10018_out0 = v$MUX1_11637_out0;
assign v$SEL2_6033_out0 = v$OUT_10013_out0[22:0];
assign v$SEL2_6034_out0 = v$OUT_10018_out0[22:0];
assign v$MUX2_2973_out0 = v$IS$SUM$0_15623_out0 ? v$C5_15619_out0 : v$SEL2_6033_out0;
assign v$MUX2_2974_out0 = v$IS$SUM$0_15624_out0 ? v$C5_15620_out0 : v$SEL2_6034_out0;
assign v$MUX6_12770_out0 = v$IS$SUB_13067_out0 ? v$MUX2_2973_out0 : v$SEL3_14249_out0;
assign v$MUX6_12771_out0 = v$IS$SUB_13068_out0 ? v$MUX2_2974_out0 : v$SEL3_14250_out0;
assign v$OUT1_10407_out0 = v$MUX6_12770_out0;
assign v$OUT1_10408_out0 = v$MUX6_12771_out0;
assign v$MANTISA$RESULT_6546_out0 = v$OUT1_10407_out0;
assign v$MANTISA$RESULT_6547_out0 = v$OUT1_10408_out0;
assign v$SEL10_3207_out0 = v$MANTISA$RESULT_6546_out0[22:13];
assign v$SEL10_3208_out0 = v$MANTISA$RESULT_6547_out0[22:13];
assign v$SEL7_3274_out0 = v$MANTISA$RESULT_6546_out0[22:13];
assign v$SEL7_3275_out0 = v$MANTISA$RESULT_6547_out0[22:13];
assign v$_7021_out0 = { v$MANTISA$RESULT_6546_out0,v$OUT_14778_out0 };
assign v$_7022_out0 = { v$MANTISA$RESULT_6547_out0,v$OUT_14779_out0 };
assign v$_15351_out0 = { v$MANTISA$RESULT_6546_out0,v$OUT_16097_out0 };
assign v$_15352_out0 = { v$MANTISA$RESULT_6547_out0,v$OUT_16098_out0 };
assign v$_11383_out0 = { v$SEL10_3207_out0,v$OUT_6193_out0 };
assign v$_11384_out0 = { v$SEL10_3208_out0,v$OUT_6194_out0 };
assign v$_15153_out0 = { v$SEL7_3274_out0,v$OUT_170_out0 };
assign v$_15154_out0 = { v$SEL7_3275_out0,v$OUT_171_out0 };
assign v$_56_out0 = { v$C9_3300_out0,v$_11383_out0 };
assign v$_57_out0 = { v$C9_3301_out0,v$_11384_out0 };
assign v$_11831_out0 = { v$C7_1708_out0,v$_15153_out0 };
assign v$_11832_out0 = { v$C7_1709_out0,v$_15154_out0 };
assign v$MUX12_15140_out0 = v$IS$32$BIT_10862_out0 ? v$_7021_out0 : v$_11831_out0;
assign v$MUX12_15141_out0 = v$IS$32$BIT_10863_out0 ? v$_7022_out0 : v$_11832_out0;
assign v$MUX6_17434_out0 = v$IS$32$BIT_10862_out0 ? v$_15351_out0 : v$_56_out0;
assign v$MUX6_17435_out0 = v$IS$32$BIT_10863_out0 ? v$_15352_out0 : v$_57_out0;
assign v$_16507_out0 = { v$MUX12_15140_out0,v$SEL13_17581_out0 };
assign v$_16508_out0 = { v$MUX12_15141_out0,v$SEL13_17582_out0 };
assign v$_16799_out0 = { v$MUX6_17434_out0,v$SUBTRACTION$SIGN_11872_out0 };
assign v$_16800_out0 = { v$MUX6_17435_out0,v$SUBTRACTION$SIGN_11873_out0 };
assign v$MUX1_13555_out0 = v$IS$SUB_4443_out0 ? v$_16799_out0 : v$_16507_out0;
assign v$MUX1_13556_out0 = v$IS$SUB_4444_out0 ? v$_16800_out0 : v$_16508_out0;
assign v$MUX7_4863_out0 = v$IS$SUM$0_897_out0 ? v$C5_4112_out0 : v$MUX1_13555_out0;
assign v$MUX7_4864_out0 = v$IS$SUM$0_898_out0 ? v$C5_4113_out0 : v$MUX1_13556_out0;
assign v$OUT1_17809_out0 = v$MUX7_4863_out0;
assign v$OUT1_17810_out0 = v$MUX7_4864_out0;
assign v$MUX2_16229_out0 = v$G2_3724_out0 ? v$OUT1_17809_out0 : v$C4_14026_out0;
assign v$MUX2_16230_out0 = v$G2_3725_out0 ? v$OUT1_17810_out0 : v$C4_14027_out0;
assign v$MUX4_1257_out0 = v$FINISHED_8010_out0 ? v$OUT_3364_out0 : v$MUX2_16229_out0;
assign v$MUX4_1258_out0 = v$MUL_17035_out0 ? v$OUT_3365_out0 : v$MUX2_16230_out0;
assign v$SEL4_9556_out0 = v$MUX4_1257_out0[15:0];
assign v$SEL4_9557_out0 = v$MUX4_1258_out0[15:0];
assign v$SEL5_13590_out0 = v$MUX4_1257_out0[31:16];
assign v$SEL5_13591_out0 = v$MUX4_1258_out0[31:16];
assign v$MUX3_18386_out0 = v$G12_11978_out0 ? v$REG3_11767_out0 : v$SEL5_13590_out0;
assign v$MUX3_18387_out0 = v$G12_11979_out0 ? v$REG3_11768_out0 : v$SEL5_13591_out0;
assign v$OUT_1321_out0 = v$MUX3_18386_out0;
assign v$OUT_1322_out0 = v$MUX3_18387_out0;
assign v$FPU$OUT_17011_out0 = v$OUT_1321_out0;
assign v$FPU$OUT_17012_out0 = v$OUT_1322_out0;
assign v$MUX6_7439_out0 = v$G21_18680_out0 ? v$FPU$OUT_17011_out0 : v$MUX4_45_out0;
assign v$MUX6_7440_out0 = v$G21_18681_out0 ? v$FPU$OUT_17012_out0 : v$MUX4_46_out0;
assign v$DIN3_14419_out0 = v$MUX6_7440_out0;
assign v$MUX14_18722_out0 = v$FINISHED_13867_out0 ? v$FPU$OUT_17011_out0 : v$MUX6_7439_out0;
assign v$DIN3_14418_out0 = v$MUX14_18722_out0;


endmodule
